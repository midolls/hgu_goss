* NGSPICE file created from hgu_vgen_vref.ext - technology: sky130A

*.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 Y VGND 0.0998f
C1 VGND A 0.04f
C2 VPB Y 0.0177f
C3 VPB A 0.0451f
C4 VGND VPWR 0.0338f
C5 Y A 0.0476f
C6 VPB VPWR 0.0545f
C7 Y VPWR 0.128f
C8 A VPWR 0.037f
C9 VPB VGND 0.00948f
C10 VGND VNB 0.251f
C11 Y VNB 0.0961f
C12 VPWR VNB 0.219f
C13 A VNB 0.167f
C14 VPB VNB 0.339f
.ends

.subckt pfet_01v8_w500_l500_nf2 a_n29_0# a_129_0# a_n129_n26# w_n224_n36# a_n187_0#
+ a_29_n26# VSUBS
X0 a_129_0# a_29_n26# a_n29_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_0# a_n129_n26# a_n187_0# w_n224_n36# sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
C0 a_n187_0# a_n29_0# 0.0184f
C1 a_n29_0# a_n129_n26# 0.00388f
C2 a_n29_0# a_129_0# 0.0184f
C3 w_n224_n36# a_n187_0# 0.00201f
C4 w_n224_n36# a_n129_n26# 0.0302f
C5 a_n29_0# a_29_n26# 0.00388f
C6 a_n187_0# a_n129_n26# 0.00388f
C7 w_n224_n36# a_129_0# 0.002f
C8 w_n224_n36# a_29_n26# 0.0301f
C9 a_n129_n26# a_29_n26# 0.0143f
C10 a_29_n26# a_129_0# 0.00388f
C11 w_n224_n36# a_n29_0# 0.00149f
C12 a_129_0# VSUBS 0.0383f
C13 a_n29_0# VSUBS 0.0212f
C14 a_n187_0# VSUBS 0.0382f
C15 a_29_n26# VSUBS 0.114f
C16 a_n129_n26# VSUBS 0.114f
C17 w_n224_n36# VSUBS 0.233f
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 A VPWR 0.016f
C1 VPWR VGND 0.072f
C2 VPWR X 0.333f
C3 VPWR VPB 0.0711f
C4 A VGND 0.0194f
C5 VPWR a_27_47# 0.218f
C6 A X 4.66e-19
C7 VGND X 0.23f
C8 A VPB 0.0361f
C9 VGND VPB 0.00796f
C10 A a_27_47# 0.17f
C11 a_27_47# VGND 0.163f
C12 VPB X 0.00899f
C13 a_27_47# X 0.207f
C14 a_27_47# VPB 0.132f
C15 VGND VNB 0.378f
C16 X VNB 0.039f
C17 VPWR VNB 0.325f
C18 A VNB 0.14f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.461f
.ends

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VPWR X a_240_47# VNB VPB a_629_47#
+ a_523_47# a_346_47# a_63_47#
X0 X a_629_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 a_523_47# a_346_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2 VGND a_240_47# a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_240_47# a_63_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VPWR a_240_47# a_346_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND A a_63_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR A a_63_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VPWR a_523_47# a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND a_523_47# a_629_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_523_47# a_346_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X10 a_240_47# a_63_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X11 X a_629_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
C0 a_523_47# a_629_47# 0.322f
C1 VGND A 0.0175f
C2 a_629_47# a_240_47# 7.09e-19
C3 a_523_47# X 0.00484f
C4 a_629_47# VPWR 0.13f
C5 VGND a_346_47# 0.121f
C6 VPWR X 0.0861f
C7 VPB VGND 0.00789f
C8 a_63_47# a_240_47# 0.16f
C9 a_63_47# VPWR 0.15f
C10 a_523_47# a_240_47# 0.0145f
C11 a_523_47# VPWR 0.081f
C12 a_629_47# VPB 0.0445f
C13 VPWR a_240_47# 0.0828f
C14 VPB X 0.0189f
C15 a_63_47# A 0.245f
C16 a_63_47# VPB 0.0507f
C17 a_523_47# a_346_47# 0.16f
C18 a_240_47# A 0.0146f
C19 VPWR A 0.0174f
C20 a_240_47# a_346_47# 0.319f
C21 a_523_47# VPB 0.116f
C22 VPWR a_346_47# 0.127f
C23 VPB a_240_47# 0.116f
C24 a_629_47# VGND 0.124f
C25 VPB VPWR 0.0985f
C26 X VGND 0.0832f
C27 A a_346_47# 6.53e-19
C28 a_63_47# VGND 0.144f
C29 VPB A 0.104f
C30 VPB a_346_47# 0.0439f
C31 a_523_47# VGND 0.0787f
C32 a_629_47# X 0.136f
C33 VGND a_240_47# 0.0806f
C34 VPWR VGND 0.0902f
C35 VGND VNB 0.539f
C36 X VNB 0.1f
C37 VPWR VNB 0.446f
C38 A VNB 0.198f
C39 VPB VNB 0.959f
C40 a_629_47# VNB 0.129f
C41 a_523_47# VNB 0.162f
C42 a_346_47# VNB 0.109f
C43 a_240_47# VNB 0.153f
C44 a_63_47# VNB 0.167f
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 nmoscap_top nmoscap_bot pwell sky130_fd_pr__cap_var_lvt w=16.4 l=16
X1 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=17.2 w=17.2
C0 mimcap_top nmoscap_bot 0.225f
C1 nmoscap_bot mimcap_bot 21.2f
C2 mimcap_top mimcap_bot 31.6f
C3 nmoscap_top nmoscap_bot 0.281p
C4 nmoscap_top mimcap_top 2.63f
C5 nmoscap_top mimcap_bot 19.2f
C6 mimcap_top pwell 2.84f
C7 mimcap_bot pwell 3.75f
C8 nmoscap_top pwell 8.6f
C9 nmoscap_bot pwell 40.7f
.ends

.subckt nfet_01v8_w500_l500_nf2 a_n129_n76# a_n29_n50# a_n187_n50# a_29_n76# a_129_n50#
+ VSUBS
X0 a_129_n50# a_29_n76# a_n29_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n76# a_n187_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
C0 a_n29_n50# a_129_n50# 0.0184f
C1 a_n29_n50# a_n129_n76# 0.00388f
C2 a_29_n76# a_129_n50# 0.00388f
C3 a_n129_n76# a_n187_n50# 0.00388f
C4 a_n29_n50# a_n187_n50# 0.0184f
C5 a_29_n76# a_n129_n76# 0.0143f
C6 a_29_n76# a_n29_n50# 0.00388f
C7 a_129_n50# VSUBS 0.0402f
C8 a_n29_n50# VSUBS 0.0227f
C9 a_n187_n50# VSUBS 0.0402f
C10 a_29_n76# VSUBS 0.144f
C11 a_n129_n76# VSUBS 0.144f
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 VPWR VGND 0.0322f
C1 VPWR VPB 0.0509f
C2 Y B 0.0481f
C3 Y a_113_47# 0.00937f
C4 B A 0.051f
C5 Y VGND 0.139f
C6 Y VPB 0.00618f
C7 A VGND 0.00949f
C8 A VPB 0.0379f
C9 B VGND 0.0544f
C10 B VPB 0.0391f
C11 a_113_47# VGND 0.0019f
C12 Y VPWR 0.211f
C13 A VPWR 0.0444f
C14 VPB VGND 0.0044f
C15 Y A 0.0855f
C16 B VPWR 0.0478f
C17 VPWR a_113_47# 1.78e-19
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt hgu_vgen_vref clk vcm VSS VDD
Xsky130_fd_sc_hd__inv_1_4 clk VSS VDD sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__inv_1
Xpfet_01v8_w500_l500_nf2_0 mimtop2 vcm phi1_n VDD vcm phi1_n VSS pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_1 mimtop1 vcm phi1_n VDD vcm phi1_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_0 sky130_fd_sc_hd__inv_1_2/A VSS VDD phi1 VSS VDD sky130_fd_sc_hd__buf_4_0/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_2 mimtop2 mimbot1 phi2_n VDD mimbot1 phi2_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_1 sky130_fd_sc_hd__inv_1_2/Y VSS VDD phi1_n VSS VDD sky130_fd_sc_hd__buf_4_1/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xpfet_01v8_w500_l500_nf2_3 VDD mimtop1 phi2_n VDD mimtop1 phi2_n VSS pfet_01v8_w500_l500_nf2
Xpfet_01v8_w500_l500_nf2_4 mimbot1 VSS phi1_n VDD VSS phi1_n VSS pfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__buf_4_2 sky130_fd_sc_hd__inv_1_3/A VSS VDD phi2 VSS VDD sky130_fd_sc_hd__buf_4_2/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_4_3 sky130_fd_sc_hd__inv_1_3/Y VSS VDD phi2_n VSS VDD sky130_fd_sc_hd__buf_4_3/a_27_47#
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dlymetal6s6s_1_0 sky130_fd_sc_hd__nand2_1_0/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_1 sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_2 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_3 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_0/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_5 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VSS VDD sky130_fd_sc_hd__inv_1_1/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xsky130_fd_sc_hd__dlymetal6s6s_1_4 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_5/A
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VSS VDD sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47#
+ sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|0] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|1] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|2] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|3] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7|4] vcm VSS mimtop2 VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|0] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|1] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|2] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|3] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[0|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[1|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[2|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[3|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[4|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[5|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[6|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_3[7|4] vcm VSS mimtop1 mimbot1 VSS adc_noise_decoup_cell1
Xnfet_01v8_w500_l500_nf2_0 phi1 mimtop2 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_1 phi1 mimtop1 vcm phi1 vcm VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_0 clk sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__nand2_1_0/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_2 phi2 mimtop2 mimbot1 phi2 mimbot1 VSS nfet_01v8_w500_l500_nf2
Xnfet_01v8_w500_l500_nf2_3 phi2 VDD mimtop1 phi2 mimtop1 VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_4/Y
+ VSS VDD sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xnfet_01v8_w500_l500_nf2_4 phi1 mimbot1 VSS phi1 VSS VSS nfet_01v8_w500_l500_nf2
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VSS VDD sky130_fd_sc_hd__inv_1_2/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A VSS VDD sky130_fd_sc_hd__inv_1_3/A
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VSS VDD sky130_fd_sc_hd__inv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A VSS VDD sky130_fd_sc_hd__inv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__inv_1
X0 VDD.t5 VSS sky130_fd_pr__cap_mim_m3_1 l=0 w=0
X1 vcm.t0 VSS.t1 error sky130_fd_pr__cap_var_lvt w=0 l=0
X2 vcm.t62 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X3 vcm.t67 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X4 vcm.t78 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X5 mimtop2 VSS.t0 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
X6 vcm.t25 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X7 vcm.t58 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X8 vcm.t74 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X9 vcm.t43 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X10 vcm.t54 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X11 vcm.t70 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X12 vcm.t50 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X13 vcm.t61 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X14 vcm.t66 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X15 vcm.t20 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X16 vcm.t46 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X17 vcm.t77 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X18 VDD.t3 VSS sky130_fd_pr__cap_mim_m3_1 l=0 w=0
X19 vcm.t2 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X20 vcm.t36 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X21 vcm.t42 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X22 VDD.t0 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X23 VDD.t4 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X24 vcm.t53 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X25 vcm.t12 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X26 vcm.t69 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X27 vcm.t23 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X28 vcm.t28 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X29 vcm.t39 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X30 vcm.t60 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X31 vcm.t76 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X32 VDD.t2 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X33 vcm.t1 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X34 vcm.t19 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X35 vcm.t35 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X36 vcm.t45 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X37 vcm.t4 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X38 sky130_fd_sc_hd__nand2_1_0/Y clk.t3 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
X39 vcm.t15 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X40 vcm.t31 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X41 vcm.t52 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X42 vcm.t63 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X43 vcm.t68 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X44 vcm.t11 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X45 vcm.t22 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X46 vcm.t27 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X47 vcm.t79 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X48 vcm.t7 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X49 vcm.t18 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X50 vcm.t38 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X51 vcm.t44 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X52 vcm.t55 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X53 vcm.t71 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X54 sky130_fd_sc_hd__inv_1_4/Y clk.t0 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0 l=0
X55 vcm.t3 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X56 vcm.t14 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X57 VDD.t1 VSS sky130_fd_pr__cap_mim_m3_1 l=0 w=0
X58 vcm.t30 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X59 vcm.t34 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X60 vcm.t21 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X61 vcm.t37 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X62 vcm.t47 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X63 vcm.t6 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X64 vcm.t17 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X65 vcm.t57 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X66 vcm.t13 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X67 vcm.t29 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X68 vcm.t33 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X69 vcm.t73 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X70 vcm.t8 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X71 vcm.t49 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X72 vcm.t5 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X73 vcm.t16 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X74 vcm.t24 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X75 vcm.t65 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X76 vcm.t32 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X77 vcm.t56 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X78 vcm.t72 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X79 vcm.t10 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X80 vcm.t41 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X81 VDD clk.t2 sky130_fd_sc_hd__nand2_1_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
X82 vcm.t48 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X83 vcm.t59 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X84 vcm.t64 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X85 sky130_fd_sc_hd__inv_1_4/Y clk.t1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=0 l=0
X86 vcm.t26 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X87 vcm.t75 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X88 vcm.t9 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X89 vcm.t40 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
X90 vcm.t51 VSS error sky130_fd_pr__cap_var_lvt w=0 l=0
R0 clk.n1 clk.t1 229.433
R1 clk.n0 clk.t2 229.04
R2 clk.n1 clk.t0 158.886
R3 clk.n0 clk.t3 158.46
R4 clk.n7 clk 38.8978
R5 clk.n8 clk.n0 8.7103
R6 clk.n2 clk.n1 7.39078
R7 clk.n4 clk.n3 3.46717
R8 clk clk.n8 3.16209
R9 clk.n6 clk.n4 3.03598
R10 clk.n7 clk.n6 2.61367
R11 clk.n8 clk.n7 2.26586
R12 clk.n4 clk.n2 1.06717
R13 clk.n3 clk 1.06717
R14 clk.n6 clk.n5 0.00666568
R15 VSS.n4945 VSS.n4944 34571.4
R16 VSS.n4814 VSS.n4812 34571.4
R17 VSS.n5108 VSS.n5107 34571.4
R18 VSS.n10411 VSS.n10410 32675.1
R19 VSS.n10530 VSS.n10524 32675.1
R20 VSS.n10522 VSS.n10520 32675.1
R21 VSS.n10515 VSS.n10253 32675.1
R22 VSS.n11347 VSS.n11346 23783
R23 VSS.n5108 VSS.n4745 22403.2
R24 VSS.n10202 VSS.n10201 21511.1
R25 VSS.n10484 VSS.n10483 21511.1
R26 VSS.n10189 VSS.n3684 21511.1
R27 VSS.n4877 VSS.n4872 21511.1
R28 VSS.n4953 VSS.n4951 21511.1
R29 VSS.n4809 VSS.n4801 21511.1
R30 VSS.n4875 VSS.n4551 21511.1
R31 VSS.n4903 VSS.n4900 21511.1
R32 VSS.n4560 VSS.n4559 21511.1
R33 VSS.n4764 VSS.n4763 21511.1
R34 VSS.n10187 VSS.n4555 21511.1
R35 VSS.n5169 VSS.n5168 21511.1
R36 VSS.n5092 VSS.n5091 21511.1
R37 VSS.n10362 VSS.n10281 21511.1
R38 VSS.n12493 VSS.n3599 21511.1
R39 VSS.n10358 VSS.n10282 21511.1
R40 VSS.n10511 VSS.n10254 21511.1
R41 VSS.n10517 VSS.n10252 21511.1
R42 VSS.n10241 VSS.n10240 21511.1
R43 VSS.n10247 VSS.n10246 21511.1
R44 VSS.n10250 VSS.n10249 21511.1
R45 VSS.n10504 VSS.n10255 21511.1
R46 VSS.n10305 VSS.n3600 21511.1
R47 VSS.n12485 VSS.n12484 21511.1
R48 VSS.n12506 VSS.n12505 21511.1
R49 VSS.n10206 VSS.n10205 21511.1
R50 VSS.n11436 VSS.n11435 21511.1
R51 VSS.n11347 VSS.n3638 20274.5
R52 VSS.n10410 VSS.n10409 20235.8
R53 VSS.n5094 VSS.n5093 18464.3
R54 VSS.n4814 VSS.n4813 18464.3
R55 VSS.n5101 VSS.n5100 18464.3
R56 VSS.n10530 VSS.n10529 17458.2
R57 VSS.n10506 VSS.n10505 17451.5
R58 VSS.n10510 VSS.n10509 17451.5
R59 VSS.n10522 VSS.n10521 17451.5
R60 VSS.n10516 VSS.n10515 17451.5
R61 VSS.n4896 VSS.n4889 17285.7
R62 VSS.n4866 VSS.n4865 17285.7
R63 VSS.n4880 VSS.n4879 17285.7
R64 VSS.n4557 VSS.n4556 17285.7
R65 VSS.n4855 VSS.n4854 17285.7
R66 VSS.n5060 VSS.n5059 17285.7
R67 VSS.n5065 VSS.n5064 17285.7
R68 VSS.n5174 VSS.n5173 17285.7
R69 VSS.n4843 VSS.n4777 17285.7
R70 VSS.n5051 VSS.n5050 17285.7
R71 VSS.n5039 VSS.n5037 17285.7
R72 VSS.n5164 VSS.n4728 17285.7
R73 VSS.n5162 VSS.n4730 17285.7
R74 VSS.n4837 VSS.n4836 17285.7
R75 VSS.n5030 VSS.n5029 17285.7
R76 VSS.n4993 VSS.n4992 17285.7
R77 VSS.n4998 VSS.n4996 17285.7
R78 VSS.n5150 VSS.n4733 17285.7
R79 VSS.n4825 VSS.n4785 17285.7
R80 VSS.n5020 VSS.n5019 17285.7
R81 VSS.n5009 VSS.n4976 17285.7
R82 VSS.n5007 VSS.n5006 17285.7
R83 VSS.n5143 VSS.n4736 17285.7
R84 VSS.n4929 VSS.n4928 17285.7
R85 VSS.n4969 VSS.n4968 17285.7
R86 VSS.n4794 VSS.n4793 17285.7
R87 VSS.n4791 VSS.n4790 17285.7
R88 VSS.n5136 VSS.n5133 17285.7
R89 VSS.n4937 VSS.n4802 17285.7
R90 VSS.n4959 VSS.n4958 17285.7
R91 VSS.n5089 VSS.n4748 17285.7
R92 VSS.n5124 VSS.n4742 17285.7
R93 VSS.n5122 VSS.n4744 17285.7
R94 VSS.n10292 VSS.n10291 17285.7
R95 VSS.n10294 VSS.n10225 17285.7
R96 VSS.n10345 VSS.n10344 17285.7
R97 VSS.n12519 VSS.n3591 17285.7
R98 VSS.n10429 VSS.n10271 17285.7
R99 VSS.n10220 VSS.n10219 17285.7
R100 VSS.n10327 VSS.n10326 17285.7
R101 VSS.n10336 VSS.n10330 17285.7
R102 VSS.n10334 VSS.n10333 17285.7
R103 VSS.n10397 VSS.n10269 17285.7
R104 VSS.n10455 VSS.n10454 17285.7
R105 VSS.n10449 VSS.n10448 17285.7
R106 VSS.n10446 VSS.n3378 17285.7
R107 VSS.n12533 VSS.n12532 17285.7
R108 VSS.n10464 VSS.n10265 17285.7
R109 VSS.n10476 VSS.n10475 17285.7
R110 VSS.n10473 VSS.n10472 17285.7
R111 VSS.n12546 VSS.n12545 17285.7
R112 VSS.n10499 VSS.n10256 17285.7
R113 VSS.n10489 VSS.n10487 17285.7
R114 VSS.n10244 VSS.n10243 17285.7
R115 VSS.n10537 VSS.n10536 17285.7
R116 VSS.n10284 VSS.n10283 17285.7
R117 VSS.n10288 VSS.n10287 17285.7
R118 VSS.n12512 VSS.n12510 17285.7
R119 VSS.n10369 VSS.n10368 17285.7
R120 VSS.n11479 VSS.n3604 17283.5
R121 VSS.n10171 VSS.n3685 14040.1
R122 VSS.n10511 VSS.n10510 12405.6
R123 VSS.n10517 VSS.n10516 12405.6
R124 VSS.n10521 VSS.n10250 12405.6
R125 VSS.n10505 VSS.n10504 12405.6
R126 VSS.n4951 VSS.n4808 12320
R127 VSS.n5093 VSS.n5092 12320
R128 VSS.n5102 VSS.n5101 12320
R129 VSS.n10176 VSS.n4560 11061.4
R130 VSS.n4896 VSS.n4895 11000
R131 VSS.n4855 VSS.n4774 11000
R132 VSS.n5059 VSS.n4774 11000
R133 VSS.n4766 VSS.n4720 11000
R134 VSS.n5173 VSS.n4720 11000
R135 VSS.n5052 VSS.n4777 11000
R136 VSS.n5052 VSS.n5051 11000
R137 VSS.n5050 VSS.n5049 11000
R138 VSS.n5039 VSS.n5038 11000
R139 VSS.n5038 VSS.n4728 11000
R140 VSS.n5164 VSS.n5163 11000
R141 VSS.n5163 VSS.n5162 11000
R142 VSS.n4837 VSS.n4782 11000
R143 VSS.n5029 VSS.n4782 11000
R144 VSS.n5031 VSS.n5030 11000
R145 VSS.n4994 VSS.n4993 11000
R146 VSS.n4996 VSS.n4994 11000
R147 VSS.n4998 VSS.n4997 11000
R148 VSS.n4997 VSS.n4733 11000
R149 VSS.n5021 VSS.n4785 11000
R150 VSS.n5021 VSS.n5020 11000
R151 VSS.n5019 VSS.n5018 11000
R152 VSS.n5009 VSS.n5008 11000
R153 VSS.n5008 VSS.n5007 11000
R154 VSS.n5006 VSS.n5005 11000
R155 VSS.n5005 VSS.n4736 11000
R156 VSS.n4929 VSS.n4799 11000
R157 VSS.n4968 VSS.n4799 11000
R158 VSS.n4970 VSS.n4969 11000
R159 VSS.n4793 VSS.n4792 11000
R160 VSS.n4792 VSS.n4791 11000
R161 VSS.n4790 VSS.n4739 11000
R162 VSS.n5133 VSS.n4739 11000
R163 VSS.n4960 VSS.n4802 11000
R164 VSS.n4960 VSS.n4959 11000
R165 VSS.n4952 VSS.n4748 11000
R166 VSS.n5090 VSS.n5089 11000
R167 VSS.n5090 VSS.n4742 11000
R168 VSS.n5124 VSS.n5123 11000
R169 VSS.n5123 VSS.n5122 11000
R170 VSS.n10293 VSS.n10292 11000
R171 VSS.n10294 VSS.n10293 11000
R172 VSS.n10569 VSS.n10225 11000
R173 VSS.n10569 VSS.n10568 11000
R174 VSS.n10346 VSS.n10227 11000
R175 VSS.n10346 VSS.n10345 11000
R176 VSS.n10344 VSS.n10343 11000
R177 VSS.n10343 VSS.n3591 11000
R178 VSS.n10430 VSS.n10429 11000
R179 VSS.n10430 VSS.n10219 11000
R180 VSS.n10572 VSS.n10220 11000
R181 VSS.n10328 VSS.n10327 11000
R182 VSS.n10330 VSS.n10328 11000
R183 VSS.n10336 VSS.n10335 11000
R184 VSS.n10335 VSS.n10334 11000
R185 VSS.n10456 VSS.n10269 11000
R186 VSS.n10456 VSS.n10455 11000
R187 VSS.n10449 VSS.n10443 11000
R188 VSS.n10448 VSS.n10447 11000
R189 VSS.n10447 VSS.n10446 11000
R190 VSS.n12534 VSS.n3378 11000
R191 VSS.n12534 VSS.n12533 11000
R192 VSS.n10465 VSS.n10464 11000
R193 VSS.n10466 VSS.n10465 11000
R194 VSS.n10477 VSS.n10469 11000
R195 VSS.n10477 VSS.n10476 11000
R196 VSS.n10475 VSS.n10474 11000
R197 VSS.n10474 VSS.n10473 11000
R198 VSS.n10472 VSS.n3375 11000
R199 VSS.n12545 VSS.n3375 11000
R200 VSS.n10499 VSS.n10498 11000
R201 VSS.n10498 VSS.n10497 11000
R202 VSS.n10486 VSS.n10259 11000
R203 VSS.n10487 VSS.n10486 11000
R204 VSS.n10489 VSS.n10488 11000
R205 VSS.n10488 VSS.n10243 11000
R206 VSS.n10535 VSS.n10244 11000
R207 VSS.n10536 VSS.n10535 11000
R208 VSS.n10285 VSS.n10284 11000
R209 VSS.n10287 VSS.n10285 11000
R210 VSS.n10301 VSS.n10300 11000
R211 VSS.n10311 VSS.n10302 11000
R212 VSS.n10311 VSS.n10310 11000
R213 VSS.n10307 VSS.n3595 11000
R214 VSS.n12510 VSS.n3595 11000
R215 VSS.n10368 VSS.n10367 11000
R216 VSS.n10367 VSS.n10366 11000
R217 VSS.n10361 VSS.n10277 11000
R218 VSS.n10361 VSS.n10360 11000
R219 VSS.n12498 VSS.n12497 11000
R220 VSS.n12499 VSS.n12498 11000
R221 VSS.n12501 VSS.n3597 11000
R222 VSS.n12300 VSS.n3597 11000
R223 VSS.n10300 VSS.n10299 10951.1
R224 VSS.n10569 VSS.n10224 10951.1
R225 VSS.n10570 VSS.n10569 10951.1
R226 VSS.n10573 VSS.n10572 10951.1
R227 VSS.n10443 VSS.n10442 10951.1
R228 VSS.n10457 VSS.n10456 10951.1
R229 VSS.n10465 VSS.n10263 10951.1
R230 VSS.n10293 VSS.n10217 10951.1
R231 VSS.n10430 VSS.n10218 10951.1
R232 VSS.n10285 VSS.n10213 10951.1
R233 VSS.n10293 VSS.n10214 10951.1
R234 VSS.n10367 VSS.n10209 10951.1
R235 VSS.n10285 VSS.n10210 10951.1
R236 VSS.n10189 VSS.n10188 10951.1
R237 VSS.n11429 VSS.n3684 10951.1
R238 VSS.n4872 VSS.n4870 10951.1
R239 VSS.n4877 VSS.n4876 10951.1
R240 VSS.n4870 VSS.n4869 10951.1
R241 VSS.n4846 VSS.n4782 10951.1
R242 VSS.n5052 VSS.n4776 10951.1
R243 VSS.n5053 VSS.n5052 10951.1
R244 VSS.n5055 VSS.n4774 10951.1
R245 VSS.n4953 VSS.n4952 10951.1
R246 VSS.n4960 VSS.n4801 10951.1
R247 VSS.n4971 VSS.n4970 10951.1
R248 VSS.n4961 VSS.n4960 10951.1
R249 VSS.n4963 VSS.n4799 10951.1
R250 VSS.n4828 VSS.n4799 10951.1
R251 VSS.n5021 VSS.n4784 10951.1
R252 VSS.n5018 VSS.n5017 10951.1
R253 VSS.n5032 VSS.n5031 10951.1
R254 VSS.n5022 VSS.n5021 10951.1
R255 VSS.n5024 VSS.n4782 10951.1
R256 VSS.n4891 VSS.n4774 10951.1
R257 VSS.n4895 VSS.n4894 10951.1
R258 VSS.n5049 VSS.n5048 10951.1
R259 VSS.n4876 VSS.n4875 10951.1
R260 VSS.n10196 VSS.n4551 10951.1
R261 VSS.n4903 VSS.n4902 10951.1
R262 VSS.n4723 VSS.n4722 10951.1
R263 VSS.n4722 VSS.n4559 10951.1
R264 VSS.n4555 VSS.n4554 10951.1
R265 VSS.n10188 VSS.n10187 10951.1
R266 VSS.n5163 VSS.n4729 10951.1
R267 VSS.n4994 VSS.n4757 10951.1
R268 VSS.n5038 VSS.n4761 10951.1
R269 VSS.n5005 VSS.n5004 10951.1
R270 VSS.n4997 VSS.n4983 10951.1
R271 VSS.n4792 VSS.n4750 10951.1
R272 VSS.n5008 VSS.n4754 10951.1
R273 VSS.n5091 VSS.n5090 10951.1
R274 VSS.n5123 VSS.n4743 10951.1
R275 VSS.n5129 VSS.n4739 10951.1
R276 VSS.n10362 VSS.n10361 10951.1
R277 VSS.n12498 VSS.n3599 10951.1
R278 VSS.n10361 VSS.n10358 10951.1
R279 VSS.n10300 VSS.n10282 10951.1
R280 VSS.n10431 VSS.n10430 10951.1
R281 VSS.n10456 VSS.n10268 10951.1
R282 VSS.n10465 VSS.n10264 10951.1
R283 VSS.n10498 VSS.n10257 10951.1
R284 VSS.n10478 VSS.n10477 10951.1
R285 VSS.n10343 VSS.n10342 10951.1
R286 VSS.n10335 VSS.n10320 10951.1
R287 VSS.n10328 VSS.n10230 10951.1
R288 VSS.n10447 VSS.n10234 10951.1
R289 VSS.n12535 VSS.n12534 10951.1
R290 VSS.n12541 VSS.n3375 10951.1
R291 VSS.n10474 VSS.n10238 10951.1
R292 VSS.n10498 VSS.n10255 10951.1
R293 VSS.n12498 VSS.n3600 10951.1
R294 VSS.n10311 VSS.n10305 10951.1
R295 VSS.n10312 VSS.n10311 10951.1
R296 VSS.n10347 VSS.n10346 10951.1
R297 VSS.n12485 VSS.n3597 10951.1
R298 VSS.n12505 VSS.n3597 10951.1
R299 VSS.n10167 VSS.n10166 9232.14
R300 VSS.n5176 VSS.n5174 9232.14
R301 VSS.n5156 VSS.n4730 9232.14
R302 VSS.n5150 VSS.n5149 9232.14
R303 VSS.n5143 VSS.n5142 9232.14
R304 VSS.n5136 VSS.n5135 9232.14
R305 VSS.n5115 VSS.n4744 9232.14
R306 VSS.n12519 VSS.n12518 9232.14
R307 VSS.n10333 VSS.n10332 9232.14
R308 VSS.n12532 VSS.n12531 9232.14
R309 VSS.n12547 VSS.n12546 9232.14
R310 VSS.n10539 VSS.n10537 9232.14
R311 VSS.n12512 VSS.n12511 9232.14
R312 VSS.n12306 VSS.n12305 9232.14
R313 VSS VSS.n3687 7931.8
R314 VSS VSS 7754.79
R315 VSS VSS 7754.79
R316 VSS.n10174 VSS.n3685 6319.07
R317 VSS.n10175 VSS.n3685 6267.1
R318 VSS.n10371 VSS.n10204 6020.82
R319 VSS.n11445 VSS.n3678 6020.82
R320 VSS.n4819 VSS.n4811 4827.93
R321 VSS.n4822 VSS.n4821 4827.93
R322 VSS.n4926 VSS.n4925 4827.93
R323 VSS.n4923 VSS.n4922 4827.93
R324 VSS.n4920 VSS.n4919 4827.93
R325 VSS.n4917 VSS.n4916 4827.93
R326 VSS.n4914 VSS.n4913 4827.93
R327 VSS.n4911 VSS.n4910 4827.93
R328 VSS.n10377 VSS.n10376 4827.93
R329 VSS.n10382 VSS.n10381 4827.93
R330 VSS.n10388 VSS.n10386 4827.93
R331 VSS.n10393 VSS.n10272 4827.93
R332 VSS.n10396 VSS.n10395 4827.93
R333 VSS.n10402 VSS.n10401 4827.93
R334 VSS.n10405 VSS.n10404 4827.93
R335 VSS.n10409 VSS.n10408 4827.93
R336 VSS.n11480 VSS.n11479 4810.3
R337 VSS.n5115 VSS.n5114 4376.55
R338 VSS.n5116 VSS.n5115 4376.55
R339 VSS.n5135 VSS.n5134 4376.55
R340 VSS.n5135 VSS.n4737 4376.55
R341 VSS.n5142 VSS.n5141 4376.55
R342 VSS.n5142 VSS.n4734 4376.55
R343 VSS.n5149 VSS.n5148 4376.55
R344 VSS.n5149 VSS.n4731 4376.55
R345 VSS.n5156 VSS.n5155 4376.55
R346 VSS.n5157 VSS.n5156 4376.55
R347 VSS.n5176 VSS.n5175 4376.55
R348 VSS.n5177 VSS.n5176 4376.55
R349 VSS.n10166 VSS.n4561 4376.55
R350 VSS.n12305 VSS.n12303 4376.55
R351 VSS.n12305 VSS.n12304 4376.55
R352 VSS.n12511 VSS.n3592 4376.55
R353 VSS.n12518 VSS.n12517 4376.55
R354 VSS.n12518 VSS.n3589 4376.55
R355 VSS.n10332 VSS.n3588 4376.55
R356 VSS.n10332 VSS.n3586 4376.55
R357 VSS.n12531 VSS.n3380 4376.55
R358 VSS.n12531 VSS.n12530 4376.55
R359 VSS.n12548 VSS.n12547 4376.55
R360 VSS.n12547 VSS.n3320 4376.55
R361 VSS.n10540 VSS.n10539 4376.55
R362 VSS.n10539 VSS.n10538 4376.55
R363 VSS.n10527 VSS.n10525 3774.78
R364 VSS.n12482 VSS.n3603 3288.62
R365 VSS.n10599 VSS.n10598 3147.35
R366 VSS.n10597 VSS.n10596 3147.35
R367 VSS.n11440 VSS.n11439 3147.35
R368 VSS.n11442 VSS.n11441 3147.35
R369 VSS.n11448 VSS.n11447 3147.35
R370 VSS.n11486 VSS.n3638 3085.55
R371 VSS.n4820 VSS.n4819 3072.32
R372 VSS.n4821 VSS.n4820 3072.32
R373 VSS.n4823 VSS.n4822 3072.32
R374 VSS.n4926 VSS.n4823 3072.32
R375 VSS.n4925 VSS.n4924 3072.32
R376 VSS.n4924 VSS.n4923 3072.32
R377 VSS.n4922 VSS.n4921 3072.32
R378 VSS.n4921 VSS.n4920 3072.32
R379 VSS.n4919 VSS.n4918 3072.32
R380 VSS.n4918 VSS.n4917 3072.32
R381 VSS.n4916 VSS.n4915 3072.32
R382 VSS.n4915 VSS.n4914 3072.32
R383 VSS.n4913 VSS.n4912 3072.32
R384 VSS.n4912 VSS.n4911 3072.32
R385 VSS.n10377 VSS.n10276 3072.32
R386 VSS.n10381 VSS.n10276 3072.32
R387 VSS.n10382 VSS.n10274 3072.32
R388 VSS.n10386 VSS.n10274 3072.32
R389 VSS.n10388 VSS.n10387 3072.32
R390 VSS.n10387 VSS.n10272 3072.32
R391 VSS.n10394 VSS.n10393 3072.32
R392 VSS.n10395 VSS.n10394 3072.32
R393 VSS.n10400 VSS.n10396 3072.32
R394 VSS.n10401 VSS.n10400 3072.32
R395 VSS.n10403 VSS.n10402 3072.32
R396 VSS.n10404 VSS.n10403 3072.32
R397 VSS.n10407 VSS.n10405 3072.32
R398 VSS.n10408 VSS.n10407 3072.32
R399 VSS.n4545 VSS.n4544 3014.53
R400 VSS.n10176 VSS.n3685 2895.44
R401 VSS.n4910 VSS.n4909 2574.58
R402 VSS.n10372 VSS.n10371 1881.22
R403 VSS.n10599 VSS.n10204 1881.22
R404 VSS.n10598 VSS.n10597 1881.22
R405 VSS.n10596 VSS.n10595 1881.22
R406 VSS.n11439 VSS.n3680 1881.22
R407 VSS.n11441 VSS.n11440 1881.22
R408 VSS.n11442 VSS.n3678 1881.22
R409 VSS.n11448 VSS.n11445 1881.22
R410 VSS VSS.n11345 1694.25
R411 VSS VSS 1567.82
R412 VSS.n11446 VSS.n3677 1544.68
R413 VSS.n11275 VSS.n11274 1544.5
R414 VSS.n11261 VSS 1266.45
R415 VSS.n11453 VSS.n11452 1250.46
R416 VSS.n4735 VSS 1088
R417 VSS.n4732 VSS 1088
R418 VSS.n5180 VSS 1088
R419 VSS.n10163 VSS 1088
R420 VSS.n10173 VSS 1088
R421 VSS.n12479 VSS 1088
R422 VSS.n3590 VSS 1088
R423 VSS.n14486 VSS 1088
R424 VSS.n12552 VSS 1088
R425 VSS.n3374 VSS 1088
R426 VSS.n11447 VSS.n11446 1073.06
R427 VSS.n11452 VSS.n3603 1043.16
R428 VSS.n3677 VSS.n3603 918.338
R429 VSS VSS.n11260 881.011
R430 VSS.n13603 VSS.n13485 880.317
R431 VSS.n14016 VSS.n1720 880.317
R432 VSS.n12796 VSS.n2935 880.317
R433 VSS.n10891 VSS.n3898 880.317
R434 VSS.n10987 VSS.n3859 880.317
R435 VSS.n11042 VSS.n3830 880.317
R436 VSS.n9577 VSS.n7555 880.317
R437 VSS.n8826 VSS.n8183 880.317
R438 VSS.n8788 VSS.n8215 880.317
R439 VSS.n6761 VSS.n6230 880.317
R440 VSS.n8114 VSS.n8034 880.317
R441 VSS.n8893 VSS.n7953 880.317
R442 VSS.n9516 VSS.n9016 880.317
R443 VSS.n9838 VSS.n7180 880.317
R444 VSS.n7367 VSS.n7208 880.317
R445 VSS.n9265 VSS.n9165 880.317
R446 VSS.n8958 VSS.n7814 880.317
R447 VSS.n8985 VSS.n7631 880.317
R448 VSS.n7775 VSS.n7666 880.317
R449 VSS.n7137 VSS.n7087 880.317
R450 VSS.n8932 VSS.n7877 880.317
R451 VSS.n6854 VSS.n6626 880.317
R452 VSS.n6921 VSS.n6578 880.317
R453 VSS.n7040 VSS.n6516 880.317
R454 VSS.n7053 VSS.n6289 880.317
R455 VSS.n6421 VSS.n6314 880.317
R456 VSS.n6786 VSS.n6674 880.317
R457 VSS.n10776 VSS.n4114 880.317
R458 VSS.n4405 VSS.n4404 880.317
R459 VSS.n4344 VSS.n4234 880.317
R460 VSS.n1165 VSS.n879 880.317
R461 VSS.n14229 VSS.n14228 880.317
R462 VSS.n1151 VSS.n602 880.317
R463 VSS.n13045 VSS.n2478 880.317
R464 VSS.n13101 VSS.n2356 880.317
R465 VSS.n2342 VSS.n1928 880.317
R466 VSS.n14115 VSS.n650 880.317
R467 VSS.n14079 VSS.n1661 880.317
R468 VSS.n13643 VSS.n13221 880.317
R469 VSS.n1435 VSS.n818 880.317
R470 VSS.n2245 VSS.n2005 880.317
R471 VSS.n2180 VSS.n2080 880.317
R472 VSS.n13188 VSS.n1849 880.317
R473 VSS.n13935 VSS.n1777 880.317
R474 VSS.n2319 VSS.n1972 880.317
R475 VSS.n12985 VSS.n2584 880.317
R476 VSS.n12949 VSS.n2688 880.317
R477 VSS.n12908 VSS.n2765 880.317
R478 VSS.n12872 VSS.n2868 880.317
R479 VSS.n12730 VSS.n2955 880.317
R480 VSS.n13024 VSS.n2524 880.317
R481 VSS.n4909 VSS.n4908 851.542
R482 VSS.n13583 VSS.n13484 754.287
R483 VSS.n1764 VSS.n1719 754.287
R484 VSS.n12781 VSS.n12780 754.287
R485 VSS.n10876 VSS.n10875 754.287
R486 VSS.n10947 VSS.n10946 754.287
R487 VSS.n11027 VSS.n11026 754.287
R488 VSS.n8279 VSS.n7569 754.287
R489 VSS.n8822 VSS.n8184 754.287
R490 VSS.n8383 VSS.n8188 754.287
R491 VSS.n8784 VSS.n8216 754.287
R492 VSS.n8779 VSS.n8777 754.287
R493 VSS.n6744 VSS.n6743 754.287
R494 VSS.n8151 VSS.n8150 754.287
R495 VSS.n8041 VSS.n8038 754.287
R496 VSS.n8876 VSS.n8875 754.287
R497 VSS.n9289 VSS.n9017 754.287
R498 VSS.n7182 VSS.n7181 754.287
R499 VSS.n7266 VSS.n7263 754.287
R500 VSS.n9213 VSS.n9212 754.287
R501 VSS.n7909 VSS.n7852 754.287
R502 VSS.n7638 VSS.n7637 754.287
R503 VSS.n7673 VSS.n7672 754.287
R504 VSS.n7093 VSS.n7090 754.287
R505 VSS.n7993 VSS.n7942 754.287
R506 VSS.n6633 VSS.n6630 754.287
R507 VSS.n6585 VSS.n6582 754.287
R508 VSS.n6944 VSS.n6541 754.287
R509 VSS.n6487 VSS.n6484 754.287
R510 VSS.n6320 VSS.n6317 754.287
R511 VSS.n6684 VSS.n6677 754.287
R512 VSS.n4453 VSS.n4452 754.287
R513 VSS.n4378 VSS.n4165 754.287
R514 VSS.n4267 VSS.n4233 754.287
R515 VSS.n886 VSS.n883 754.287
R516 VSS.n14201 VSS.n14200 754.287
R517 VSS.n2399 VSS.n549 754.287
R518 VSS.n1134 VSS.n1133 754.287
R519 VSS.n2486 VSS.n2483 754.287
R520 VSS.n2453 VSS.n2452 754.287
R521 VSS.n13093 VSS.n2372 754.287
R522 VSS.n1934 VSS.n1931 754.287
R523 VSS.n1459 VSS.n651 754.287
R524 VSS.n1668 VSS.n1667 754.287
R525 VSS.n13227 VSS.n13224 754.287
R526 VSS.n1190 VSS.n842 754.287
R527 VSS.n2008 VSS.n2006 754.287
R528 VSS.n2083 VSS.n2081 754.287
R529 VSS.n1857 VSS.n1854 754.287
R530 VSS.n13927 VSS.n1793 754.287
R531 VSS.n1975 VSS.n1967 754.287
R532 VSS.n2587 VSS.n2585 754.287
R533 VSS.n2695 VSS.n2694 754.287
R534 VSS.n2768 VSS.n2766 754.287
R535 VSS.n2875 VSS.n2874 754.287
R536 VSS.n12722 VSS.n2971 754.287
R537 VSS.n2527 VSS.n2519 754.287
R538 VSS.n13584 VSS.n13502 750
R539 VSS.n1765 VSS.n1737 750
R540 VSS.n12785 VSS.n12783 750
R541 VSS.n10880 VSS.n10878 750
R542 VSS.n10944 VSS.n10943 750
R543 VSS.n11031 VSS.n11029 750
R544 VSS.n9555 VSS.n9554 750
R545 VSS.n8817 VSS.n8816 750
R546 VSS.n8243 VSS.n8242 750
R547 VSS.n6741 VSS.n6711 750
R548 VSS.n8116 VSS.n8115 750
R549 VSS.n8873 VSS.n7968 750
R550 VSS.n9515 VSS.n9513 750
R551 VSS.n9837 VSS.n9835 750
R552 VSS.n7369 VSS.n7368 750
R553 VSS.n9241 VSS.n9240 750
R554 VSS.n8948 VSS.n8947 750
R555 VSS.n8984 VSS.n7632 750
R556 VSS.n7774 VSS.n7667 750
R557 VSS.n7139 VSS.n7138 750
R558 VSS.n8923 VSS.n8922 750
R559 VSS.n6856 VSS.n6855 750
R560 VSS.n6923 VSS.n6922 750
R561 VSS.n6996 VSS.n6995 750
R562 VSS.n7055 VSS.n7054 750
R563 VSS.n6423 VSS.n6422 750
R564 VSS.n6788 VSS.n6787 750
R565 VSS.n4450 VSS.n4449 750
R566 VSS.n4380 VSS.n4379 750
R567 VSS.n4268 VSS.n4251 750
R568 VSS.n1167 VSS.n1166 750
R569 VSS.n2402 VSS.n2401 750
R570 VSS.n1131 VSS.n929 750
R571 VSS.n13047 VSS.n13046 750
R572 VSS.n13094 VSS.n2363 750
R573 VSS.n2344 VSS.n2343 750
R574 VSS.n14114 VSS.n14112 750
R575 VSS.n14078 VSS.n1662 750
R576 VSS.n13645 VSS.n13644 750
R577 VSS.n1411 VSS.n1410 750
R578 VSS.n2244 VSS.n2242 750
R579 VSS.n2179 VSS.n2177 750
R580 VSS.n13190 VSS.n13189 750
R581 VSS.n13928 VSS.n1784 750
R582 VSS.n2318 VSS.n1973 750
R583 VSS.n12984 VSS.n12982 750
R584 VSS.n12948 VSS.n2689 750
R585 VSS.n12907 VSS.n12905 750
R586 VSS.n12871 VSS.n2869 750
R587 VSS.n12723 VSS.n2962 750
R588 VSS.n13023 VSS.n2525 750
R589 VSS.n4864 VSS.n4546 745.378
R590 VSS.n10199 VSS.n10198 745.378
R591 VSS.n3683 VSS.n3682 745.378
R592 VSS VSS 733.333
R593 VSS.n11348 VSS.n11347 708.047
R594 VSS VSS.n4735 688
R595 VSS VSS.n4732 688
R596 VSS.n5180 VSS 688
R597 VSS VSS.n10163 688
R598 VSS VSS.n10173 688
R599 VSS VSS.n3590 688
R600 VSS.n12549 VSS.n3374 673.318
R601 VSS.n14487 VSS.n14486 656.076
R602 VSS.n12552 VSS.n3319 656.076
R603 VSS.n12479 VSS.n3605 656
R604 VSS.n11348 VSS 632.184
R605 VSS.n11345 VSS 623.755
R606 VSS.n11276 VSS.n11275 617.899
R607 VSS.n11487 VSS.n11486 617.899
R608 VSS.n11349 VSS.n11348 613.249
R609 VSS.n11345 VSS.n3695 613.249
R610 VSS.n11486 VSS.n3639 613.249
R611 VSS VSS.n11485 460.231
R612 VSS.n10527 VSS.n10526 445.471
R613 VSS.n11446 VSS.n3602 435.765
R614 VSS.n11309 VSS.n11308 433.748
R615 VSS.n4902 VSS.n4547 389.642
R616 VSS.n4901 VSS.n4548 389.642
R617 VSS.n10197 VSS.n10196 389.642
R618 VSS.n10195 VSS.n10194 389.642
R619 VSS.n11430 VSS.n11429 389.642
R620 VSS.n11413 VSS.n3687 306.625
R621 VSS.n4817 VSS.n4816 274.635
R622 VSS.n10375 VSS.n10374 274.635
R623 VSS.n10631 VSS.n4543 257.318
R624 VSS.n10603 VSS.n10200 257.318
R625 VSS.n10420 VSS.n10418 257.318
R626 VSS.n4860 VSS.n4859 257.318
R627 VSS.n4933 VSS.n4927 257.318
R628 VSS.n4949 VSS.n4948 257.318
R629 VSS.n5098 VSS.n5096 257.318
R630 VSS.n4943 VSS.n4942 257.318
R631 VSS.n4936 VSS.n4935 257.318
R632 VSS.n4834 VSS.n4833 257.318
R633 VSS.n4841 VSS.n4840 257.318
R634 VSS.n4852 VSS.n4851 257.318
R635 VSS.n4887 VSS.n4862 257.318
R636 VSS.n4907 VSS 257.318
R637 VSS VSS.n4905 257.318
R638 VSS.n10193 VSS 257.318
R639 VSS VSS.n4552 257.318
R640 VSS VSS.n10175 257.318
R641 VSS.n5106 VSS.n5105 257.318
R642 VSS.n12489 VSS.n12483 257.318
R643 VSS.n10391 VSS.n10390 257.318
R644 VSS.n10385 VSS.n10384 257.318
R645 VSS.n10380 VSS.n10379 257.318
R646 VSS.n10594 VSS.n10592 257.318
R647 VSS.n11443 VSS.n3679 257.318
R648 VSS.n12492 VSS.n12491 257.318
R649 VSS.n10426 VSS.n10425 257.318
R650 VSS.n10423 VSS.n10422 257.318
R651 VSS.n10416 VSS.n10415 257.318
R652 VSS VSS.n10413 257.318
R653 VSS.n10507 VSS 257.318
R654 VSS.n10513 VSS 257.318
R655 VSS.n10519 VSS 257.318
R656 VSS VSS.n10532 257.318
R657 VSS.n11433 VSS.n11432 257.318
R658 VSS.n11451 VSS 257.318
R659 VSS VSS.n3681 257.318
R660 VSS VSS.n10203 257.318
R661 VSS.n10630 VSS.n10605 257.318
R662 VSS.n5110 VSS 240.076
R663 VSS VSS.n5119 240.076
R664 VSS.n5138 VSS 240.076
R665 VSS.n5145 VSS 240.076
R666 VSS.n5152 VSS 240.076
R667 VSS VSS.n5159 240.076
R668 VSS VSS.n5179 240.076
R669 VSS.n10169 VSS 240.076
R670 VSS.n12308 VSS 240.076
R671 VSS.n12514 VSS 240.076
R672 VSS.n12525 VSS 240.076
R673 VSS.n12521 VSS 240.076
R674 VSS.n11433 VSS 240
R675 VSS.n10549 VSS.n10242 240
R676 VSS.n10481 VSS.n10480 240
R677 VSS VSS.n10416 240
R678 VSS.n12508 VSS.n3596 240
R679 VSS.n5126 VSS.n4741 240
R680 VSS.n5087 VSS.n5085 240
R681 VSS.n5131 VSS.n4740 240
R682 VSS.n10181 VSS.n4558 240
R683 VSS.n10185 VSS.n4553 240
R684 VSS.n5046 VSS.n5042 240
R685 VSS.n5074 VSS.n4758 240
R686 VSS.n5082 VSS.n4751 240
R687 VSS.n4887 VSS 240
R688 VSS.n4833 VSS 240
R689 VSS.n4942 VSS 240
R690 VSS.n4936 VSS 240
R691 VSS.n5105 VSS 240
R692 VSS.n5096 VSS 240
R693 VSS VSS.n4810 240
R694 VSS.n4949 VSS 240
R695 VSS VSS 240
R696 VSS VSS.n4956 240
R697 VSS VSS.n5085 240
R698 VSS.n4956 VSS.n4806 240
R699 VSS VSS.n4806 240
R700 VSS VSS.n4800 240
R701 VSS VSS.n4933 240
R702 VSS VSS.n4826 240
R703 VSS.n4827 VSS 240
R704 VSS.n4965 VSS 240
R705 VSS.n4973 VSS.n4797 240
R706 VSS VSS.n5012 240
R707 VSS.n4973 VSS 240
R708 VSS VSS.n4797 240
R709 VSS VSS.n5082 240
R710 VSS VSS.n5078 240
R711 VSS.n5002 VSS.n4981 240
R712 VSS.n4989 VSS.n4985 240
R713 VSS VSS.n4985 240
R714 VSS VSS.n5002 240
R715 VSS.n5078 VSS.n5077 240
R716 VSS.n5077 VSS 240
R717 VSS.n5015 VSS.n5012 240
R718 VSS VSS.n5015 240
R719 VSS VSS.n4783 240
R720 VSS.n4840 VSS 240
R721 VSS.n4851 VSS 240
R722 VSS VSS.n4775 240
R723 VSS.n4859 VSS 240
R724 VSS.n4890 VSS 240
R725 VSS VSS.n4886 240
R726 VSS.n5057 VSS 240
R727 VSS VSS.n4844 240
R728 VSS.n4845 VSS 240
R729 VSS.n5026 VSS 240
R730 VSS.n5034 VSS.n4780 240
R731 VSS.n5034 VSS 240
R732 VSS VSS 240
R733 VSS VSS.n4780 240
R734 VSS VSS.n5074 240
R735 VSS VSS.n5070 240
R736 VSS.n5166 VSS.n4727 240
R737 VSS.n5171 VSS.n4726 240
R738 VSS.n5171 VSS 240
R739 VSS.n5166 VSS 240
R740 VSS.n5070 VSS.n5069 240
R741 VSS.n5069 VSS 240
R742 VSS VSS.n5042 240
R743 VSS VSS.n5046 240
R744 VSS.n5062 VSS.n4772 240
R745 VSS.n4771 VSS.n4769 240
R746 VSS VSS.n4771 240
R747 VSS.n5062 VSS 240
R748 VSS VSS.n4772 240
R749 VSS VSS 240
R750 VSS VSS.n4883 240
R751 VSS.n4883 VSS.n4867 240
R752 VSS VSS.n4867 240
R753 VSS.n4898 VSS.n4886 240
R754 VSS.n4898 VSS 240
R755 VSS VSS.n4553 240
R756 VSS VSS.n10185 240
R757 VSS VSS.n10181 240
R758 VSS.n4558 VSS 240
R759 VSS VSS.n4726 240
R760 VSS VSS.n4769 240
R761 VSS VSS.n4727 240
R762 VSS VSS.n4989 240
R763 VSS VSS.n4758 240
R764 VSS VSS.n4981 240
R765 VSS VSS.n4740 240
R766 VSS VSS.n4751 240
R767 VSS.n5131 VSS 240
R768 VSS.n5126 VSS 240
R769 VSS VSS.n5087 240
R770 VSS VSS.n4741 240
R771 VSS VSS.n5113 240
R772 VSS VSS.n4738 240
R773 VSS.n10426 VSS 240
R774 VSS.n10390 VSS 240
R775 VSS.n10384 VSS 240
R776 VSS.n10379 VSS 240
R777 VSS.n10592 VSS 240
R778 VSS VSS.n3679 240
R779 VSS VSS.n10279 240
R780 VSS.n12492 VSS 240
R781 VSS VSS.n3598 240
R782 VSS VSS.n12489 240
R783 VSS.n12299 VSS 240
R784 VSS VSS.n3594 240
R785 VSS VSS.n3605 240
R786 VSS VSS.n12480 240
R787 VSS.n12508 VSS 240
R788 VSS.n12503 VSS 240
R789 VSS VSS.n3601 240
R790 VSS VSS.n10278 240
R791 VSS VSS.n10207 240
R792 VSS VSS.n10589 240
R793 VSS VSS.n10211 240
R794 VSS VSS.n10585 240
R795 VSS VSS.n10223 240
R796 VSS VSS 240
R797 VSS VSS.n10215 240
R798 VSS VSS.n10581 240
R799 VSS VSS.n10577 240
R800 VSS VSS.n10221 240
R801 VSS.n10270 VSS 240
R802 VSS VSS.n10423 240
R803 VSS VSS.n10420 240
R804 VSS VSS.n10462 240
R805 VSS.n10258 VSS 240
R806 VSS VSS.n10262 240
R807 VSS VSS.n10267 240
R808 VSS.n10434 VSS 240
R809 VSS VSS.n10452 240
R810 VSS.n10452 VSS.n10451 240
R811 VSS.n10451 VSS 240
R812 VSS.n10222 VSS.n10221 240
R813 VSS VSS.n10222 240
R814 VSS VSS.n10226 240
R815 VSS.n10290 VSS 240
R816 VSS VSS.n10355 240
R817 VSS VSS.n10351 240
R818 VSS.n10565 VSS.n10228 240
R819 VSS.n10340 VSS.n10318 240
R820 VSS VSS.n10340 240
R821 VSS.n10228 VSS 240
R822 VSS VSS.n10565 240
R823 VSS.n10561 VSS.n10231 240
R824 VSS VSS.n10324 240
R825 VSS VSS 240
R826 VSS VSS.n10231 240
R827 VSS VSS.n10561 240
R828 VSS.n10557 VSS.n10235 240
R829 VSS.n12538 VSS 240
R830 VSS VSS.n10235 240
R831 VSS VSS.n10557 240
R832 VSS VSS.n10553 240
R833 VSS VSS.n3376 240
R834 VSS.n10553 VSS.n10552 240
R835 VSS.n10552 VSS 240
R836 VSS.n10480 VSS 240
R837 VSS VSS 240
R838 VSS.n10481 VSS 240
R839 VSS.n10494 VSS.n10492 240
R840 VSS.n10492 VSS 240
R841 VSS VSS.n10494 240
R842 VSS.n10242 VSS 240
R843 VSS VSS.n10549 240
R844 VSS VSS 240
R845 VSS VSS.n10545 240
R846 VSS.n10545 VSS.n10544 240
R847 VSS.n10544 VSS 240
R848 VSS.n12543 VSS.n3376 240
R849 VSS.n12543 VSS 240
R850 VSS.n12538 VSS.n12537 240
R851 VSS.n12537 VSS 240
R852 VSS.n10324 VSS.n10321 240
R853 VSS VSS.n10321 240
R854 VSS.n10501 VSS 240
R855 VSS VSS 240
R856 VSS VSS.n20 240
R857 VSS VSS.n21 240
R858 VSS VSS.n10541 240
R859 VSS.n12551 VSS 240
R860 VSS.n12529 VSS 240
R861 VSS VSS.n12528 240
R862 VSS VSS.n12524 240
R863 VSS VSS.n10318 240
R864 VSS VSS.n3596 240
R865 VSS.n10306 VSS 240
R866 VSS VSS.n10603 240
R867 VSS.n8782 VSS.n8781 236.089
R868 VSS.n6740 VSS.n6231 236.089
R869 VSS.n8148 VSS.n8118 236.089
R870 VSS.n8872 VSS.n8871 236.089
R871 VSS.n8820 VSS.n8819 236.089
R872 VSS.n9559 VSS.n9557 236.089
R873 VSS.n9511 VSS.n9510 236.089
R874 VSS.n9833 VSS.n9832 236.089
R875 VSS.n7372 VSS.n7371 236.089
R876 VSS.n9245 VSS.n9243 236.089
R877 VSS.n8952 VSS.n8950 236.089
R878 VSS.n7806 VSS.n7805 236.089
R879 VSS.n7727 VSS.n7726 236.089
R880 VSS.n7142 VSS.n7141 236.089
R881 VSS.n8926 VSS.n8925 236.089
R882 VSS.n6904 VSS.n6858 236.089
R883 VSS.n6977 VSS.n6925 236.089
R884 VSS.n7000 VSS.n6998 236.089
R885 VSS.n7058 VSS.n7057 236.089
R886 VSS.n6426 VSS.n6425 236.089
R887 VSS.n6791 VSS.n6790 236.089
R888 VSS.n6394 VSS.n3838 236.089
R889 VSS.n10919 VSS.n3880 236.089
R890 VSS.n7340 VSS.n3906 236.089
R891 VSS.n4271 VSS.n4270 236.089
R892 VSS.n4383 VSS.n4382 236.089
R893 VSS.n10772 VSS.n10771 236.089
R894 VSS.n14198 VSS.n604 236.089
R895 VSS.n13050 VSS.n13049 236.089
R896 VSS.n13096 VSS.n13092 236.089
R897 VSS.n2347 VSS.n2346 236.089
R898 VSS.n2398 VSS.n582 236.089
R899 VSS.n1392 VSS.n1169 236.089
R900 VSS.n14110 VSS.n14109 236.089
R901 VSS.n13695 VSS.n1670 236.089
R902 VSS.n13648 VSS.n13647 236.089
R903 VSS.n1415 VSS.n1413 236.089
R904 VSS.n2240 VSS.n2239 236.089
R905 VSS.n2175 VSS.n2174 236.089
R906 VSS.n13193 VSS.n13192 236.089
R907 VSS.n13930 VSS.n13926 236.089
R908 VSS.n2278 VSS.n2277 236.089
R909 VSS.n12980 VSS.n12979 236.089
R910 VSS.n2812 VSS.n2697 236.089
R911 VSS.n12903 VSS.n12902 236.089
R912 VSS.n12636 VSS.n2877 236.089
R913 VSS.n12725 VSS.n12721 236.089
R914 VSS.n2632 VSS.n2529 236.089
R915 VSS.n12760 VSS.n12759 236.089
R916 VSS.n1768 VSS.n1767 236.089
R917 VSS.n13586 VSS.n13582 236.089
R918 VSS.n4908 VSS.n4546 232.895
R919 VSS.n4864 VSS.n4547 232.895
R920 VSS.n4902 VSS.n4901 232.895
R921 VSS.n10199 VSS.n4548 232.895
R922 VSS.n10198 VSS.n10197 232.895
R923 VSS.n10196 VSS.n10195 232.895
R924 VSS.n10194 VSS.n3682 232.895
R925 VSS.n11430 VSS.n3683 232.895
R926 VSS.n10600 VSS 225.319
R927 VSS.n4550 VSS 225.319
R928 VSS VSS.n10417 225.319
R929 VSS.n4861 VSS 225.319
R930 VSS.n4824 VSS 225.319
R931 VSS VSS.n4815 225.319
R932 VSS.n4818 VSS 225.319
R933 VSS.n5099 VSS 225.319
R934 VSS.n5095 VSS 225.319
R935 VSS.n4946 VSS 225.319
R936 VSS VSS.n4934 225.319
R937 VSS.n4835 VSS 225.319
R938 VSS.n4842 VSS 225.319
R939 VSS.n4853 VSS 225.319
R940 VSS.n4863 VSS 225.319
R941 VSS VSS.n4906 225.319
R942 VSS VSS.n4549 225.319
R943 VSS VSS.n10192 225.319
R944 VSS.n10177 VSS 225.319
R945 VSS.n5109 VSS 225.319
R946 VSS.n5154 VSS.n5153 225.319
R947 VSS VSS.n10174 225.319
R948 VSS.n10392 VSS 225.319
R949 VSS.n10389 VSS 225.319
R950 VSS.n10383 VSS 225.319
R951 VSS.n10378 VSS 225.319
R952 VSS VSS.n10373 225.319
R953 VSS VSS.n10593 225.319
R954 VSS.n11444 VSS 225.319
R955 VSS VSS.n12490 225.319
R956 VSS.n12481 VSS 225.319
R957 VSS VSS.n10424 225.319
R958 VSS VSS.n10421 225.319
R959 VSS VSS.n10414 225.319
R960 VSS VSS.n10412 225.319
R961 VSS.n10508 VSS 225.319
R962 VSS.n10514 VSS 225.319
R963 VSS.n10523 VSS 225.319
R964 VSS VSS.n10531 225.319
R965 VSS VSS.n11431 225.319
R966 VSS VSS.n11450 225.319
R967 VSS.n11449 VSS 225.319
R968 VSS.n11438 VSS 225.319
R969 VSS VSS.n10604 225.319
R970 VSS.n5112 VSS.n5111 208.076
R971 VSS.n5118 VSS.n5117 208.076
R972 VSS.n12298 VSS.n12297 208.076
R973 VSS.n12527 VSS.n12526 208.076
R974 VSS.n12523 VSS.n12522 208.076
R975 VSS VSS.n4807 208
R976 VSS VSS.n4807 208
R977 VSS VSS.n4931 208
R978 VSS VSS.n4931 208
R979 VSS VSS.n4966 208
R980 VSS VSS.n4966 208
R981 VSS VSS.n4795 208
R982 VSS VSS.n4795 208
R983 VSS VSS.n5080 208
R984 VSS VSS.n5080 208
R985 VSS VSS.n4857 208
R986 VSS VSS.n4857 208
R987 VSS VSS.n5027 208
R988 VSS VSS.n5027 208
R989 VSS VSS.n4990 208
R990 VSS VSS.n4990 208
R991 VSS VSS.n5072 208
R992 VSS VSS.n5072 208
R993 VSS VSS.n5044 208
R994 VSS VSS.n5044 208
R995 VSS VSS.n4868 208
R996 VSS VSS.n4868 208
R997 VSS VSS.n10183 208
R998 VSS VSS.n10183 208
R999 VSS VSS.n10179 208
R1000 VSS VSS.n10179 208
R1001 VSS.n5140 VSS.n5139 208
R1002 VSS.n5147 VSS.n5146 208
R1003 VSS.n5158 VSS.n4718 208
R1004 VSS.n5178 VSS.n4563 208
R1005 VSS.n10172 VSS.n10170 208
R1006 VSS VSS.n12487 208
R1007 VSS VSS.n12487 208
R1008 VSS.n12302 VSS 208
R1009 VSS.n12302 VSS 208
R1010 VSS.n12516 VSS.n12515 208
R1011 VSS VSS.n10587 208
R1012 VSS VSS.n10587 208
R1013 VSS VSS.n10583 208
R1014 VSS VSS.n10583 208
R1015 VSS VSS.n10579 208
R1016 VSS VSS.n10579 208
R1017 VSS VSS.n10266 208
R1018 VSS VSS.n10266 208
R1019 VSS.n10436 VSS 208
R1020 VSS.n10436 VSS 208
R1021 VSS VSS.n10353 208
R1022 VSS VSS.n10353 208
R1023 VSS VSS.n10349 208
R1024 VSS VSS.n10349 208
R1025 VSS VSS.n10563 208
R1026 VSS VSS.n10563 208
R1027 VSS VSS.n10559 208
R1028 VSS VSS.n10559 208
R1029 VSS VSS.n10555 208
R1030 VSS VSS.n10555 208
R1031 VSS VSS.n10260 208
R1032 VSS VSS.n10260 208
R1033 VSS VSS.n10547 208
R1034 VSS VSS.n10547 208
R1035 VSS.n10631 VSS.n10630 208
R1036 VSS.n11498 VSS.n11497 203.197
R1037 VSS.n11486 VSS 183.333
R1038 VSS.n11428 VSS.n11427 169.403
R1039 VSS.n11311 VSS.n11310 140.675
R1040 VSS.n11428 VSS.n3685 137.083
R1041 VSS.n11429 VSS.n11428 132.845
R1042 VSS.n4747 VSS 112.659
R1043 VSS VSS.n4940 112.659
R1044 VSS.n5088 VSS 112.659
R1045 VSS.n4972 VSS 112.659
R1046 VSS.n4957 VSS 112.659
R1047 VSS.n4964 VSS 112.659
R1048 VSS.n4939 VSS 112.659
R1049 VSS.n4830 VSS 112.659
R1050 VSS.n5016 VSS 112.659
R1051 VSS.n5151 VSS 112.659
R1052 VSS VSS.n5000 112.659
R1053 VSS.n4977 VSS 112.659
R1054 VSS VSS.n5075 112.659
R1055 VSS VSS.n5010 112.659
R1056 VSS.n5033 VSS 112.659
R1057 VSS.n4787 VSS 112.659
R1058 VSS.n5025 VSS 112.659
R1059 VSS VSS.n4831 112.659
R1060 VSS VSS.n4838 112.659
R1061 VSS VSS.n4849 112.659
R1062 VSS.n4893 VSS 112.659
R1063 VSS.n5061 VSS 112.659
R1064 VSS.n5056 VSS 112.659
R1065 VSS.n4779 VSS 112.659
R1066 VSS.n4848 VSS 112.659
R1067 VSS.n5047 VSS 112.659
R1068 VSS VSS.n4719 112.659
R1069 VSS.n5170 VSS 112.659
R1070 VSS.n5165 VSS 112.659
R1071 VSS VSS.n5067 112.659
R1072 VSS VSS.n5040 112.659
R1073 VSS.n10186 VSS 112.659
R1074 VSS.n5066 VSS 112.659
R1075 VSS VSS.n4881 112.659
R1076 VSS VSS.n4873 112.659
R1077 VSS VSS.n4884 112.659
R1078 VSS.n4904 VSS 112.659
R1079 VSS.n4897 VSS 112.659
R1080 VSS.n10191 VSS 112.659
R1081 VSS.n10168 VSS 112.659
R1082 VSS VSS.n4724 112.659
R1083 VSS VSS.n4767 112.659
R1084 VSS VSS.n5160 112.659
R1085 VSS VSS.n4987 112.659
R1086 VSS.n4999 VSS 112.659
R1087 VSS.n5144 VSS 112.659
R1088 VSS.n5003 VSS 112.659
R1089 VSS.n4789 VSS 112.659
R1090 VSS VSS.n5083 112.659
R1091 VSS.n5137 VSS 112.659
R1092 VSS.n5130 VSS 112.659
R1093 VSS.n5125 VSS 112.659
R1094 VSS VSS.n5120 112.659
R1095 VSS VSS.n5103 112.659
R1096 VSS VSS.n10216 112.659
R1097 VSS VSS.n10212 112.659
R1098 VSS VSS.n10208 112.659
R1099 VSS VSS.n10590 112.659
R1100 VSS.n10363 VSS 112.659
R1101 VSS.n12495 VSS 112.659
R1102 VSS.n12513 VSS 112.659
R1103 VSS.n12507 VSS 112.659
R1104 VSS.n12502 VSS 112.659
R1105 VSS.n10304 VSS 112.659
R1106 VSS.n12496 VSS 112.659
R1107 VSS VSS.n10356 112.659
R1108 VSS VSS.n10364 112.659
R1109 VSS.n10289 VSS 112.659
R1110 VSS.n10296 VSS 112.659
R1111 VSS VSS.n10575 112.659
R1112 VSS.n10433 VSS 112.659
R1113 VSS.n10428 VSS 112.659
R1114 VSS VSS.n10398 112.659
R1115 VSS VSS.n10495 112.659
R1116 VSS VSS.n10460 112.659
R1117 VSS.n10468 VSS 112.659
R1118 VSS.n10459 VSS 112.659
R1119 VSS.n10479 VSS 112.659
R1120 VSS VSS.n10236 112.659
R1121 VSS.n10441 VSS 112.659
R1122 VSS VSS.n10232 112.659
R1123 VSS.n10574 VSS 112.659
R1124 VSS VSS.n10566 112.659
R1125 VSS VSS.n10297 112.659
R1126 VSS VSS.n10338 112.659
R1127 VSS.n10314 VSS 112.659
R1128 VSS.n10337 VSS 112.659
R1129 VSS VSS.n10444 112.659
R1130 VSS.n10471 VSS 112.659
R1131 VSS VSS.n10550 112.659
R1132 VSS.n10470 VSS 112.659
R1133 VSS VSS.n10490 112.659
R1134 VSS.n10512 VSS 112.659
R1135 VSS.n10518 VSS 112.659
R1136 VSS VSS.n10533 112.659
R1137 VSS VSS.n10542 112.659
R1138 VSS.n10248 VSS 112.659
R1139 VSS VSS.n3321 112.659
R1140 VSS.n12542 VSS 112.659
R1141 VSS.n3379 VSS 112.659
R1142 VSS.n12536 VSS 112.659
R1143 VSS VSS.n3587 112.659
R1144 VSS.n10503 VSS 112.659
R1145 VSS.n10500 VSS 112.659
R1146 VSS.n12520 VSS 112.659
R1147 VSS.n10341 VSS 112.659
R1148 VSS VSS.n10308 112.659
R1149 VSS.n11437 VSS 112.659
R1150 VSS VSS.n10601 112.659
R1151 VSS.n3676 VSS.n3675 89.977
R1152 VSS.n11232 VSS.n11231 89.977
R1153 VSS.n13589 VSS.n13586 84.2672
R1154 VSS.n1767 VSS.n1763 84.2672
R1155 VSS.n12760 VSS.n2930 84.2672
R1156 VSS.n12902 VSS.n2842 84.2672
R1157 VSS.n2812 VSS.n2811 84.2672
R1158 VSS.n3906 VSS.n3893 84.2672
R1159 VSS.n10942 VSS.n10919 84.2672
R1160 VSS.n3838 VSS.n3825 84.2672
R1161 VSS.n6977 VSS.n6561 84.2672
R1162 VSS.n9562 VSS.n9559 84.2672
R1163 VSS.n8820 VSS.n8185 84.2672
R1164 VSS.n8782 VSS.n8217 84.2672
R1165 VSS.n8781 VSS.n8218 84.2672
R1166 VSS.n8781 VSS.n8219 84.2672
R1167 VSS.n8782 VSS.n8194 84.2672
R1168 VSS.n6231 VSS.n6213 84.2672
R1169 VSS.n6740 VSS.n6692 84.2672
R1170 VSS.n6745 VSS.n6740 84.2672
R1171 VSS.n9972 VSS.n6231 84.2672
R1172 VSS.n8148 VSS.n8016 84.2672
R1173 VSS.n8118 VSS.n8036 84.2672
R1174 VSS.n8118 VSS.n8037 84.2672
R1175 VSS.n8148 VSS.n8147 84.2672
R1176 VSS.n8871 VSS.n8001 84.2672
R1177 VSS.n8872 VSS.n7948 84.2672
R1178 VSS.n8877 VSS.n8872 84.2672
R1179 VSS.n8871 VSS.n8870 84.2672
R1180 VSS.n8819 VSS.n8186 84.2672
R1181 VSS.n8819 VSS.n8187 84.2672
R1182 VSS.n8820 VSS.n8162 84.2672
R1183 VSS.n9557 VSS.n7567 84.2672
R1184 VSS.n9557 VSS.n7568 84.2672
R1185 VSS.n9559 VSS.n7551 84.2672
R1186 VSS.n9510 VSS.n9291 84.2672
R1187 VSS.n9511 VSS.n8994 84.2672
R1188 VSS.n9511 VSS.n9290 84.2672
R1189 VSS.n9510 VSS.n9509 84.2672
R1190 VSS.n9832 VSS.n7184 84.2672
R1191 VSS.n9833 VSS.n7158 84.2672
R1192 VSS.n9833 VSS.n7183 84.2672
R1193 VSS.n9832 VSS.n9831 84.2672
R1194 VSS.n7372 VSS.n7260 84.2672
R1195 VSS.n7371 VSS.n7261 84.2672
R1196 VSS.n7371 VSS.n7262 84.2672
R1197 VSS.n7372 VSS.n7190 84.2672
R1198 VSS.n9245 VSS.n9160 84.2672
R1199 VSS.n9243 VSS.n9187 84.2672
R1200 VSS.n9243 VSS.n9188 84.2672
R1201 VSS.n9246 VSS.n9245 84.2672
R1202 VSS.n8952 VSS.n7849 84.2672
R1203 VSS.n8950 VSS.n7850 84.2672
R1204 VSS.n8950 VSS.n7851 84.2672
R1205 VSS.n8954 VSS.n8952 84.2672
R1206 VSS.n7805 VSS.n7640 84.2672
R1207 VSS.n8983 VSS.n7806 84.2672
R1208 VSS.n7806 VSS.n7636 84.2672
R1209 VSS.n7805 VSS.n7804 84.2672
R1210 VSS.n7726 VSS.n7675 84.2672
R1211 VSS.n7773 VSS.n7727 84.2672
R1212 VSS.n7727 VSS.n7671 84.2672
R1213 VSS.n7726 VSS.n7725 84.2672
R1214 VSS.n7142 VSS.n7070 84.2672
R1215 VSS.n7141 VSS.n7088 84.2672
R1216 VSS.n7141 VSS.n7089 84.2672
R1217 VSS.n9887 VSS.n7142 84.2672
R1218 VSS.n8926 VSS.n7939 84.2672
R1219 VSS.n8925 VSS.n7940 84.2672
R1220 VSS.n8925 VSS.n7941 84.2672
R1221 VSS.n8926 VSS.n7872 84.2672
R1222 VSS.n6904 VSS.n6609 84.2672
R1223 VSS.n6858 VSS.n6628 84.2672
R1224 VSS.n6858 VSS.n6629 84.2672
R1225 VSS.n6904 VSS.n6903 84.2672
R1226 VSS.n6925 VSS.n6580 84.2672
R1227 VSS.n6925 VSS.n6581 84.2672
R1228 VSS.n6977 VSS.n6976 84.2672
R1229 VSS.n7000 VSS.n6538 84.2672
R1230 VSS.n6998 VSS.n6539 84.2672
R1231 VSS.n6998 VSS.n6540 84.2672
R1232 VSS.n7036 VSS.n7000 84.2672
R1233 VSS.n7058 VSS.n6481 84.2672
R1234 VSS.n7057 VSS.n6482 84.2672
R1235 VSS.n7057 VSS.n6483 84.2672
R1236 VSS.n7058 VSS.n6271 84.2672
R1237 VSS.n6426 VSS.n6297 84.2672
R1238 VSS.n6425 VSS.n6315 84.2672
R1239 VSS.n6425 VSS.n6316 84.2672
R1240 VSS.n6449 VSS.n6426 84.2672
R1241 VSS.n6835 VSS.n6791 84.2672
R1242 VSS.n6790 VSS.n6675 84.2672
R1243 VSS.n6790 VSS.n6676 84.2672
R1244 VSS.n6791 VSS.n6657 84.2672
R1245 VSS.n6394 VSS.n6347 84.2672
R1246 VSS.n6395 VSS.n6394 84.2672
R1247 VSS.n11025 VSS.n3838 84.2672
R1248 VSS.n3880 VSS.n3853 84.2672
R1249 VSS.n10984 VSS.n3880 84.2672
R1250 VSS.n10919 VSS.n10900 84.2672
R1251 VSS.n7340 VSS.n7293 84.2672
R1252 VSS.n7341 VSS.n7340 84.2672
R1253 VSS.n10874 VSS.n3906 84.2672
R1254 VSS.n10771 VSS.n4132 84.2672
R1255 VSS.n4382 VSS.n4377 84.2672
R1256 VSS.n4270 VSS.n4266 84.2672
R1257 VSS.n4271 VSS.n4262 84.2672
R1258 VSS.n4298 VSS.n4271 84.2672
R1259 VSS.n4270 VSS.n4230 84.2672
R1260 VSS.n4383 VSS.n4201 84.2672
R1261 VSS.n4401 VSS.n4383 84.2672
R1262 VSS.n4382 VSS.n4162 84.2672
R1263 VSS.n10772 VSS.n4131 84.2672
R1264 VSS.n10773 VSS.n10772 84.2672
R1265 VSS.n10771 VSS.n10770 84.2672
R1266 VSS.n1392 VSS.n862 84.2672
R1267 VSS.n14198 VSS.n584 84.2672
R1268 VSS.n2398 VSS.n545 84.2672
R1269 VSS.n910 VSS.n604 84.2672
R1270 VSS.n1135 VSS.n604 84.2672
R1271 VSS.n14198 VSS.n14197 84.2672
R1272 VSS.n13050 VSS.n2480 84.2672
R1273 VSS.n13049 VSS.n2481 84.2672
R1274 VSS.n13049 VSS.n2482 84.2672
R1275 VSS.n13050 VSS.n2461 84.2672
R1276 VSS.n13092 VSS.n2392 84.2672
R1277 VSS.n13096 VSS.n2391 84.2672
R1278 VSS.n13097 VSS.n13096 84.2672
R1279 VSS.n13092 VSS.n13091 84.2672
R1280 VSS.n2347 VSS.n1911 84.2672
R1281 VSS.n2346 VSS.n1929 84.2672
R1282 VSS.n2346 VSS.n1930 84.2672
R1283 VSS.n13128 VSS.n2347 84.2672
R1284 VSS.n14157 VSS.n582 84.2672
R1285 VSS.n14225 VSS.n582 84.2672
R1286 VSS.n2403 VSS.n2398 84.2672
R1287 VSS.n1169 VSS.n881 84.2672
R1288 VSS.n1169 VSS.n882 84.2672
R1289 VSS.n1392 VSS.n1391 84.2672
R1290 VSS.n14109 VSS.n1461 84.2672
R1291 VSS.n14110 VSS.n628 84.2672
R1292 VSS.n14110 VSS.n1460 84.2672
R1293 VSS.n14109 VSS.n14108 84.2672
R1294 VSS.n13695 VSS.n13694 84.2672
R1295 VSS.n14077 VSS.n1670 84.2672
R1296 VSS.n1670 VSS.n1666 84.2672
R1297 VSS.n13695 VSS.n13652 84.2672
R1298 VSS.n13648 VSS.n13204 84.2672
R1299 VSS.n13647 VSS.n13222 84.2672
R1300 VSS.n13647 VSS.n13223 84.2672
R1301 VSS.n13898 VSS.n13648 84.2672
R1302 VSS.n1415 VSS.n813 84.2672
R1303 VSS.n1413 VSS.n840 84.2672
R1304 VSS.n1413 VSS.n841 84.2672
R1305 VSS.n1416 VSS.n1415 84.2672
R1306 VSS.n2239 VSS.n2054 84.2672
R1307 VSS.n2240 VSS.n1983 84.2672
R1308 VSS.n2240 VSS.n2053 84.2672
R1309 VSS.n2239 VSS.n2238 84.2672
R1310 VSS.n2174 VSS.n2103 84.2672
R1311 VSS.n2175 VSS.n2058 84.2672
R1312 VSS.n2175 VSS.n2102 84.2672
R1313 VSS.n2174 VSS.n2173 84.2672
R1314 VSS.n13193 VSS.n1851 84.2672
R1315 VSS.n13192 VSS.n1852 84.2672
R1316 VSS.n13192 VSS.n1853 84.2672
R1317 VSS.n13193 VSS.n1831 84.2672
R1318 VSS.n13926 VSS.n1813 84.2672
R1319 VSS.n13930 VSS.n1812 84.2672
R1320 VSS.n13931 VSS.n13930 84.2672
R1321 VSS.n13926 VSS.n13925 84.2672
R1322 VSS.n2277 VSS.n1977 84.2672
R1323 VSS.n2317 VSS.n2278 84.2672
R1324 VSS.n2278 VSS.n1948 84.2672
R1325 VSS.n2277 VSS.n2276 84.2672
R1326 VSS.n12979 VSS.n2661 84.2672
R1327 VSS.n12980 VSS.n2562 84.2672
R1328 VSS.n12980 VSS.n2660 84.2672
R1329 VSS.n12979 VSS.n12978 84.2672
R1330 VSS.n12947 VSS.n2697 84.2672
R1331 VSS.n2697 VSS.n2693 84.2672
R1332 VSS.n2812 VSS.n2770 84.2672
R1333 VSS.n12903 VSS.n2743 84.2672
R1334 VSS.n12903 VSS.n2841 84.2672
R1335 VSS.n12902 VSS.n12901 84.2672
R1336 VSS.n12636 VSS.n12635 84.2672
R1337 VSS.n12870 VSS.n2877 84.2672
R1338 VSS.n2877 VSS.n2873 84.2672
R1339 VSS.n12636 VSS.n3036 84.2672
R1340 VSS.n12721 VSS.n3018 84.2672
R1341 VSS.n12725 VSS.n3017 84.2672
R1342 VSS.n12726 VSS.n12725 84.2672
R1343 VSS.n12721 VSS.n12720 84.2672
R1344 VSS.n2632 VSS.n2590 84.2672
R1345 VSS.n13022 VSS.n2529 84.2672
R1346 VSS.n2529 VSS.n2500 84.2672
R1347 VSS.n2632 VSS.n2631 84.2672
R1348 VSS.n12759 VSS.n2943 84.2672
R1349 VSS.n12759 VSS.n2944 84.2672
R1350 VSS.n12779 VSS.n12760 84.2672
R1351 VSS.n1768 VSS.n1759 84.2672
R1352 VSS.n13963 VSS.n1768 84.2672
R1353 VSS.n1767 VSS.n1716 84.2672
R1354 VSS.n13582 VSS.n13510 84.2672
R1355 VSS.n13582 VSS.n13511 84.2672
R1356 VSS.n13586 VSS.n13481 84.2672
R1357 VSS.n13568 VSS.n13565 68.5719
R1358 VSS.n13566 VSS.n13561 68.5719
R1359 VSS.n13576 VSS.n13558 68.5719
R1360 VSS.n13579 VSS.n13578 68.5719
R1361 VSS.n13555 VSS.n13554 68.5719
R1362 VSS.n13516 VSS.n13513 68.5719
R1363 VSS.n13526 VSS.n13518 68.5719
R1364 VSS.n13524 VSS.n13523 68.5719
R1365 VSS.n13495 VSS.n13494 68.5719
R1366 VSS.n13499 VSS.n13489 68.5719
R1367 VSS.n13499 VSS.n13490 68.5719
R1368 VSS.n13605 VSS.n13483 68.5719
R1369 VSS.n13587 VSS.n13502 68.5719
R1370 VSS.n13601 VSS.n13506 68.5719
R1371 VSS.n13508 VSS.n13505 68.5719
R1372 VSS.n13594 VSS.n13593 68.5719
R1373 VSS.n13951 VSS.n13949 68.5719
R1374 VSS.n13956 VSS.n13944 68.5719
R1375 VSS.n13960 VSS.n13958 68.5719
R1376 VSS.n13964 VSS.n1769 68.5719
R1377 VSS.n13969 VSS.n13968 68.5719
R1378 VSS.n13985 VSS.n13971 68.5719
R1379 VSS.n13983 VSS.n13982 68.5719
R1380 VSS.n13976 VSS.n13974 68.5719
R1381 VSS.n1730 VSS.n1729 68.5719
R1382 VSS.n1734 VSS.n1724 68.5719
R1383 VSS.n1734 VSS.n1725 68.5719
R1384 VSS.n14018 VSS.n1718 68.5719
R1385 VSS.n1761 VSS.n1737 68.5719
R1386 VSS.n14014 VSS.n1741 68.5719
R1387 VSS.n1743 VSS.n1740 68.5719
R1388 VSS.n14007 VSS.n14006 68.5719
R1389 VSS.n12743 VSS.n12738 68.5719
R1390 VSS.n12747 VSS.n12745 68.5719
R1391 VSS.n12753 VSS.n2947 68.5719
R1392 VSS.n12756 VSS.n12755 68.5719
R1393 VSS.n2978 VSS.n2977 68.5719
R1394 VSS.n2994 VSS.n2980 68.5719
R1395 VSS.n2992 VSS.n2991 68.5719
R1396 VSS.n2985 VSS.n2983 68.5719
R1397 VSS.n12768 VSS.n12767 68.5719
R1398 VSS.n12763 VSS.n2940 68.5719
R1399 VSS.n12773 VSS.n2940 68.5719
R1400 VSS.n12776 VSS.n12775 68.5719
R1401 VSS.n12785 VSS.n12784 68.5719
R1402 VSS.n12798 VSS.n2932 68.5719
R1403 VSS.n12794 VSS.n2934 68.5719
R1404 VSS.n12788 VSS.n12787 68.5719
R1405 VSS.n2600 VSS.n2598 68.5719
R1406 VSS.n2604 VSS.n2593 68.5719
R1407 VSS.n2638 VSS.n2606 68.5719
R1408 VSS.n2636 VSS.n2635 68.5719
R1409 VSS.n2626 VSS.n2608 68.5719
R1410 VSS.n2628 VSS.n2625 68.5719
R1411 VSS.n2623 VSS.n2611 68.5719
R1412 VSS.n2618 VSS.n2616 68.5719
R1413 VSS.n2020 VSS.n2018 68.5719
R1414 VSS.n2024 VSS.n2013 68.5719
R1415 VSS.n2031 VSS.n2026 68.5719
R1416 VSS.n2029 VSS.n2028 68.5719
R1417 VSS.n2271 VSS.n1980 68.5719
R1418 VSS.n2273 VSS.n2270 68.5719
R1419 VSS.n2268 VSS.n2256 68.5719
R1420 VSS.n2263 VSS.n2261 68.5719
R1421 VSS.n829 VSS.n828 68.5719
R1422 VSS.n833 VSS.n824 68.5719
R1423 VSS.n1437 VSS.n816 68.5719
R1424 VSS.n835 VSS.n817 68.5719
R1425 VSS.n1433 VSS.n839 68.5719
R1426 VSS.n1428 VSS.n838 68.5719
R1427 VSS.n1426 VSS.n1425 68.5719
R1428 VSS.n1421 VSS.n1420 68.5719
R1429 VSS.n7287 VSS.n7282 68.5719
R1430 VSS.n7290 VSS.n7289 68.5719
R1431 VSS.n7347 VSS.n7345 68.5719
R1432 VSS.n7343 VSS.n7292 68.5719
R1433 VSS.n7336 VSS.n7335 68.5719
R1434 VSS.n7298 VSS.n7295 68.5719
R1435 VSS.n7308 VSS.n7300 68.5719
R1436 VSS.n7306 VSS.n7305 68.5719
R1437 VSS.n10863 VSS.n10862 68.5719
R1438 VSS.n10858 VSS.n3903 68.5719
R1439 VSS.n10868 VSS.n3903 68.5719
R1440 VSS.n10871 VSS.n10870 68.5719
R1441 VSS.n10880 VSS.n10879 68.5719
R1442 VSS.n10893 VSS.n3895 68.5719
R1443 VSS.n10889 VSS.n3897 68.5719
R1444 VSS.n10883 VSS.n10882 68.5719
R1445 VSS.n10974 VSS.n10973 68.5719
R1446 VSS.n10970 VSS.n10969 68.5719
R1447 VSS.n10981 VSS.n10980 68.5719
R1448 VSS.n10985 VSS.n3878 68.5719
R1449 VSS.n3861 VSS.n3860 68.5719
R1450 VSS.n10989 VSS.n3855 68.5719
R1451 VSS.n3866 VSS.n3857 68.5719
R1452 VSS.n3871 VSS.n3865 68.5719
R1453 VSS.n10909 VSS.n10907 68.5719
R1454 VSS.n10913 VSS.n10902 68.5719
R1455 VSS.n10914 VSS.n10913 68.5719
R1456 VSS.n10949 VSS.n10916 68.5719
R1457 VSS.n10943 VSS.n10918 68.5719
R1458 VSS.n10938 VSS.n10923 68.5719
R1459 VSS.n10936 VSS.n10935 68.5719
R1460 VSS.n10933 VSS.n10926 68.5719
R1461 VSS.n6341 VSS.n6336 68.5719
R1462 VSS.n6344 VSS.n6343 68.5719
R1463 VSS.n6401 VSS.n6399 68.5719
R1464 VSS.n6397 VSS.n6346 68.5719
R1465 VSS.n6390 VSS.n6389 68.5719
R1466 VSS.n6352 VSS.n6349 68.5719
R1467 VSS.n6362 VSS.n6354 68.5719
R1468 VSS.n6360 VSS.n6359 68.5719
R1469 VSS.n11014 VSS.n11013 68.5719
R1470 VSS.n11009 VSS.n3835 68.5719
R1471 VSS.n11019 VSS.n3835 68.5719
R1472 VSS.n11022 VSS.n11021 68.5719
R1473 VSS.n11031 VSS.n11030 68.5719
R1474 VSS.n11044 VSS.n3827 68.5719
R1475 VSS.n11040 VSS.n3829 68.5719
R1476 VSS.n11034 VSS.n11033 68.5719
R1477 VSS.n6823 VSS.n6821 68.5719
R1478 VSS.n6828 VSS.n6816 68.5719
R1479 VSS.n6832 VSS.n6830 68.5719
R1480 VSS.n6836 VSS.n6792 68.5719
R1481 VSS.n6841 VSS.n6840 68.5719
R1482 VSS.n6843 VSS.n6660 68.5719
R1483 VSS.n6672 VSS.n6663 68.5719
R1484 VSS.n6668 VSS.n6667 68.5719
R1485 VSS.n7925 VSS.n7924 68.5719
R1486 VSS.n7930 VSS.n7929 68.5719
R1487 VSS.n7934 VSS.n7933 68.5719
R1488 VSS.n7938 VSS.n7937 68.5719
R1489 VSS.n8930 VSS.n8929 68.5719
R1490 VSS.n8934 VSS.n7874 68.5719
R1491 VSS.n7886 VSS.n7876 68.5719
R1492 VSS.n7880 VSS.n7879 68.5719
R1493 VSS.n9176 VSS.n9175 68.5719
R1494 VSS.n9180 VSS.n9171 68.5719
R1495 VSS.n9267 VSS.n9163 68.5719
R1496 VSS.n9182 VSS.n9164 68.5719
R1497 VSS.n9263 VSS.n9186 68.5719
R1498 VSS.n9258 VSS.n9185 68.5719
R1499 VSS.n9256 VSS.n9255 68.5719
R1500 VSS.n9251 VSS.n9250 68.5719
R1501 VSS.n8273 VSS.n8272 68.5719
R1502 VSS.n8277 VSS.n8276 68.5719
R1503 VSS.n8282 VSS.n8281 68.5719
R1504 VSS.n9554 VSS.n9553 68.5719
R1505 VSS.n9551 VSS.n7572 68.5719
R1506 VSS.n7584 VSS.n7576 68.5719
R1507 VSS.n7582 VSS.n7581 68.5719
R1508 VSS.n8498 VSS.n8497 68.5719
R1509 VSS.n8502 VSS.n8501 68.5719
R1510 VSS.n8506 VSS.n8505 68.5719
R1511 VSS.n8824 VSS.n8823 68.5719
R1512 VSS.n8828 VSS.n8164 68.5719
R1513 VSS.n8175 VSS.n8166 68.5719
R1514 VSS.n8169 VSS.n8168 68.5719
R1515 VSS.n8377 VSS.n8376 68.5719
R1516 VSS.n8381 VSS.n8380 68.5719
R1517 VSS.n8386 VSS.n8385 68.5719
R1518 VSS.n8816 VSS.n8815 68.5719
R1519 VSS.n8813 VSS.n8191 68.5719
R1520 VSS.n8807 VSS.n8806 68.5719
R1521 VSS.n8804 VSS.n8799 68.5719
R1522 VSS.n8397 VSS.n8396 68.5719
R1523 VSS.n8401 VSS.n8400 68.5719
R1524 VSS.n8405 VSS.n8404 68.5719
R1525 VSS.n8786 VSS.n8785 68.5719
R1526 VSS.n8790 VSS.n8196 68.5719
R1527 VSS.n8207 VSS.n8198 68.5719
R1528 VSS.n8201 VSS.n8200 68.5719
R1529 VSS.n8253 VSS.n8248 68.5719
R1530 VSS.n8254 VSS.n8253 68.5719
R1531 VSS.n8258 VSS.n8257 68.5719
R1532 VSS.n8775 VSS.n8244 68.5719
R1533 VSS.n8242 VSS.n8241 68.5719
R1534 VSS.n8239 VSS.n8221 68.5719
R1535 VSS.n8234 VSS.n8233 68.5719
R1536 VSS.n8231 VSS.n8225 68.5719
R1537 VSS.n8857 VSS.n8851 68.5719
R1538 VSS.n8861 VSS.n8859 68.5719
R1539 VSS.n8865 VSS.n8005 68.5719
R1540 VSS.n8869 VSS.n8867 68.5719
R1541 VSS.n8069 VSS.n8068 68.5719
R1542 VSS.n8071 VSS.n8066 68.5719
R1543 VSS.n8064 VSS.n8053 68.5719
R1544 VSS.n8060 VSS.n8058 68.5719
R1545 VSS.n9960 VSS.n9958 68.5719
R1546 VSS.n9965 VSS.n9953 68.5719
R1547 VSS.n9969 VSS.n9967 68.5719
R1548 VSS.n9973 VSS.n6232 68.5719
R1549 VSS.n9978 VSS.n9977 68.5719
R1550 VSS.n9980 VSS.n6216 68.5719
R1551 VSS.n6223 VSS.n6222 68.5719
R1552 VSS.n6228 VSS.n6220 68.5719
R1553 VSS.n6756 VSS.n6755 68.5719
R1554 VSS.n6752 VSS.n6751 68.5719
R1555 VSS.n6748 VSS.n6747 68.5719
R1556 VSS.n6711 VSS.n6710 68.5719
R1557 VSS.n6764 VSS.n6763 68.5719
R1558 VSS.n6708 VSS.n6696 68.5719
R1559 VSS.n6702 VSS.n6700 68.5719
R1560 VSS.n8028 VSS.n8022 68.5719
R1561 VSS.n8032 VSS.n8023 68.5719
R1562 VSS.n8154 VSS.n8153 68.5719
R1563 VSS.n8126 VSS.n8120 68.5719
R1564 VSS.n8143 VSS.n8128 68.5719
R1565 VSS.n8141 VSS.n8140 68.5719
R1566 VSS.n8137 VSS.n8136 68.5719
R1567 VSS.n8109 VSS.n8108 68.5719
R1568 VSS.n8105 VSS.n8104 68.5719
R1569 VSS.n8101 VSS.n8100 68.5719
R1570 VSS.n8115 VSS.n8040 68.5719
R1571 VSS.n8090 VSS.n8046 68.5719
R1572 VSS.n8084 VSS.n8083 68.5719
R1573 VSS.n8080 VSS.n8079 68.5719
R1574 VSS.n8888 VSS.n8887 68.5719
R1575 VSS.n8884 VSS.n8883 68.5719
R1576 VSS.n8880 VSS.n8879 68.5719
R1577 VSS.n7968 VSS.n7967 68.5719
R1578 VSS.n8896 VSS.n8895 68.5719
R1579 VSS.n7965 VSS.n7952 68.5719
R1580 VSS.n7959 VSS.n7957 68.5719
R1581 VSS.n9588 VSS.n9579 68.5719
R1582 VSS.n9591 VSS.n9590 68.5719
R1583 VSS.n9593 VSS.n7554 68.5719
R1584 VSS.n7557 VSS.n7554 68.5719
R1585 VSS.n9561 VSS.n9560 68.5719
R1586 VSS.n9566 VSS.n9565 68.5719
R1587 VSS.n9569 VSS.n9568 68.5719
R1588 VSS.n9575 VSS.n7563 68.5719
R1589 VSS.n9277 VSS.n9276 68.5719
R1590 VSS.n9283 VSS.n9282 68.5719
R1591 VSS.n9286 VSS.n9285 68.5719
R1592 VSS.n9515 VSS.n9514 68.5719
R1593 VSS.n9518 VSS.n8996 68.5719
R1594 VSS.n9013 VSS.n8998 68.5719
R1595 VSS.n9007 VSS.n9006 68.5719
R1596 VSS.n9501 VSS.n9491 68.5719
R1597 VSS.n9504 VSS.n9503 68.5719
R1598 VSS.n9506 VSS.n9489 68.5719
R1599 VSS.n9489 VSS.n9319 68.5719
R1600 VSS.n9314 VSS.n9313 68.5719
R1601 VSS.n9310 VSS.n9309 68.5719
R1602 VSS.n9307 VSS.n9295 68.5719
R1603 VSS.n9302 VSS.n9300 68.5719
R1604 VSS.n9818 VSS.n9816 68.5719
R1605 VSS.n9823 VSS.n9811 68.5719
R1606 VSS.n9828 VSS.n9825 68.5719
R1607 VSS.n9826 VSS.n7188 68.5719
R1608 VSS.n7222 VSS.n7221 68.5719
R1609 VSS.n7225 VSS.n7222 68.5719
R1610 VSS.n7237 VSS.n7227 68.5719
R1611 VSS.n7235 VSS.n7234 68.5719
R1612 VSS.n7232 VSS.n7229 68.5719
R1613 VSS.n9475 VSS.n9474 68.5719
R1614 VSS.n9482 VSS.n9477 68.5719
R1615 VSS.n9479 VSS.n9478 68.5719
R1616 VSS.n9837 VSS.n9836 68.5719
R1617 VSS.n9840 VSS.n7160 68.5719
R1618 VSS.n7177 VSS.n7162 68.5719
R1619 VSS.n7171 VSS.n7170 68.5719
R1620 VSS.n7200 VSS.n7199 68.5719
R1621 VSS.n7206 VSS.n7197 68.5719
R1622 VSS.n7196 VSS.n7192 68.5719
R1623 VSS.n7376 VSS.n7375 68.5719
R1624 VSS.n7259 VSS.n7258 68.5719
R1625 VSS.n7256 VSS.n7212 68.5719
R1626 VSS.n7247 VSS.n7214 68.5719
R1627 VSS.n7249 VSS.n7246 68.5719
R1628 VSS.n7356 VSS.n7355 68.5719
R1629 VSS.n7360 VSS.n7359 68.5719
R1630 VSS.n7366 VSS.n7275 68.5719
R1631 VSS.n7366 VSS.n7276 68.5719
R1632 VSS.n7368 VSS.n7265 68.5719
R1633 VSS.n7317 VSS.n7316 68.5719
R1634 VSS.n7326 VSS.n7325 68.5719
R1635 VSS.n7321 VSS.n7319 68.5719
R1636 VSS.n9201 VSS.n9191 68.5719
R1637 VSS.n9205 VSS.n9203 68.5719
R1638 VSS.n9210 VSS.n9189 68.5719
R1639 VSS.n9240 VSS.n9239 68.5719
R1640 VSS.n9237 VSS.n9216 68.5719
R1641 VSS.n9228 VSS.n9220 68.5719
R1642 VSS.n9226 VSS.n9225 68.5719
R1643 VSS.n7835 VSS.n7834 68.5719
R1644 VSS.n7840 VSS.n7839 68.5719
R1645 VSS.n7842 VSS.n7829 68.5719
R1646 VSS.n8956 VSS.n7830 68.5719
R1647 VSS.n7848 VSS.n7827 68.5719
R1648 VSS.n7845 VSS.n7827 68.5719
R1649 VSS.n8960 VSS.n7812 68.5719
R1650 VSS.n7820 VSS.n7813 68.5719
R1651 VSS.n7824 VSS.n7818 68.5719
R1652 VSS.n7904 VSS.n7903 68.5719
R1653 VSS.n7914 VSS.n7906 68.5719
R1654 VSS.n7912 VSS.n7911 68.5719
R1655 VSS.n8947 VSS.n8946 68.5719
R1656 VSS.n8944 VSS.n7855 68.5719
R1657 VSS.n7867 VSS.n7859 68.5719
R1658 VSS.n7865 VSS.n7864 68.5719
R1659 VSS.n7791 VSS.n7789 68.5719
R1660 VSS.n7796 VSS.n7784 68.5719
R1661 VSS.n7801 VSS.n7798 68.5719
R1662 VSS.n7799 VSS.n7644 68.5719
R1663 VSS.n7735 VSS.n7734 68.5719
R1664 VSS.n7738 VSS.n7735 68.5719
R1665 VSS.n7750 VSS.n7740 68.5719
R1666 VSS.n7748 VSS.n7747 68.5719
R1667 VSS.n7745 VSS.n7742 68.5719
R1668 VSS.n7622 VSS.n7621 68.5719
R1669 VSS.n8987 VSS.n7613 68.5719
R1670 VSS.n7634 VSS.n7615 68.5719
R1671 VSS.n8984 VSS.n7633 68.5719
R1672 VSS.n8979 VSS.n8967 68.5719
R1673 VSS.n8969 VSS.n8968 68.5719
R1674 VSS.n8973 VSS.n8972 68.5719
R1675 VSS.n7712 VSS.n7710 68.5719
R1676 VSS.n7717 VSS.n7705 68.5719
R1677 VSS.n7722 VSS.n7719 68.5719
R1678 VSS.n7720 VSS.n7703 68.5719
R1679 VSS.n7698 VSS.n7697 68.5719
R1680 VSS.n7697 VSS.n7676 68.5719
R1681 VSS.n7692 VSS.n7691 68.5719
R1682 VSS.n7689 VSS.n7679 68.5719
R1683 VSS.n7684 VSS.n7683 68.5719
R1684 VSS.n7657 VSS.n7656 68.5719
R1685 VSS.n7777 VSS.n7648 68.5719
R1686 VSS.n7669 VSS.n7650 68.5719
R1687 VSS.n7774 VSS.n7668 68.5719
R1688 VSS.n7769 VSS.n7757 68.5719
R1689 VSS.n7759 VSS.n7758 68.5719
R1690 VSS.n7763 VSS.n7762 68.5719
R1691 VSS.n9875 VSS.n9873 68.5719
R1692 VSS.n9880 VSS.n9868 68.5719
R1693 VSS.n9884 VSS.n9882 68.5719
R1694 VSS.n9888 VSS.n7143 68.5719
R1695 VSS.n9893 VSS.n9892 68.5719
R1696 VSS.n9895 VSS.n7073 68.5719
R1697 VSS.n7080 VSS.n7079 68.5719
R1698 VSS.n7085 VSS.n7077 68.5719
R1699 VSS.n7125 VSS.n7124 68.5719
R1700 VSS.n7130 VSS.n7129 68.5719
R1701 VSS.n7136 VSS.n7119 68.5719
R1702 VSS.n7136 VSS.n7120 68.5719
R1703 VSS.n7138 VSS.n7092 68.5719
R1704 VSS.n7114 VSS.n7098 68.5719
R1705 VSS.n7109 VSS.n7108 68.5719
R1706 VSS.n7103 VSS.n7102 68.5719
R1707 VSS.n7983 VSS.n7982 68.5719
R1708 VSS.n7990 VSS.n7979 68.5719
R1709 VSS.n7996 VSS.n7992 68.5719
R1710 VSS.n7994 VSS.n7993 68.5719
R1711 VSS.n8922 VSS.n8921 68.5719
R1712 VSS.n8919 VSS.n7945 68.5719
R1713 VSS.n8913 VSS.n8912 68.5719
R1714 VSS.n8910 VSS.n8905 68.5719
R1715 VSS.n6801 VSS.n6800 68.5719
R1716 VSS.n6808 VSS.n6803 68.5719
R1717 VSS.n6805 VSS.n6804 68.5719
R1718 VSS.n6855 VSS.n6632 68.5719
R1719 VSS.n6852 VSS.n6642 68.5719
R1720 VSS.n6652 VSS.n6646 68.5719
R1721 VSS.n6649 VSS.n6647 68.5719
R1722 VSS.n6890 VSS.n6888 68.5719
R1723 VSS.n6895 VSS.n6883 68.5719
R1724 VSS.n6900 VSS.n6897 68.5719
R1725 VSS.n6898 VSS.n6860 68.5719
R1726 VSS.n6908 VSS.n6907 68.5719
R1727 VSS.n6910 VSS.n6612 68.5719
R1728 VSS.n6624 VSS.n6615 68.5719
R1729 VSS.n6620 VSS.n6619 68.5719
R1730 VSS.n6869 VSS.n6868 68.5719
R1731 VSS.n6876 VSS.n6871 68.5719
R1732 VSS.n6873 VSS.n6872 68.5719
R1733 VSS.n6922 VSS.n6584 68.5719
R1734 VSS.n6919 VSS.n6594 68.5719
R1735 VSS.n6604 VSS.n6598 68.5719
R1736 VSS.n6601 VSS.n6599 68.5719
R1737 VSS.n6963 VSS.n6961 68.5719
R1738 VSS.n6968 VSS.n6956 68.5719
R1739 VSS.n6973 VSS.n6970 68.5719
R1740 VSS.n6971 VSS.n6927 68.5719
R1741 VSS.n6981 VSS.n6980 68.5719
R1742 VSS.n6983 VSS.n6564 68.5719
R1743 VSS.n6576 VSS.n6567 68.5719
R1744 VSS.n6572 VSS.n6571 68.5719
R1745 VSS.n7005 VSS.n7004 68.5719
R1746 VSS.n7011 VSS.n7010 68.5719
R1747 VSS.n7008 VSS.n6531 68.5719
R1748 VSS.n7038 VSS.n6532 68.5719
R1749 VSS.n6537 VSS.n6529 68.5719
R1750 VSS.n6534 VSS.n6529 68.5719
R1751 VSS.n7042 VSS.n6514 68.5719
R1752 VSS.n6522 VSS.n6515 68.5719
R1753 VSS.n6526 VSS.n6520 68.5719
R1754 VSS.n6939 VSS.n6938 68.5719
R1755 VSS.n6949 VSS.n6941 68.5719
R1756 VSS.n6947 VSS.n6946 68.5719
R1757 VSS.n6995 VSS.n6994 68.5719
R1758 VSS.n6992 VSS.n6544 68.5719
R1759 VSS.n6556 VSS.n6548 68.5719
R1760 VSS.n6554 VSS.n6553 68.5719
R1761 VSS.n6282 VSS.n6281 68.5719
R1762 VSS.n6286 VSS.n6277 68.5719
R1763 VSS.n6287 VSS.n6273 68.5719
R1764 VSS.n7062 VSS.n7061 68.5719
R1765 VSS.n6480 VSS.n6479 68.5719
R1766 VSS.n6479 VSS.n6478 68.5719
R1767 VSS.n6476 VSS.n6294 68.5719
R1768 VSS.n6470 VSS.n6466 68.5719
R1769 VSS.n6468 VSS.n6467 68.5719
R1770 VSS.n7022 VSS.n7021 68.5719
R1771 VSS.n7029 VSS.n7024 68.5719
R1772 VSS.n7026 VSS.n7025 68.5719
R1773 VSS.n7054 VSS.n6486 68.5719
R1774 VSS.n7051 VSS.n6496 68.5719
R1775 VSS.n6506 VSS.n6500 68.5719
R1776 VSS.n6503 VSS.n6501 68.5719
R1777 VSS.n6437 VSS.n6435 68.5719
R1778 VSS.n6442 VSS.n6430 68.5719
R1779 VSS.n6446 VSS.n6444 68.5719
R1780 VSS.n6450 VSS.n6427 68.5719
R1781 VSS.n6455 VSS.n6454 68.5719
R1782 VSS.n6457 VSS.n6300 68.5719
R1783 VSS.n6307 VSS.n6306 68.5719
R1784 VSS.n6312 VSS.n6304 68.5719
R1785 VSS.n6410 VSS.n6409 68.5719
R1786 VSS.n6414 VSS.n6413 68.5719
R1787 VSS.n6420 VSS.n6329 68.5719
R1788 VSS.n6420 VSS.n6330 68.5719
R1789 VSS.n6422 VSS.n6319 68.5719
R1790 VSS.n6371 VSS.n6370 68.5719
R1791 VSS.n6380 VSS.n6379 68.5719
R1792 VSS.n6375 VSS.n6373 68.5719
R1793 VSS.n6722 VSS.n6721 68.5719
R1794 VSS.n6728 VSS.n6727 68.5719
R1795 VSS.n6734 VSS.n6733 68.5719
R1796 VSS.n6731 VSS.n6684 68.5719
R1797 VSS.n6787 VSS.n6679 68.5719
R1798 VSS.n6784 VSS.n6688 68.5719
R1799 VSS.n6778 VSS.n6777 68.5719
R1800 VSS.n6774 VSS.n6773 68.5719
R1801 VSS.n4125 VSS.n4121 68.5719
R1802 VSS.n4120 VSS.n4110 68.5719
R1803 VSS.n10778 VSS.n4112 68.5719
R1804 VSS.n10774 VSS.n4129 68.5719
R1805 VSS.n4416 VSS.n4415 68.5719
R1806 VSS.n4429 VSS.n4418 68.5719
R1807 VSS.n4426 VSS.n4419 68.5719
R1808 VSS.n4421 VSS.n4420 68.5719
R1809 VSS.n4389 VSS.n4388 68.5719
R1810 VSS.n4394 VSS.n4393 68.5719
R1811 VSS.n4398 VSS.n4397 68.5719
R1812 VSS.n4402 VSS.n4198 68.5719
R1813 VSS.n4200 VSS.n4195 68.5719
R1814 VSS.n4211 VSS.n4195 68.5719
R1815 VSS.n4222 VSS.n4221 68.5719
R1816 VSS.n4219 VSS.n4218 68.5719
R1817 VSS.n4215 VSS.n4187 68.5719
R1818 VSS.n10757 VSS.n10755 68.5719
R1819 VSS.n10762 VSS.n10750 68.5719
R1820 VSS.n10763 VSS.n10762 68.5719
R1821 VSS.n10767 VSS.n10766 68.5719
R1822 VSS.n4449 VSS.n4448 68.5719
R1823 VSS.n4446 VSS.n4136 68.5719
R1824 VSS.n4149 VSS.n4148 68.5719
R1825 VSS.n4146 VSS.n4141 68.5719
R1826 VSS.n4175 VSS.n4171 68.5719
R1827 VSS.n4173 VSS.n4172 68.5719
R1828 VSS.n4407 VSS.n4164 68.5719
R1829 VSS.n4362 VSS.n4361 68.5719
R1830 VSS.n4373 VSS.n4186 68.5719
R1831 VSS.n4363 VSS.n4186 68.5719
R1832 VSS.n4367 VSS.n4366 68.5719
R1833 VSS.n4286 VSS.n4284 68.5719
R1834 VSS.n4291 VSS.n4279 68.5719
R1835 VSS.n4295 VSS.n4293 68.5719
R1836 VSS.n4299 VSS.n4272 68.5719
R1837 VSS.n4304 VSS.n4303 68.5719
R1838 VSS.n4320 VSS.n4306 68.5719
R1839 VSS.n4318 VSS.n4317 68.5719
R1840 VSS.n4311 VSS.n4309 68.5719
R1841 VSS.n4244 VSS.n4243 68.5719
R1842 VSS.n4248 VSS.n4238 68.5719
R1843 VSS.n4248 VSS.n4239 68.5719
R1844 VSS.n4346 VSS.n4232 68.5719
R1845 VSS.n4264 VSS.n4251 68.5719
R1846 VSS.n4342 VSS.n4255 68.5719
R1847 VSS.n4257 VSS.n4254 68.5719
R1848 VSS.n4335 VSS.n4334 68.5719
R1849 VSS.n944 VSS.n943 68.5719
R1850 VSS.n948 VSS.n947 68.5719
R1851 VSS.n952 VSS.n951 68.5719
R1852 VSS.n1166 VSS.n885 68.5719
R1853 VSS.n1163 VSS.n895 68.5719
R1854 VSS.n905 VSS.n899 68.5719
R1855 VSS.n902 VSS.n900 68.5719
R1856 VSS.n596 VSS.n590 68.5719
R1857 VSS.n600 VSS.n591 68.5719
R1858 VSS.n14204 VSS.n14203 68.5719
R1859 VSS.n14176 VSS.n606 68.5719
R1860 VSS.n14193 VSS.n14178 68.5719
R1861 VSS.n14191 VSS.n14190 68.5719
R1862 VSS.n14187 VSS.n14186 68.5719
R1863 VSS.n14213 VSS.n14212 68.5719
R1864 VSS.n14218 VSS.n14217 68.5719
R1865 VSS.n14222 VSS.n14221 68.5719
R1866 VSS.n14226 VSS.n580 68.5719
R1867 VSS.n14156 VSS.n577 68.5719
R1868 VSS.n14159 VSS.n577 68.5719
R1869 VSS.n14170 VSS.n14169 68.5719
R1870 VSS.n14167 VSS.n14166 68.5719
R1871 VSS.n14163 VSS.n569 68.5719
R1872 VSS.n562 VSS.n561 68.5719
R1873 VSS.n568 VSS.n558 68.5719
R1874 VSS.n568 VSS.n559 68.5719
R1875 VSS.n14232 VSS.n14231 68.5719
R1876 VSS.n2406 VSS.n2405 68.5719
R1877 VSS.n2416 VSS.n554 68.5719
R1878 VSS.n2413 VSS.n554 68.5719
R1879 VSS.n2411 VSS.n2410 68.5719
R1880 VSS.n1146 VSS.n1145 68.5719
R1881 VSS.n1142 VSS.n1141 68.5719
R1882 VSS.n1138 VSS.n1137 68.5719
R1883 VSS.n929 VSS.n928 68.5719
R1884 VSS.n1154 VSS.n1153 68.5719
R1885 VSS.n926 VSS.n914 68.5719
R1886 VSS.n920 VSS.n918 68.5719
R1887 VSS.n13116 VSS.n13114 68.5719
R1888 VSS.n13121 VSS.n13109 68.5719
R1889 VSS.n13125 VSS.n13123 68.5719
R1890 VSS.n13129 VSS.n2348 68.5719
R1891 VSS.n13134 VSS.n13133 68.5719
R1892 VSS.n13136 VSS.n1914 68.5719
R1893 VSS.n1921 VSS.n1920 68.5719
R1894 VSS.n1926 VSS.n1918 68.5719
R1895 VSS.n2470 VSS.n2469 68.5719
R1896 VSS.n2476 VSS.n2467 68.5719
R1897 VSS.n13056 VSS.n2464 68.5719
R1898 VSS.n13054 VSS.n13053 68.5719
R1899 VSS.n12415 VSS.n12414 68.5719
R1900 VSS.n12417 VSS.n12413 68.5719
R1901 VSS.n12411 VSS.n12400 68.5719
R1902 VSS.n12407 VSS.n12405 68.5719
R1903 VSS.n13034 VSS.n13033 68.5719
R1904 VSS.n13038 VSS.n13037 68.5719
R1905 VSS.n13044 VSS.n2495 68.5719
R1906 VSS.n13044 VSS.n2496 68.5719
R1907 VSS.n13046 VSS.n2485 68.5719
R1908 VSS.n2536 VSS.n2535 68.5719
R1909 VSS.n2545 VSS.n2544 68.5719
R1910 VSS.n2540 VSS.n2538 68.5719
R1911 VSS.n2439 VSS.n2438 68.5719
R1912 VSS.n2443 VSS.n2442 68.5719
R1913 VSS.n2450 VSS.n2393 68.5719
R1914 VSS.n13070 VSS.n2457 68.5719
R1915 VSS.n13087 VSS.n13072 68.5719
R1916 VSS.n13085 VSS.n13084 68.5719
R1917 VSS.n13081 VSS.n13080 68.5719
R1918 VSS.n2369 VSS.n2365 68.5719
R1919 VSS.n13103 VSS.n2354 68.5719
R1920 VSS.n13100 VSS.n2355 68.5719
R1921 VSS.n13100 VSS.n2371 68.5719
R1922 VSS.n2373 VSS.n2363 68.5719
R1923 VSS.n2387 VSS.n2375 68.5719
R1924 VSS.n2385 VSS.n2384 68.5719
R1925 VSS.n2379 VSS.n2378 68.5719
R1926 VSS.n2337 VSS.n2336 68.5719
R1927 VSS.n2333 VSS.n2332 68.5719
R1928 VSS.n2329 VSS.n2328 68.5719
R1929 VSS.n2343 VSS.n1933 68.5719
R1930 VSS.n2294 VSS.n2293 68.5719
R1931 VSS.n2290 VSS.n2289 68.5719
R1932 VSS.n2286 VSS.n2285 68.5719
R1933 VSS.n1383 VSS.n1373 68.5719
R1934 VSS.n1386 VSS.n1385 68.5719
R1935 VSS.n1388 VSS.n1371 68.5719
R1936 VSS.n1371 VSS.n1171 68.5719
R1937 VSS.n1396 VSS.n1395 68.5719
R1938 VSS.n1398 VSS.n865 68.5719
R1939 VSS.n872 VSS.n871 68.5719
R1940 VSS.n877 VSS.n869 68.5719
R1941 VSS.n1447 VSS.n1446 68.5719
R1942 VSS.n1453 VSS.n1452 68.5719
R1943 VSS.n1456 VSS.n1455 68.5719
R1944 VSS.n14114 VSS.n14113 68.5719
R1945 VSS.n14117 VSS.n630 68.5719
R1946 VSS.n647 VSS.n632 68.5719
R1947 VSS.n641 VSS.n640 68.5719
R1948 VSS.n14100 VSS.n14090 68.5719
R1949 VSS.n14103 VSS.n14102 68.5719
R1950 VSS.n14105 VSS.n14088 68.5719
R1951 VSS.n14088 VSS.n1465 68.5719
R1952 VSS.n1688 VSS.n1686 68.5719
R1953 VSS.n1691 VSS.n1690 68.5719
R1954 VSS.n1693 VSS.n1683 68.5719
R1955 VSS.n1681 VSS.n1676 68.5719
R1956 VSS.n13661 VSS.n13659 68.5719
R1957 VSS.n13665 VSS.n13654 68.5719
R1958 VSS.n13668 VSS.n13667 68.5719
R1959 VSS.n13699 VSS.n13698 68.5719
R1960 VSS.n13693 VSS.n13692 68.5719
R1961 VSS.n13692 VSS.n13691 68.5719
R1962 VSS.n13689 VSS.n13674 68.5719
R1963 VSS.n13683 VSS.n13679 68.5719
R1964 VSS.n13681 VSS.n13680 68.5719
R1965 VSS.n1652 VSS.n1651 68.5719
R1966 VSS.n14081 VSS.n1643 68.5719
R1967 VSS.n1664 VSS.n1645 68.5719
R1968 VSS.n14078 VSS.n1663 68.5719
R1969 VSS.n14073 VSS.n14061 68.5719
R1970 VSS.n14063 VSS.n14062 68.5719
R1971 VSS.n14067 VSS.n14066 68.5719
R1972 VSS.n13886 VSS.n13884 68.5719
R1973 VSS.n13891 VSS.n13879 68.5719
R1974 VSS.n13895 VSS.n13893 68.5719
R1975 VSS.n13899 VSS.n13649 68.5719
R1976 VSS.n13904 VSS.n13903 68.5719
R1977 VSS.n13906 VSS.n13207 68.5719
R1978 VSS.n13214 VSS.n13213 68.5719
R1979 VSS.n13219 VSS.n13211 68.5719
R1980 VSS.n13632 VSS.n13631 68.5719
R1981 VSS.n13636 VSS.n13635 68.5719
R1982 VSS.n13642 VSS.n13236 68.5719
R1983 VSS.n13642 VSS.n13237 68.5719
R1984 VSS.n13644 VSS.n13226 68.5719
R1985 VSS.n13535 VSS.n13534 68.5719
R1986 VSS.n13544 VSS.n13543 68.5719
R1987 VSS.n13539 VSS.n13537 68.5719
R1988 VSS.n1184 VSS.n1183 68.5719
R1989 VSS.n1188 VSS.n1187 68.5719
R1990 VSS.n1193 VSS.n1192 68.5719
R1991 VSS.n1410 VSS.n1409 68.5719
R1992 VSS.n1407 VSS.n845 68.5719
R1993 VSS.n857 VSS.n849 68.5719
R1994 VSS.n855 VSS.n854 68.5719
R1995 VSS.n2225 VSS.n2223 68.5719
R1996 VSS.n2230 VSS.n2218 68.5719
R1997 VSS.n2235 VSS.n2232 68.5719
R1998 VSS.n2233 VSS.n2215 68.5719
R1999 VSS.n2210 VSS.n2209 68.5719
R2000 VSS.n2209 VSS.n2055 68.5719
R2001 VSS.n2202 VSS.n2192 68.5719
R2002 VSS.n2200 VSS.n2199 68.5719
R2003 VSS.n2197 VSS.n2194 68.5719
R2004 VSS.n2041 VSS.n2040 68.5719
R2005 VSS.n2047 VSS.n2046 68.5719
R2006 VSS.n2050 VSS.n2049 68.5719
R2007 VSS.n2244 VSS.n2243 68.5719
R2008 VSS.n2247 VSS.n1985 68.5719
R2009 VSS.n2002 VSS.n1987 68.5719
R2010 VSS.n1996 VSS.n1995 68.5719
R2011 VSS.n2160 VSS.n2158 68.5719
R2012 VSS.n2165 VSS.n2153 68.5719
R2013 VSS.n2170 VSS.n2167 68.5719
R2014 VSS.n2168 VSS.n2131 68.5719
R2015 VSS.n2126 VSS.n2125 68.5719
R2016 VSS.n2125 VSS.n2104 68.5719
R2017 VSS.n2120 VSS.n2119 68.5719
R2018 VSS.n2117 VSS.n2107 68.5719
R2019 VSS.n2112 VSS.n2111 68.5719
R2020 VSS.n2090 VSS.n2089 68.5719
R2021 VSS.n2096 VSS.n2095 68.5719
R2022 VSS.n2099 VSS.n2098 68.5719
R2023 VSS.n2179 VSS.n2178 68.5719
R2024 VSS.n2182 VSS.n2060 68.5719
R2025 VSS.n2077 VSS.n2062 68.5719
R2026 VSS.n2071 VSS.n2070 68.5719
R2027 VSS.n1842 VSS.n1841 68.5719
R2028 VSS.n1846 VSS.n1837 68.5719
R2029 VSS.n1847 VSS.n1833 68.5719
R2030 VSS.n13197 VSS.n13196 68.5719
R2031 VSS.n12650 VSS.n12649 68.5719
R2032 VSS.n12653 VSS.n12650 68.5719
R2033 VSS.n12665 VSS.n12655 68.5719
R2034 VSS.n12663 VSS.n12662 68.5719
R2035 VSS.n12660 VSS.n12657 68.5719
R2036 VSS.n2139 VSS.n2138 68.5719
R2037 VSS.n2146 VSS.n2141 68.5719
R2038 VSS.n2143 VSS.n2142 68.5719
R2039 VSS.n13189 VSS.n1856 68.5719
R2040 VSS.n13186 VSS.n1866 68.5719
R2041 VSS.n1876 VSS.n1870 68.5719
R2042 VSS.n1873 VSS.n1871 68.5719
R2043 VSS.n1827 VSS.n1824 68.5719
R2044 VSS.n1825 VSS.n1820 68.5719
R2045 VSS.n13920 VSS.n1817 68.5719
R2046 VSS.n13924 VSS.n13922 68.5719
R2047 VSS.n12688 VSS.n12687 68.5719
R2048 VSS.n12690 VSS.n12685 68.5719
R2049 VSS.n12683 VSS.n12672 68.5719
R2050 VSS.n12679 VSS.n12677 68.5719
R2051 VSS.n1790 VSS.n1786 68.5719
R2052 VSS.n13937 VSS.n1775 68.5719
R2053 VSS.n13934 VSS.n1776 68.5719
R2054 VSS.n13934 VSS.n1792 68.5719
R2055 VSS.n1794 VSS.n1784 68.5719
R2056 VSS.n1808 VSS.n1796 68.5719
R2057 VSS.n1806 VSS.n1805 68.5719
R2058 VSS.n1800 VSS.n1799 68.5719
R2059 VSS.n1959 VSS.n1958 68.5719
R2060 VSS.n1965 VSS.n1956 68.5719
R2061 VSS.n2321 VSS.n1951 68.5719
R2062 VSS.n1967 VSS.n1952 68.5719
R2063 VSS.n2318 VSS.n1974 68.5719
R2064 VSS.n2314 VSS.n2313 68.5719
R2065 VSS.n2310 VSS.n2309 68.5719
R2066 VSS.n2305 VSS.n2304 68.5719
R2067 VSS.n2648 VSS.n2647 68.5719
R2068 VSS.n2654 VSS.n2653 68.5719
R2069 VSS.n2657 VSS.n2656 68.5719
R2070 VSS.n12984 VSS.n12983 68.5719
R2071 VSS.n12987 VSS.n2564 68.5719
R2072 VSS.n2581 VSS.n2566 68.5719
R2073 VSS.n2575 VSS.n2574 68.5719
R2074 VSS.n12965 VSS.n12963 68.5719
R2075 VSS.n12970 VSS.n12958 68.5719
R2076 VSS.n12975 VSS.n12972 68.5719
R2077 VSS.n12973 VSS.n2665 68.5719
R2078 VSS.n2718 VSS.n2717 68.5719
R2079 VSS.n2720 VSS.n2715 68.5719
R2080 VSS.n2713 VSS.n2702 68.5719
R2081 VSS.n2709 VSS.n2707 68.5719
R2082 VSS.n2679 VSS.n2678 68.5719
R2083 VSS.n12951 VSS.n2670 68.5719
R2084 VSS.n2691 VSS.n2672 68.5719
R2085 VSS.n12948 VSS.n2690 68.5719
R2086 VSS.n12943 VSS.n12931 68.5719
R2087 VSS.n12933 VSS.n12932 68.5719
R2088 VSS.n12937 VSS.n12936 68.5719
R2089 VSS.n2776 VSS.n2775 68.5719
R2090 VSS.n2783 VSS.n2772 68.5719
R2091 VSS.n2786 VSS.n2785 68.5719
R2092 VSS.n2817 VSS.n2815 68.5719
R2093 VSS.n2810 VSS.n2809 68.5719
R2094 VSS.n2807 VSS.n2790 68.5719
R2095 VSS.n2798 VSS.n2792 68.5719
R2096 VSS.n2800 VSS.n2797 68.5719
R2097 VSS.n2829 VSS.n2828 68.5719
R2098 VSS.n2835 VSS.n2834 68.5719
R2099 VSS.n2838 VSS.n2837 68.5719
R2100 VSS.n12907 VSS.n12906 68.5719
R2101 VSS.n12910 VSS.n2745 68.5719
R2102 VSS.n2762 VSS.n2747 68.5719
R2103 VSS.n2756 VSS.n2755 68.5719
R2104 VSS.n12888 VSS.n12886 68.5719
R2105 VSS.n12893 VSS.n12881 68.5719
R2106 VSS.n12898 VSS.n12895 68.5719
R2107 VSS.n12896 VSS.n2846 68.5719
R2108 VSS.n2898 VSS.n2897 68.5719
R2109 VSS.n2900 VSS.n2895 68.5719
R2110 VSS.n2893 VSS.n2882 68.5719
R2111 VSS.n2889 VSS.n2887 68.5719
R2112 VSS.n3045 VSS.n3043 68.5719
R2113 VSS.n3049 VSS.n3038 68.5719
R2114 VSS.n3052 VSS.n3051 68.5719
R2115 VSS.n12640 VSS.n12639 68.5719
R2116 VSS.n12634 VSS.n12633 68.5719
R2117 VSS.n12633 VSS.n12632 68.5719
R2118 VSS.n12630 VSS.n3058 68.5719
R2119 VSS.n12624 VSS.n12620 68.5719
R2120 VSS.n12622 VSS.n12621 68.5719
R2121 VSS.n2859 VSS.n2858 68.5719
R2122 VSS.n12874 VSS.n2850 68.5719
R2123 VSS.n2871 VSS.n2852 68.5719
R2124 VSS.n12871 VSS.n2870 68.5719
R2125 VSS.n12866 VSS.n12854 68.5719
R2126 VSS.n12856 VSS.n12855 68.5719
R2127 VSS.n12860 VSS.n12859 68.5719
R2128 VSS.n3032 VSS.n3029 68.5719
R2129 VSS.n3030 VSS.n3025 68.5719
R2130 VSS.n12715 VSS.n3022 68.5719
R2131 VSS.n12719 VSS.n12717 68.5719
R2132 VSS.n3079 VSS.n3078 68.5719
R2133 VSS.n3081 VSS.n3076 68.5719
R2134 VSS.n3074 VSS.n3063 68.5719
R2135 VSS.n3070 VSS.n3068 68.5719
R2136 VSS.n2968 VSS.n2964 68.5719
R2137 VSS.n12732 VSS.n2953 68.5719
R2138 VSS.n12729 VSS.n2954 68.5719
R2139 VSS.n12729 VSS.n2970 68.5719
R2140 VSS.n2972 VSS.n2962 68.5719
R2141 VSS.n3013 VSS.n3001 68.5719
R2142 VSS.n3011 VSS.n3010 68.5719
R2143 VSS.n3005 VSS.n3004 68.5719
R2144 VSS.n2511 VSS.n2510 68.5719
R2145 VSS.n2517 VSS.n2508 68.5719
R2146 VSS.n13026 VSS.n2503 68.5719
R2147 VSS.n2519 VSS.n2504 68.5719
R2148 VSS.n13023 VSS.n2526 68.5719
R2149 VSS.n13019 VSS.n13018 68.5719
R2150 VSS.n13015 VSS.n13014 68.5719
R2151 VSS.n13010 VSS.n13009 68.5719
R2152 VSS.n11321 VSS.n11320 66.4303
R2153 VSS.n8270 VSS.n8266 64.2862
R2154 VSS.n8492 VSS.n8178 64.2862
R2155 VSS.n8374 VSS.n8370 64.2862
R2156 VSS.n8391 VSS.n8210 64.2862
R2157 VSS.n6760 VSS.n6715 64.2862
R2158 VSS.n8024 VSS.n8020 64.2862
R2159 VSS.n8113 VSS.n8095 64.2862
R2160 VSS.n8892 VSS.n7972 64.2862
R2161 VSS.n9583 VSS.n9582 64.2862
R2162 VSS.n9274 VSS.n9004 64.2862
R2163 VSS.n9495 VSS.n9494 64.2862
R2164 VSS.n9471 VSS.n7168 64.2862
R2165 VSS.n9195 VSS.n9194 64.2862
R2166 VSS.n7900 VSS.n7899 64.2862
R2167 VSS.n7626 VSS.n7620 64.2862
R2168 VSS.n7661 VSS.n7655 64.2862
R2169 VSS.n6797 VSS.n6638 64.2862
R2170 VSS.n6865 VSS.n6590 64.2862
R2171 VSS.n6935 VSS.n6934 64.2862
R2172 VSS.n7018 VSS.n6492 64.2862
R2173 VSS.n4180 VSS.n4169 64.2862
R2174 VSS.n938 VSS.n891 64.2862
R2175 VSS.n592 VSS.n588 64.2862
R2176 VSS.n1150 VSS.n933 64.2862
R2177 VSS.n2435 VSS.n2434 64.2862
R2178 VSS.n2341 VSS.n1943 64.2862
R2179 VSS.n1377 VSS.n1376 64.2862
R2180 VSS.n1444 VSS.n638 64.2862
R2181 VSS.n14094 VSS.n14093 64.2862
R2182 VSS.n1656 VSS.n1650 64.2862
R2183 VSS.n1181 VSS.n1177 64.2862
R2184 VSS.n2038 VSS.n1993 64.2862
R2185 VSS.n2087 VSS.n2068 64.2862
R2186 VSS.n2135 VSS.n1862 64.2862
R2187 VSS.n2645 VSS.n2572 64.2862
R2188 VSS.n2683 VSS.n2677 64.2862
R2189 VSS.n2826 VSS.n2753 64.2862
R2190 VSS.n2863 VSS.n2857 64.2862
R2191 VSS.n11414 VSS.n11413 44.424
R2192 VSS.n10529 VSS.n10527 40.4
R2193 VSS.n11499 VSS.n11496 38.9511
R2194 VSS.n11377 VSS.n11376 34.6358
R2195 VSS.n11395 VSS.n11394 34.6358
R2196 VSS.n11252 VSS.n11216 34.6358
R2197 VSS.n3656 VSS.n3644 34.6358
R2198 VSS.n3667 VSS.n3666 34.6358
R2199 VSS.n3672 VSS.n3671 34.6358
R2200 VSS.n11242 VSS.n11241 34.6358
R2201 VSS.n11237 VSS.n11219 34.6358
R2202 VSS.n5110 VSS 34.5605
R2203 VSS.n5112 VSS 34.5605
R2204 VSS.n5119 VSS 34.5605
R2205 VSS.n5117 VSS 34.5605
R2206 VSS.n5138 VSS 34.5605
R2207 VSS.n5145 VSS 34.5605
R2208 VSS.n5152 VSS 34.5605
R2209 VSS.n5159 VSS 34.5605
R2210 VSS.n5179 VSS 34.5605
R2211 VSS.n10169 VSS 34.5605
R2212 VSS.n12297 VSS 34.5605
R2213 VSS.n12308 VSS 34.5605
R2214 VSS.n12514 VSS 34.5605
R2215 VSS.n14487 VSS 34.5605
R2216 VSS.n3319 VSS 34.5605
R2217 VSS.n12527 VSS 34.5605
R2218 VSS.n12525 VSS 34.5605
R2219 VSS.n12523 VSS 34.5605
R2220 VSS.n12521 VSS 34.5605
R2221 VSS.n11255 VSS.n11213 28.9887
R2222 VSS.n11254 VSS.n11253 28.9887
R2223 VSS.n11248 VSS.n11247 28.9887
R2224 VSS.n11246 VSS.n11218 28.9887
R2225 VSS.n3661 VSS.n3660 28.9887
R2226 VSS.n3662 VSS.n3642 28.9887
R2227 VSS.n11312 VSS.n11307 26.9663
R2228 VSS.n11224 VSS.n11221 24.921
R2229 VSS.n11350 VSS.n11349 23.7181
R2230 VSS.n11352 VSS.n3695 23.7181
R2231 VSS.n11359 VSS.n11358 23.7181
R2232 VSS.n11413 VSS.n3686 23.7181
R2233 VSS.n11260 VSS.n11259 23.7181
R2234 VSS.n3647 VSS.n3639 23.7181
R2235 VSS.n11282 VSS.n11281 23.4463
R2236 VSS.n11310 VSS.n11309 23.4463
R2237 VSS.n11358 VSS.n3693 22.2123
R2238 VSS.n11264 VSS.n11263 20.3989
R2239 VSS.n11301 VSS.n11298 19.3944
R2240 VSS.n3636 VSS.n3633 19.3944
R2241 VSS.n11271 VSS.n11203 19.0674
R2242 VSS.n10632 VSS 18.3101
R2243 VSS VSS.n10628 18.3101
R2244 VSS.n11230 VSS.n11227 17.7168
R2245 VSS.n11424 VSS.n11420 17.7168
R2246 VSS.n11425 VSS.n11424 17.7168
R2247 VSS.n10529 VSS.n10528 17.6755
R2248 VSS.n11482 VSS.n11478 17.649
R2249 VSS.n3671 VSS.n3641 17.3181
R2250 VSS.n3675 VSS.n3640 17.3181
R2251 VSS.n11238 VSS.n11237 17.3181
R2252 VSS.n11233 VSS.n11232 17.3181
R2253 VSS VSS.n4543 17.3181
R2254 VSS VSS.n10600 17.3181
R2255 VSS.n4550 VSS 17.3181
R2256 VSS.n10200 VSS 17.3181
R2257 VSS.n10417 VSS 17.3181
R2258 VSS.n10418 VSS 17.3181
R2259 VSS VSS.n4861 17.3181
R2260 VSS VSS.n4860 17.3181
R2261 VSS VSS.n4824 17.3181
R2262 VSS.n4927 VSS 17.3181
R2263 VSS.n4815 VSS 17.3181
R2264 VSS.n4816 VSS 17.3181
R2265 VSS.n4818 VSS 17.3181
R2266 VSS VSS.n4817 17.3181
R2267 VSS.n5099 VSS 17.3181
R2268 VSS VSS.n5098 17.3181
R2269 VSS VSS.n5095 17.3181
R2270 VSS.n4948 VSS 17.3181
R2271 VSS.n4943 VSS 17.3181
R2272 VSS VSS.n4946 17.3181
R2273 VSS.n4935 VSS 17.3181
R2274 VSS.n4934 VSS 17.3181
R2275 VSS VSS.n4834 17.3181
R2276 VSS VSS.n4835 17.3181
R2277 VSS VSS.n4841 17.3181
R2278 VSS VSS.n4842 17.3181
R2279 VSS VSS.n4852 17.3181
R2280 VSS VSS.n4853 17.3181
R2281 VSS VSS.n4862 17.3181
R2282 VSS VSS.n4863 17.3181
R2283 VSS.n4907 VSS 17.3181
R2284 VSS.n4906 VSS 17.3181
R2285 VSS.n4905 VSS 17.3181
R2286 VSS VSS.n4549 17.3181
R2287 VSS.n10193 VSS 17.3181
R2288 VSS.n10192 VSS 17.3181
R2289 VSS VSS.n4552 17.3181
R2290 VSS VSS.n10177 17.3181
R2291 VSS.n5106 VSS 17.3181
R2292 VSS VSS.n5109 17.3181
R2293 VSS.n10174 VSS 17.3181
R2294 VSS.n10175 VSS 17.3181
R2295 VSS.n10392 VSS 17.3181
R2296 VSS VSS.n10391 17.3181
R2297 VSS VSS.n10389 17.3181
R2298 VSS.n10385 VSS 17.3181
R2299 VSS VSS.n10383 17.3181
R2300 VSS.n10380 VSS 17.3181
R2301 VSS VSS.n10378 17.3181
R2302 VSS.n10375 VSS 17.3181
R2303 VSS.n10374 VSS 17.3181
R2304 VSS.n10373 VSS 17.3181
R2305 VSS.n10594 VSS 17.3181
R2306 VSS.n10593 VSS 17.3181
R2307 VSS VSS.n11443 17.3181
R2308 VSS.n11444 VSS 17.3181
R2309 VSS.n12491 VSS 17.3181
R2310 VSS.n12490 VSS 17.3181
R2311 VSS.n12481 VSS 17.3181
R2312 VSS.n12483 VSS 17.3181
R2313 VSS.n10425 VSS 17.3181
R2314 VSS.n10424 VSS 17.3181
R2315 VSS.n10422 VSS 17.3181
R2316 VSS.n10421 VSS 17.3181
R2317 VSS.n10415 VSS 17.3181
R2318 VSS.n10414 VSS 17.3181
R2319 VSS.n10413 VSS 17.3181
R2320 VSS.n10412 VSS 17.3181
R2321 VSS VSS.n10507 17.3181
R2322 VSS.n10508 VSS 17.3181
R2323 VSS VSS.n10513 17.3181
R2324 VSS.n10514 VSS 17.3181
R2325 VSS.n10519 VSS 17.3181
R2326 VSS VSS.n10523 17.3181
R2327 VSS.n10532 VSS 17.3181
R2328 VSS.n10531 VSS 17.3181
R2329 VSS.n11432 VSS 17.3181
R2330 VSS.n11431 VSS 17.3181
R2331 VSS.n11451 VSS 17.3181
R2332 VSS.n11450 VSS 17.3181
R2333 VSS VSS.n11449 17.3181
R2334 VSS.n3681 VSS 17.3181
R2335 VSS.n11438 VSS 17.3181
R2336 VSS.n10203 VSS 17.3181
R2337 VSS.n10604 VSS 17.3181
R2338 VSS.n10605 VSS 17.3181
R2339 VSS VSS.n4706 17.2429
R2340 VSS VSS.n12550 17.2429
R2341 VSS.n11455 VSS.n3676 16.8752
R2342 VSS.n11483 VSS.n11482 16.2614
R2343 VSS.n3637 VSS.n3636 15.952
R2344 VSS.n11302 VSS.n11301 15.7581
R2345 VSS.n11255 VSS.n11254 15.4358
R2346 VSS.n11253 VSS 15.4358
R2347 VSS.n11247 VSS.n11246 15.4358
R2348 VSS VSS.n3655 15.4358
R2349 VSS.n3662 VSS.n3661 15.4358
R2350 VSS.n3642 VSS 15.4358
R2351 VSS VSS.n11218 15.4358
R2352 VSS.n11290 VSS.n11203 14.4975
R2353 VSS.n11231 VSS.n11224 14.395
R2354 VSS.n11317 VSS.n11315 14.2324
R2355 VSS.n3695 VSS.n3694 12.8005
R2356 VSS.n11456 VSS.n11455 12.2814
R2357 VSS.n11259 VSS.n11213 9.78874
R2358 VSS.n11248 VSS.n11216 9.78874
R2359 VSS.n3660 VSS.n3644 9.78874
R2360 VSS.n5096 VSS.n4746 8.65932
R2361 VSS VSS.n4746 8.65932
R2362 VSS.n4940 VSS 8.65932
R2363 VSS.n4942 VSS.n4941 8.65932
R2364 VSS.n4941 VSS 8.65932
R2365 VSS.n4950 VSS.n4949 8.65932
R2366 VSS.n4950 VSS 8.65932
R2367 VSS.n4954 VSS.n4807 8.65932
R2368 VSS VSS.n4954 8.65932
R2369 VSS.n5088 VSS 8.65932
R2370 VSS.n4956 VSS.n4955 8.65932
R2371 VSS.n4955 VSS 8.65932
R2372 VSS.n4806 VSS.n4805 8.65932
R2373 VSS.n4805 VSS 8.65932
R2374 VSS.n4957 VSS 8.65932
R2375 VSS.n4810 VSS.n4803 8.65932
R2376 VSS VSS.n4803 8.65932
R2377 VSS.n4962 VSS.n4800 8.65932
R2378 VSS VSS.n4962 8.65932
R2379 VSS VSS.n4939 8.65932
R2380 VSS.n4938 VSS.n4936 8.65932
R2381 VSS VSS.n4938 8.65932
R2382 VSS.n4933 VSS.n4932 8.65932
R2383 VSS.n4932 VSS 8.65932
R2384 VSS VSS.n4830 8.65932
R2385 VSS.n4829 VSS.n4827 8.65932
R2386 VSS VSS.n4829 8.65932
R2387 VSS.n4931 VSS.n4930 8.65932
R2388 VSS.n4930 VSS 8.65932
R2389 VSS VSS.n4964 8.65932
R2390 VSS.n4967 VSS.n4965 8.65932
R2391 VSS.n4967 VSS 8.65932
R2392 VSS.n5016 VSS 8.65932
R2393 VSS.n4975 VSS.n4973 8.65932
R2394 VSS VSS.n4975 8.65932
R2395 VSS.n4966 VSS.n4798 8.65932
R2396 VSS VSS.n4798 8.65932
R2397 VSS VSS.n4972 8.65932
R2398 VSS.n4797 VSS.n4796 8.65932
R2399 VSS.n4796 VSS 8.65932
R2400 VSS.n4795 VSS.n4752 8.65932
R2401 VSS VSS.n4752 8.65932
R2402 VSS.n5082 VSS.n5081 8.65932
R2403 VSS.n5081 VSS 8.65932
R2404 VSS.n5080 VSS.n5079 8.65932
R2405 VSS.n5079 VSS 8.65932
R2406 VSS.n4985 VSS.n4984 8.65932
R2407 VSS.n4984 VSS 8.65932
R2408 VSS.n5000 VSS 8.65932
R2409 VSS.n5002 VSS.n5001 8.65932
R2410 VSS.n5001 VSS 8.65932
R2411 VSS VSS.n4977 8.65932
R2412 VSS.n5078 VSS.n4755 8.65932
R2413 VSS VSS.n4755 8.65932
R2414 VSS.n5077 VSS.n5076 8.65932
R2415 VSS.n5076 VSS 8.65932
R2416 VSS.n5010 VSS 8.65932
R2417 VSS.n5012 VSS.n5011 8.65932
R2418 VSS.n5011 VSS 8.65932
R2419 VSS.n5015 VSS.n5014 8.65932
R2420 VSS.n5014 VSS 8.65932
R2421 VSS VSS.n4787 8.65932
R2422 VSS.n4826 VSS.n4786 8.65932
R2423 VSS VSS.n4786 8.65932
R2424 VSS.n5023 VSS.n4783 8.65932
R2425 VSS VSS.n5023 8.65932
R2426 VSS.n4831 VSS 8.65932
R2427 VSS.n4833 VSS.n4832 8.65932
R2428 VSS.n4832 VSS 8.65932
R2429 VSS.n4840 VSS.n4839 8.65932
R2430 VSS.n4839 VSS 8.65932
R2431 VSS.n4849 VSS 8.65932
R2432 VSS.n4851 VSS.n4850 8.65932
R2433 VSS.n4850 VSS 8.65932
R2434 VSS.n4859 VSS.n4858 8.65932
R2435 VSS.n4858 VSS 8.65932
R2436 VSS.n4857 VSS.n4856 8.65932
R2437 VSS.n4856 VSS 8.65932
R2438 VSS.n4893 VSS 8.65932
R2439 VSS.n4892 VSS.n4890 8.65932
R2440 VSS VSS.n4892 8.65932
R2441 VSS.n5058 VSS.n5057 8.65932
R2442 VSS.n5058 VSS 8.65932
R2443 VSS VSS.n5056 8.65932
R2444 VSS.n5054 VSS.n4775 8.65932
R2445 VSS VSS.n5054 8.65932
R2446 VSS.n4844 VSS.n4778 8.65932
R2447 VSS VSS.n4778 8.65932
R2448 VSS VSS.n4848 8.65932
R2449 VSS.n4847 VSS.n4845 8.65932
R2450 VSS VSS.n4847 8.65932
R2451 VSS.n4838 VSS 8.65932
R2452 VSS VSS.n5025 8.65932
R2453 VSS.n5028 VSS.n5026 8.65932
R2454 VSS.n5028 VSS 8.65932
R2455 VSS.n5036 VSS.n5034 8.65932
R2456 VSS VSS.n5036 8.65932
R2457 VSS.n5027 VSS.n4781 8.65932
R2458 VSS VSS.n4781 8.65932
R2459 VSS VSS.n5033 8.65932
R2460 VSS.n4991 VSS.n4780 8.65932
R2461 VSS.n4991 VSS 8.65932
R2462 VSS.n4990 VSS.n4759 8.65932
R2463 VSS VSS.n4759 8.65932
R2464 VSS.n5074 VSS.n5073 8.65932
R2465 VSS.n5073 VSS 8.65932
R2466 VSS.n5072 VSS.n5071 8.65932
R2467 VSS.n5071 VSS 8.65932
R2468 VSS.n5172 VSS.n5171 8.65932
R2469 VSS.n5172 VSS 8.65932
R2470 VSS VSS.n5170 8.65932
R2471 VSS.n5167 VSS.n5166 8.65932
R2472 VSS.n5167 VSS 8.65932
R2473 VSS VSS.n5165 8.65932
R2474 VSS.n5070 VSS.n4762 8.65932
R2475 VSS.n4762 VSS 8.65932
R2476 VSS.n5069 VSS.n5068 8.65932
R2477 VSS.n5068 VSS 8.65932
R2478 VSS.n5040 VSS 8.65932
R2479 VSS.n5042 VSS.n5041 8.65932
R2480 VSS.n5041 VSS 8.65932
R2481 VSS.n5047 VSS 8.65932
R2482 VSS VSS.n4779 8.65932
R2483 VSS.n5046 VSS.n5045 8.65932
R2484 VSS.n5045 VSS 8.65932
R2485 VSS.n4771 VSS.n4770 8.65932
R2486 VSS.n4770 VSS 8.65932
R2487 VSS VSS.n5066 8.65932
R2488 VSS.n5063 VSS.n5062 8.65932
R2489 VSS.n5063 VSS 8.65932
R2490 VSS.n5044 VSS.n4773 8.65932
R2491 VSS VSS.n4773 8.65932
R2492 VSS VSS.n5061 8.65932
R2493 VSS.n4871 VSS.n4772 8.65932
R2494 VSS.n4871 VSS 8.65932
R2495 VSS.n4878 VSS.n4868 8.65932
R2496 VSS VSS.n4878 8.65932
R2497 VSS.n4883 VSS.n4882 8.65932
R2498 VSS.n4882 VSS 8.65932
R2499 VSS.n4874 VSS.n4867 8.65932
R2500 VSS.n4874 VSS 8.65932
R2501 VSS.n4884 VSS 8.65932
R2502 VSS.n4886 VSS.n4885 8.65932
R2503 VSS.n4885 VSS 8.65932
R2504 VSS.n4899 VSS.n4898 8.65932
R2505 VSS.n4899 VSS 8.65932
R2506 VSS VSS.n4897 8.65932
R2507 VSS.n4888 VSS.n4887 8.65932
R2508 VSS.n4888 VSS 8.65932
R2509 VSS VSS.n4904 8.65932
R2510 VSS.n4873 VSS 8.65932
R2511 VSS VSS.n10191 8.65932
R2512 VSS.n10190 VSS.n4553 8.65932
R2513 VSS VSS.n10190 8.65932
R2514 VSS.n4881 VSS 8.65932
R2515 VSS.n10186 VSS 8.65932
R2516 VSS.n10185 VSS.n10184 8.65932
R2517 VSS.n10184 VSS 8.65932
R2518 VSS.n10183 VSS.n10182 8.65932
R2519 VSS.n10182 VSS 8.65932
R2520 VSS.n10181 VSS.n10180 8.65932
R2521 VSS.n10180 VSS 8.65932
R2522 VSS.n10179 VSS.n10178 8.65932
R2523 VSS.n10178 VSS 8.65932
R2524 VSS.n10165 VSS.n4558 8.65932
R2525 VSS VSS.n10165 8.65932
R2526 VSS.n4724 VSS 8.65932
R2527 VSS.n4726 VSS.n4725 8.65932
R2528 VSS.n4725 VSS 8.65932
R2529 VSS.n4767 VSS 8.65932
R2530 VSS.n4769 VSS.n4768 8.65932
R2531 VSS.n4768 VSS 8.65932
R2532 VSS.n5067 VSS 8.65932
R2533 VSS.n5161 VSS.n4727 8.65932
R2534 VSS.n5161 VSS 8.65932
R2535 VSS.n4987 VSS 8.65932
R2536 VSS.n4989 VSS.n4988 8.65932
R2537 VSS.n4988 VSS 8.65932
R2538 VSS VSS.n4999 8.65932
R2539 VSS.n4995 VSS.n4758 8.65932
R2540 VSS.n4995 VSS 8.65932
R2541 VSS.n5075 VSS 8.65932
R2542 VSS.n4981 VSS.n4980 8.65932
R2543 VSS.n4980 VSS 8.65932
R2544 VSS.n5003 VSS 8.65932
R2545 VSS.n4979 VSS.n4740 8.65932
R2546 VSS VSS.n4979 8.65932
R2547 VSS.n4789 VSS 8.65932
R2548 VSS.n4788 VSS.n4751 8.65932
R2549 VSS VSS.n4788 8.65932
R2550 VSS.n5083 VSS 8.65932
R2551 VSS.n5085 VSS.n5084 8.65932
R2552 VSS.n5084 VSS 8.65932
R2553 VSS.n5132 VSS.n5131 8.65932
R2554 VSS.n5132 VSS 8.65932
R2555 VSS VSS.n5130 8.65932
R2556 VSS.n5128 VSS.n5126 8.65932
R2557 VSS VSS.n5128 8.65932
R2558 VSS VSS.n5125 8.65932
R2559 VSS.n5087 VSS.n5086 8.65932
R2560 VSS.n5086 VSS 8.65932
R2561 VSS VSS.n4747 8.65932
R2562 VSS.n5121 VSS.n4741 8.65932
R2563 VSS.n5121 VSS 8.65932
R2564 VSS.n5103 VSS 8.65932
R2565 VSS.n5105 VSS.n5104 8.65932
R2566 VSS.n5104 VSS 8.65932
R2567 VSS.n5120 VSS 8.65932
R2568 VSS VSS.n5137 8.65932
R2569 VSS VSS.n5144 8.65932
R2570 VSS VSS.n5151 8.65932
R2571 VSS.n5160 VSS 8.65932
R2572 VSS VSS.n4719 8.65932
R2573 VSS VSS.n10168 8.65932
R2574 VSS.n10390 VSS.n10273 8.65932
R2575 VSS.n10273 VSS 8.65932
R2576 VSS.n10384 VSS.n10275 8.65932
R2577 VSS.n10275 VSS 8.65932
R2578 VSS.n10379 VSS.n10370 8.65932
R2579 VSS.n10370 VSS 8.65932
R2580 VSS.n10592 VSS.n10591 8.65932
R2581 VSS.n10591 VSS 8.65932
R2582 VSS VSS.n10363 8.65932
R2583 VSS.n10280 VSS.n3679 8.65932
R2584 VSS.n10280 VSS 8.65932
R2585 VSS VSS.n12495 8.65932
R2586 VSS.n12494 VSS.n12492 8.65932
R2587 VSS VSS.n12494 8.65932
R2588 VSS.n12489 VSS.n12488 8.65932
R2589 VSS.n12488 VSS 8.65932
R2590 VSS.n12487 VSS.n12486 8.65932
R2591 VSS.n12486 VSS 8.65932
R2592 VSS.n12301 VSS.n12299 8.65932
R2593 VSS VSS.n12301 8.65932
R2594 VSS.n12307 VSS.n12302 8.65932
R2595 VSS VSS.n12307 8.65932
R2596 VSS VSS.n12513 8.65932
R2597 VSS.n12509 VSS.n12508 8.65932
R2598 VSS.n12509 VSS 8.65932
R2599 VSS VSS.n12507 8.65932
R2600 VSS.n12504 VSS.n12503 8.65932
R2601 VSS.n12504 VSS 8.65932
R2602 VSS VSS.n12502 8.65932
R2603 VSS.n12500 VSS.n3598 8.65932
R2604 VSS VSS.n12500 8.65932
R2605 VSS.n10303 VSS.n3601 8.65932
R2606 VSS VSS.n10303 8.65932
R2607 VSS.n12496 VSS 8.65932
R2608 VSS.n10359 VSS.n10279 8.65932
R2609 VSS.n10359 VSS 8.65932
R2610 VSS.n10357 VSS.n10278 8.65932
R2611 VSS.n10357 VSS 8.65932
R2612 VSS.n10364 VSS 8.65932
R2613 VSS.n10365 VSS.n10207 8.65932
R2614 VSS.n10365 VSS 8.65932
R2615 VSS.n10590 VSS 8.65932
R2616 VSS VSS.n10208 8.65932
R2617 VSS.n10589 VSS.n10588 8.65932
R2618 VSS.n10588 VSS 8.65932
R2619 VSS.n10286 VSS.n10211 8.65932
R2620 VSS.n10286 VSS 8.65932
R2621 VSS.n10587 VSS.n10586 8.65932
R2622 VSS.n10586 VSS 8.65932
R2623 VSS VSS.n10212 8.65932
R2624 VSS.n10585 VSS.n10584 8.65932
R2625 VSS.n10584 VSS 8.65932
R2626 VSS VSS.n10296 8.65932
R2627 VSS.n10295 VSS.n10215 8.65932
R2628 VSS VSS.n10295 8.65932
R2629 VSS.n10583 VSS.n10582 8.65932
R2630 VSS.n10582 VSS 8.65932
R2631 VSS VSS.n10216 8.65932
R2632 VSS.n10581 VSS.n10580 8.65932
R2633 VSS.n10580 VSS 8.65932
R2634 VSS.n10579 VSS.n10578 8.65932
R2635 VSS.n10578 VSS 8.65932
R2636 VSS.n10575 VSS 8.65932
R2637 VSS.n10577 VSS.n10576 8.65932
R2638 VSS.n10576 VSS 8.65932
R2639 VSS.n10432 VSS.n10270 8.65932
R2640 VSS VSS.n10432 8.65932
R2641 VSS.n10428 VSS 8.65932
R2642 VSS.n10427 VSS.n10426 8.65932
R2643 VSS VSS.n10427 8.65932
R2644 VSS.n10423 VSS.n10399 8.65932
R2645 VSS.n10399 VSS 8.65932
R2646 VSS.n10420 VSS.n10419 8.65932
R2647 VSS.n10419 VSS 8.65932
R2648 VSS.n10463 VSS.n10266 8.65932
R2649 VSS.n10463 VSS 8.65932
R2650 VSS.n10496 VSS.n10258 8.65932
R2651 VSS.n10496 VSS 8.65932
R2652 VSS.n10460 VSS 8.65932
R2653 VSS.n10462 VSS.n10461 8.65932
R2654 VSS.n10461 VSS 8.65932
R2655 VSS.n10467 VSS.n10262 8.65932
R2656 VSS VSS.n10467 8.65932
R2657 VSS VSS.n10459 8.65932
R2658 VSS.n10458 VSS.n10267 8.65932
R2659 VSS VSS.n10458 8.65932
R2660 VSS.n10398 VSS 8.65932
R2661 VSS VSS.n10433 8.65932
R2662 VSS.n10435 VSS.n10434 8.65932
R2663 VSS VSS.n10435 8.65932
R2664 VSS.n10453 VSS.n10436 8.65932
R2665 VSS.n10453 VSS 8.65932
R2666 VSS.n10452 VSS.n10438 8.65932
R2667 VSS.n10438 VSS 8.65932
R2668 VSS.n10451 VSS.n10450 8.65932
R2669 VSS.n10450 VSS 8.65932
R2670 VSS.n10441 VSS 8.65932
R2671 VSS.n10440 VSS.n10221 8.65932
R2672 VSS VSS.n10440 8.65932
R2673 VSS.n10325 VSS.n10222 8.65932
R2674 VSS.n10325 VSS 8.65932
R2675 VSS VSS.n10574 8.65932
R2676 VSS.n10571 VSS.n10223 8.65932
R2677 VSS VSS.n10571 8.65932
R2678 VSS.n10567 VSS.n10226 8.65932
R2679 VSS.n10567 VSS 8.65932
R2680 VSS.n10297 VSS 8.65932
R2681 VSS.n10298 VSS.n10290 8.65932
R2682 VSS.n10298 VSS 8.65932
R2683 VSS VSS.n10289 8.65932
R2684 VSS.n10356 VSS 8.65932
R2685 VSS.n10355 VSS.n10354 8.65932
R2686 VSS.n10354 VSS 8.65932
R2687 VSS.n10353 VSS.n10352 8.65932
R2688 VSS.n10352 VSS 8.65932
R2689 VSS.n10351 VSS.n10350 8.65932
R2690 VSS.n10350 VSS 8.65932
R2691 VSS.n10340 VSS.n10339 8.65932
R2692 VSS.n10339 VSS 8.65932
R2693 VSS VSS.n10314 8.65932
R2694 VSS.n10313 VSS.n10228 8.65932
R2695 VSS VSS.n10313 8.65932
R2696 VSS.n10349 VSS.n10348 8.65932
R2697 VSS.n10348 VSS 8.65932
R2698 VSS.n10566 VSS 8.65932
R2699 VSS.n10565 VSS.n10564 8.65932
R2700 VSS.n10564 VSS 8.65932
R2701 VSS VSS.n10337 8.65932
R2702 VSS.n10329 VSS.n10231 8.65932
R2703 VSS.n10329 VSS 8.65932
R2704 VSS.n10563 VSS.n10562 8.65932
R2705 VSS.n10562 VSS 8.65932
R2706 VSS VSS.n10232 8.65932
R2707 VSS.n10561 VSS.n10560 8.65932
R2708 VSS.n10560 VSS 8.65932
R2709 VSS.n10444 VSS 8.65932
R2710 VSS.n10445 VSS.n10235 8.65932
R2711 VSS.n10445 VSS 8.65932
R2712 VSS.n10559 VSS.n10558 8.65932
R2713 VSS.n10558 VSS 8.65932
R2714 VSS VSS.n10236 8.65932
R2715 VSS.n10557 VSS.n10556 8.65932
R2716 VSS.n10556 VSS 8.65932
R2717 VSS.n10555 VSS.n10554 8.65932
R2718 VSS.n10554 VSS 8.65932
R2719 VSS.n10471 VSS 8.65932
R2720 VSS.n10553 VSS.n10239 8.65932
R2721 VSS VSS.n10239 8.65932
R2722 VSS.n10552 VSS.n10551 8.65932
R2723 VSS.n10551 VSS 8.65932
R2724 VSS.n10470 VSS 8.65932
R2725 VSS.n10480 VSS.n10261 8.65932
R2726 VSS VSS.n10261 8.65932
R2727 VSS VSS.n10479 8.65932
R2728 VSS.n10468 VSS 8.65932
R2729 VSS.n10482 VSS.n10481 8.65932
R2730 VSS.n10482 VSS 8.65932
R2731 VSS.n10492 VSS.n10491 8.65932
R2732 VSS.n10491 VSS 8.65932
R2733 VSS.n10485 VSS.n10260 8.65932
R2734 VSS VSS.n10485 8.65932
R2735 VSS.n10495 VSS 8.65932
R2736 VSS.n10494 VSS.n10493 8.65932
R2737 VSS.n10493 VSS 8.65932
R2738 VSS.n10251 VSS.n10242 8.65932
R2739 VSS.n10251 VSS 8.65932
R2740 VSS.n10490 VSS 8.65932
R2741 VSS.n10550 VSS 8.65932
R2742 VSS.n10549 VSS.n10548 8.65932
R2743 VSS.n10548 VSS 8.65932
R2744 VSS.n10547 VSS.n10546 8.65932
R2745 VSS.n10546 VSS 8.65932
R2746 VSS.n10545 VSS.n10534 8.65932
R2747 VSS.n10534 VSS 8.65932
R2748 VSS.n10544 VSS.n10543 8.65932
R2749 VSS.n10543 VSS 8.65932
R2750 VSS VSS.n10248 8.65932
R2751 VSS.n10245 VSS.n3376 8.65932
R2752 VSS.n10245 VSS 8.65932
R2753 VSS.n12544 VSS.n12543 8.65932
R2754 VSS.n12544 VSS 8.65932
R2755 VSS VSS.n12542 8.65932
R2756 VSS.n12540 VSS.n12538 8.65932
R2757 VSS VSS.n12540 8.65932
R2758 VSS.n12537 VSS.n3377 8.65932
R2759 VSS VSS.n3377 8.65932
R2760 VSS VSS.n12536 8.65932
R2761 VSS.n10324 VSS.n10323 8.65932
R2762 VSS.n10323 VSS 8.65932
R2763 VSS.n10331 VSS.n10321 8.65932
R2764 VSS.n10331 VSS 8.65932
R2765 VSS.n10338 VSS 8.65932
R2766 VSS.n10502 VSS.n10501 8.65932
R2767 VSS VSS.n10502 8.65932
R2768 VSS VSS.n10500 8.65932
R2769 VSS.n10416 VSS.n10406 8.65932
R2770 VSS.n10406 VSS 8.65932
R2771 VSS.n10503 VSS 8.65932
R2772 VSS VSS.n10512 8.65932
R2773 VSS VSS.n10518 8.65932
R2774 VSS.n10533 VSS 8.65932
R2775 VSS.n10542 VSS 8.65932
R2776 VSS VSS.n3321 8.65932
R2777 VSS VSS.n3379 8.65932
R2778 VSS VSS.n3587 8.65932
R2779 VSS VSS.n12520 8.65932
R2780 VSS.n10318 VSS.n10317 8.65932
R2781 VSS.n10317 VSS 8.65932
R2782 VSS.n10341 VSS 8.65932
R2783 VSS.n10316 VSS.n3596 8.65932
R2784 VSS VSS.n10316 8.65932
R2785 VSS.n10308 VSS 8.65932
R2786 VSS.n10309 VSS.n10306 8.65932
R2787 VSS.n10309 VSS 8.65932
R2788 VSS.n10304 VSS 8.65932
R2789 VSS.n11434 VSS.n11433 8.65932
R2790 VSS.n11434 VSS 8.65932
R2791 VSS VSS.n11437 8.65932
R2792 VSS.n10601 VSS 8.65932
R2793 VSS.n10603 VSS.n10602 8.65932
R2794 VSS.n10602 VSS 8.65932
R2795 VSS.n13589 VSS.n13588 8.53383
R2796 VSS.n13588 VSS.n13507 8.53383
R2797 VSS.n13600 VSS.n13507 8.53383
R2798 VSS.n13600 VSS.n13599 8.53383
R2799 VSS.n13599 VSS.n13509 8.53383
R2800 VSS.n13596 VSS.n13509 8.53383
R2801 VSS.n13596 VSS.n13595 8.53383
R2802 VSS.n13595 VSS.n13592 8.53383
R2803 VSS.n1763 VSS.n1762 8.53383
R2804 VSS.n1762 VSS.n1742 8.53383
R2805 VSS.n14013 VSS.n1742 8.53383
R2806 VSS.n14013 VSS.n14012 8.53383
R2807 VSS.n14012 VSS.n1744 8.53383
R2808 VSS.n14009 VSS.n1744 8.53383
R2809 VSS.n14009 VSS.n14008 8.53383
R2810 VSS.n14008 VSS.n14005 8.53383
R2811 VSS.n2931 VSS.n2930 8.53383
R2812 VSS.n12800 VSS.n2931 8.53383
R2813 VSS.n12800 VSS.n12799 8.53383
R2814 VSS.n12799 VSS.n2933 8.53383
R2815 VSS.n12793 VSS.n2933 8.53383
R2816 VSS.n12793 VSS.n12792 8.53383
R2817 VSS.n12792 VSS.n12789 8.53383
R2818 VSS.n12790 VSS.n12789 8.53383
R2819 VSS.n2880 VSS.n2842 8.53383
R2820 VSS.n2901 VSS.n2880 8.53383
R2821 VSS.n2901 VSS.n2881 8.53383
R2822 VSS.n2892 VSS.n2881 8.53383
R2823 VSS.n2892 VSS.n2891 8.53383
R2824 VSS.n2891 VSS.n2890 8.53383
R2825 VSS.n2890 VSS.n2883 8.53383
R2826 VSS.n2885 VSS.n2883 8.53383
R2827 VSS.n2811 VSS.n2788 8.53383
R2828 VSS.n2806 VSS.n2788 8.53383
R2829 VSS.n2806 VSS.n2805 8.53383
R2830 VSS.n2805 VSS.n2804 8.53383
R2831 VSS.n2804 VSS.n2793 8.53383
R2832 VSS.n2801 VSS.n2793 8.53383
R2833 VSS.n2801 VSS.n2795 8.53383
R2834 VSS.n2795 VSS.n2794 8.53383
R2835 VSS.n3894 VSS.n3893 8.53383
R2836 VSS.n10895 VSS.n3894 8.53383
R2837 VSS.n10895 VSS.n10894 8.53383
R2838 VSS.n10894 VSS.n3896 8.53383
R2839 VSS.n10888 VSS.n3896 8.53383
R2840 VSS.n10888 VSS.n10887 8.53383
R2841 VSS.n10887 VSS.n10884 8.53383
R2842 VSS.n10885 VSS.n10884 8.53383
R2843 VSS.n10942 VSS.n10920 8.53383
R2844 VSS.n10940 VSS.n10920 8.53383
R2845 VSS.n10940 VSS.n10939 8.53383
R2846 VSS.n10939 VSS.n10924 8.53383
R2847 VSS.n10925 VSS.n10924 8.53383
R2848 VSS.n10932 VSS.n10925 8.53383
R2849 VSS.n10932 VSS.n10927 8.53383
R2850 VSS.n10930 VSS.n10927 8.53383
R2851 VSS.n3826 VSS.n3825 8.53383
R2852 VSS.n11046 VSS.n3826 8.53383
R2853 VSS.n11046 VSS.n11045 8.53383
R2854 VSS.n11045 VSS.n3828 8.53383
R2855 VSS.n11039 VSS.n3828 8.53383
R2856 VSS.n11039 VSS.n11038 8.53383
R2857 VSS.n11038 VSS.n11035 8.53383
R2858 VSS.n11036 VSS.n11035 8.53383
R2859 VSS.n6562 VSS.n6561 8.53383
R2860 VSS.n6984 VSS.n6562 8.53383
R2861 VSS.n6984 VSS.n6563 8.53383
R2862 VSS.n6575 VSS.n6563 8.53383
R2863 VSS.n6575 VSS.n6574 8.53383
R2864 VSS.n6574 VSS.n6573 8.53383
R2865 VSS.n6573 VSS.n6568 8.53383
R2866 VSS.n6569 VSS.n6568 8.53383
R2867 VSS.n9562 VSS.n7566 8.53383
R2868 VSS.n9564 VSS.n7566 8.53383
R2869 VSS.n9567 VSS.n9564 8.53383
R2870 VSS.n9570 VSS.n9567 8.53383
R2871 VSS.n9570 VSS.n7564 8.53383
R2872 VSS.n9573 VSS.n7564 8.53383
R2873 VSS.n9574 VSS.n9573 8.53383
R2874 VSS.n9574 VSS.n7562 8.53383
R2875 VSS.n8496 VSS.n8493 8.53383
R2876 VSS.n8499 VSS.n8496 8.53383
R2877 VSS.n8500 VSS.n8499 8.53383
R2878 VSS.n8503 VSS.n8500 8.53383
R2879 VSS.n8507 VSS.n8503 8.53383
R2880 VSS.n8507 VSS.n8504 8.53383
R2881 VSS.n8504 VSS.n8185 8.53383
R2882 VSS.n8373 VSS.n8369 8.53383
R2883 VSS.n8378 VSS.n8369 8.53383
R2884 VSS.n8379 VSS.n8378 8.53383
R2885 VSS.n8379 VSS.n8366 8.53383
R2886 VSS.n8387 VSS.n8366 8.53383
R2887 VSS.n8387 VSS.n8367 8.53383
R2888 VSS.n8367 VSS.n8187 8.53383
R2889 VSS.n8395 VSS.n8392 8.53383
R2890 VSS.n8398 VSS.n8395 8.53383
R2891 VSS.n8399 VSS.n8398 8.53383
R2892 VSS.n8402 VSS.n8399 8.53383
R2893 VSS.n8406 VSS.n8402 8.53383
R2894 VSS.n8406 VSS.n8403 8.53383
R2895 VSS.n8403 VSS.n8217 8.53383
R2896 VSS.n8252 VSS.n8251 8.53383
R2897 VSS.n8252 VSS.n8247 8.53383
R2898 VSS.n8259 VSS.n8247 8.53383
R2899 VSS.n8259 VSS.n8245 8.53383
R2900 VSS.n8773 VSS.n8245 8.53383
R2901 VSS.n8774 VSS.n8773 8.53383
R2902 VSS.n8774 VSS.n8219 8.53383
R2903 VSS.n8220 VSS.n8218 8.53383
R2904 VSS.n8238 VSS.n8220 8.53383
R2905 VSS.n8238 VSS.n8236 8.53383
R2906 VSS.n8236 VSS.n8235 8.53383
R2907 VSS.n8235 VSS.n8222 8.53383
R2908 VSS.n8230 VSS.n8222 8.53383
R2909 VSS.n8230 VSS.n8226 8.53383
R2910 VSS.n8228 VSS.n8226 8.53383
R2911 VSS.n8195 VSS.n8194 8.53383
R2912 VSS.n8792 VSS.n8195 8.53383
R2913 VSS.n8792 VSS.n8791 8.53383
R2914 VSS.n8791 VSS.n8197 8.53383
R2915 VSS.n8206 VSS.n8197 8.53383
R2916 VSS.n8206 VSS.n8205 8.53383
R2917 VSS.n8205 VSS.n8202 8.53383
R2918 VSS.n8203 VSS.n8202 8.53383
R2919 VSS.n6214 VSS.n6213 8.53383
R2920 VSS.n9981 VSS.n6214 8.53383
R2921 VSS.n9981 VSS.n6215 8.53383
R2922 VSS.n6221 VSS.n6215 8.53383
R2923 VSS.n6224 VSS.n6221 8.53383
R2924 VSS.n6226 VSS.n6224 8.53383
R2925 VSS.n6227 VSS.n6226 8.53383
R2926 VSS.n6227 VSS.n6219 8.53383
R2927 VSS.n6757 VSS.n6716 8.53383
R2928 VSS.n6757 VSS.n6754 8.53383
R2929 VSS.n6754 VSS.n6753 8.53383
R2930 VSS.n6753 VSS.n6750 8.53383
R2931 VSS.n6750 VSS.n6749 8.53383
R2932 VSS.n6749 VSS.n6718 8.53383
R2933 VSS.n6745 VSS.n6718 8.53383
R2934 VSS.n6693 VSS.n6692 8.53383
R2935 VSS.n6765 VSS.n6693 8.53383
R2936 VSS.n6765 VSS.n6694 8.53383
R2937 VSS.n6701 VSS.n6694 8.53383
R2938 VSS.n6707 VSS.n6701 8.53383
R2939 VSS.n6707 VSS.n6706 8.53383
R2940 VSS.n6706 VSS.n6703 8.53383
R2941 VSS.n6704 VSS.n6703 8.53383
R2942 VSS.n9961 VSS.n9956 8.53383
R2943 VSS.n9961 VSS.n9954 8.53383
R2944 VSS.n9964 VSS.n9954 8.53383
R2945 VSS.n9964 VSS.n9952 8.53383
R2946 VSS.n9970 VSS.n9952 8.53383
R2947 VSS.n9970 VSS.n6233 8.53383
R2948 VSS.n9972 VSS.n6233 8.53383
R2949 VSS.n8029 VSS.n8025 8.53383
R2950 VSS.n8030 VSS.n8029 8.53383
R2951 VSS.n8031 VSS.n8030 8.53383
R2952 VSS.n8031 VSS.n8017 8.53383
R2953 VSS.n8155 VSS.n8017 8.53383
R2954 VSS.n8155 VSS.n8018 8.53383
R2955 VSS.n8018 VSS.n8016 8.53383
R2956 VSS.n8110 VSS.n8096 8.53383
R2957 VSS.n8110 VSS.n8107 8.53383
R2958 VSS.n8107 VSS.n8106 8.53383
R2959 VSS.n8106 VSS.n8103 8.53383
R2960 VSS.n8103 VSS.n8102 8.53383
R2961 VSS.n8102 VSS.n8098 8.53383
R2962 VSS.n8098 VSS.n8037 8.53383
R2963 VSS.n8047 VSS.n8036 8.53383
R2964 VSS.n8089 VSS.n8047 8.53383
R2965 VSS.n8089 VSS.n8048 8.53383
R2966 VSS.n8085 VSS.n8048 8.53383
R2967 VSS.n8085 VSS.n8082 8.53383
R2968 VSS.n8082 VSS.n8081 8.53383
R2969 VSS.n8081 VSS.n8078 8.53383
R2970 VSS.n8078 VSS.n8077 8.53383
R2971 VSS.n8147 VSS.n8119 8.53383
R2972 VSS.n8145 VSS.n8119 8.53383
R2973 VSS.n8145 VSS.n8144 8.53383
R2974 VSS.n8144 VSS.n8129 8.53383
R2975 VSS.n8139 VSS.n8129 8.53383
R2976 VSS.n8139 VSS.n8138 8.53383
R2977 VSS.n8138 VSS.n8131 8.53383
R2978 VSS.n8134 VSS.n8131 8.53383
R2979 VSS.n8051 VSS.n8001 8.53383
R2980 VSS.n8072 VSS.n8051 8.53383
R2981 VSS.n8072 VSS.n8052 8.53383
R2982 VSS.n8063 VSS.n8052 8.53383
R2983 VSS.n8063 VSS.n8062 8.53383
R2984 VSS.n8062 VSS.n8061 8.53383
R2985 VSS.n8061 VSS.n8054 8.53383
R2986 VSS.n8056 VSS.n8054 8.53383
R2987 VSS.n8889 VSS.n7973 8.53383
R2988 VSS.n8889 VSS.n8886 8.53383
R2989 VSS.n8886 VSS.n8885 8.53383
R2990 VSS.n8885 VSS.n8882 8.53383
R2991 VSS.n8882 VSS.n8881 8.53383
R2992 VSS.n8881 VSS.n7975 8.53383
R2993 VSS.n8877 VSS.n7975 8.53383
R2994 VSS.n7949 VSS.n7948 8.53383
R2995 VSS.n8897 VSS.n7949 8.53383
R2996 VSS.n8897 VSS.n7950 8.53383
R2997 VSS.n7958 VSS.n7950 8.53383
R2998 VSS.n7964 VSS.n7958 8.53383
R2999 VSS.n7964 VSS.n7963 8.53383
R3000 VSS.n7963 VSS.n7960 8.53383
R3001 VSS.n7961 VSS.n7960 8.53383
R3002 VSS.n8856 VSS.n8852 8.53383
R3003 VSS.n8856 VSS.n8006 8.53383
R3004 VSS.n8862 VSS.n8006 8.53383
R3005 VSS.n8863 VSS.n8862 8.53383
R3006 VSS.n8864 VSS.n8863 8.53383
R3007 VSS.n8864 VSS.n8003 8.53383
R3008 VSS.n8870 VSS.n8003 8.53383
R3009 VSS.n8190 VSS.n8186 8.53383
R3010 VSS.n8812 VSS.n8190 8.53383
R3011 VSS.n8812 VSS.n8192 8.53383
R3012 VSS.n8808 VSS.n8192 8.53383
R3013 VSS.n8808 VSS.n8797 8.53383
R3014 VSS.n8803 VSS.n8797 8.53383
R3015 VSS.n8803 VSS.n8802 8.53383
R3016 VSS.n8802 VSS.n8801 8.53383
R3017 VSS.n8163 VSS.n8162 8.53383
R3018 VSS.n8830 VSS.n8163 8.53383
R3019 VSS.n8830 VSS.n8829 8.53383
R3020 VSS.n8829 VSS.n8165 8.53383
R3021 VSS.n8174 VSS.n8165 8.53383
R3022 VSS.n8174 VSS.n8173 8.53383
R3023 VSS.n8173 VSS.n8170 8.53383
R3024 VSS.n8171 VSS.n8170 8.53383
R3025 VSS.n7571 VSS.n7567 8.53383
R3026 VSS.n9550 VSS.n7571 8.53383
R3027 VSS.n9550 VSS.n7573 8.53383
R3028 VSS.n7586 VSS.n7573 8.53383
R3029 VSS.n7586 VSS.n7585 8.53383
R3030 VSS.n7585 VSS.n7577 8.53383
R3031 VSS.n7578 VSS.n7577 8.53383
R3032 VSS.n7579 VSS.n7578 8.53383
R3033 VSS.n8269 VSS.n8265 8.53383
R3034 VSS.n8274 VSS.n8265 8.53383
R3035 VSS.n8275 VSS.n8274 8.53383
R3036 VSS.n8275 VSS.n8262 8.53383
R3037 VSS.n8283 VSS.n8262 8.53383
R3038 VSS.n8283 VSS.n8263 8.53383
R3039 VSS.n8263 VSS.n7568 8.53383
R3040 VSS.n9586 VSS.n9580 8.53383
R3041 VSS.n9587 VSS.n9586 8.53383
R3042 VSS.n9587 VSS.n9578 8.53383
R3043 VSS.n9578 VSS.n7552 8.53383
R3044 VSS.n9594 VSS.n7552 8.53383
R3045 VSS.n9594 VSS.n7553 8.53383
R3046 VSS.n7553 VSS.n7551 8.53383
R3047 VSS.n9312 VSS.n9291 8.53383
R3048 VSS.n9312 VSS.n9311 8.53383
R3049 VSS.n9311 VSS.n9293 8.53383
R3050 VSS.n9306 VSS.n9293 8.53383
R3051 VSS.n9306 VSS.n9296 8.53383
R3052 VSS.n9303 VSS.n9296 8.53383
R3053 VSS.n9303 VSS.n9298 8.53383
R3054 VSS.n9298 VSS.n9297 8.53383
R3055 VSS.n8995 VSS.n8994 8.53383
R3056 VSS.n9520 VSS.n8995 8.53383
R3057 VSS.n9520 VSS.n9519 8.53383
R3058 VSS.n9519 VSS.n8997 8.53383
R3059 VSS.n9012 VSS.n8997 8.53383
R3060 VSS.n9012 VSS.n9011 8.53383
R3061 VSS.n9011 VSS.n9008 8.53383
R3062 VSS.n9009 VSS.n9008 8.53383
R3063 VSS.n9278 VSS.n9275 8.53383
R3064 VSS.n9278 VSS.n9272 8.53383
R3065 VSS.n9281 VSS.n9272 8.53383
R3066 VSS.n9284 VSS.n9281 8.53383
R3067 VSS.n9287 VSS.n9284 8.53383
R3068 VSS.n9287 VSS.n9018 8.53383
R3069 VSS.n9290 VSS.n9018 8.53383
R3070 VSS.n9499 VSS.n9492 8.53383
R3071 VSS.n9500 VSS.n9499 8.53383
R3072 VSS.n9500 VSS.n9490 8.53383
R3073 VSS.n9490 VSS.n9488 8.53383
R3074 VSS.n9507 VSS.n9488 8.53383
R3075 VSS.n9507 VSS.n9317 8.53383
R3076 VSS.n9509 VSS.n9317 8.53383
R3077 VSS.n7223 VSS.n7184 8.53383
R3078 VSS.n7224 VSS.n7223 8.53383
R3079 VSS.n7224 VSS.n7218 8.53383
R3080 VSS.n7238 VSS.n7218 8.53383
R3081 VSS.n7238 VSS.n7219 8.53383
R3082 VSS.n7228 VSS.n7219 8.53383
R3083 VSS.n7231 VSS.n7228 8.53383
R3084 VSS.n7231 VSS.n7230 8.53383
R3085 VSS.n7159 VSS.n7158 8.53383
R3086 VSS.n9842 VSS.n7159 8.53383
R3087 VSS.n9842 VSS.n9841 8.53383
R3088 VSS.n9841 VSS.n7161 8.53383
R3089 VSS.n7176 VSS.n7161 8.53383
R3090 VSS.n7176 VSS.n7175 8.53383
R3091 VSS.n7175 VSS.n7172 8.53383
R3092 VSS.n7173 VSS.n7172 8.53383
R3093 VSS.n9473 VSS.n9472 8.53383
R3094 VSS.n9476 VSS.n9473 8.53383
R3095 VSS.n9484 VSS.n9476 8.53383
R3096 VSS.n9484 VSS.n9483 8.53383
R3097 VSS.n9483 VSS.n9481 8.53383
R3098 VSS.n9481 VSS.n9480 8.53383
R3099 VSS.n9480 VSS.n7183 8.53383
R3100 VSS.n9831 VSS.n7186 8.53383
R3101 VSS.n9819 VSS.n9814 8.53383
R3102 VSS.n9819 VSS.n9812 8.53383
R3103 VSS.n9822 VSS.n9812 8.53383
R3104 VSS.n9822 VSS.n9810 8.53383
R3105 VSS.n9829 VSS.n9810 8.53383
R3106 VSS.n9829 VSS.n7186 8.53383
R3107 VSS.n7260 VSS.n7210 8.53383
R3108 VSS.n7255 VSS.n7210 8.53383
R3109 VSS.n7255 VSS.n7254 8.53383
R3110 VSS.n7254 VSS.n7253 8.53383
R3111 VSS.n7253 VSS.n7215 8.53383
R3112 VSS.n7250 VSS.n7215 8.53383
R3113 VSS.n7250 VSS.n7244 8.53383
R3114 VSS.n7244 VSS.n7243 8.53383
R3115 VSS.n7357 VSS.n7354 8.53383
R3116 VSS.n7358 VSS.n7357 8.53383
R3117 VSS.n7361 VSS.n7358 8.53383
R3118 VSS.n7361 VSS.n7277 8.53383
R3119 VSS.n7365 VSS.n7277 8.53383
R3120 VSS.n7365 VSS.n7278 8.53383
R3121 VSS.n7278 VSS.n7262 8.53383
R3122 VSS.n7314 VSS.n7261 8.53383
R3123 VSS.n7315 VSS.n7314 8.53383
R3124 VSS.n7318 VSS.n7315 8.53383
R3125 VSS.n7327 VSS.n7318 8.53383
R3126 VSS.n7327 VSS.n7324 8.53383
R3127 VSS.n7324 VSS.n7323 8.53383
R3128 VSS.n7323 VSS.n7322 8.53383
R3129 VSS.n7322 VSS.n7320 8.53383
R3130 VSS.n7203 VSS.n7198 8.53383
R3131 VSS.n7204 VSS.n7203 8.53383
R3132 VSS.n7205 VSS.n7204 8.53383
R3133 VSS.n7205 VSS.n7191 8.53383
R3134 VSS.n7378 VSS.n7191 8.53383
R3135 VSS.n7378 VSS.n7377 8.53383
R3136 VSS.n7377 VSS.n7190 8.53383
R3137 VSS.n9162 VSS.n9160 8.53383
R3138 VSS.n9177 VSS.n9172 8.53383
R3139 VSS.n9178 VSS.n9177 8.53383
R3140 VSS.n9179 VSS.n9178 8.53383
R3141 VSS.n9179 VSS.n9161 8.53383
R3142 VSS.n9268 VSS.n9161 8.53383
R3143 VSS.n9268 VSS.n9162 8.53383
R3144 VSS.n9215 VSS.n9187 8.53383
R3145 VSS.n9236 VSS.n9215 8.53383
R3146 VSS.n9236 VSS.n9217 8.53383
R3147 VSS.n9230 VSS.n9217 8.53383
R3148 VSS.n9230 VSS.n9229 8.53383
R3149 VSS.n9229 VSS.n9221 8.53383
R3150 VSS.n9222 VSS.n9221 8.53383
R3151 VSS.n9223 VSS.n9222 8.53383
R3152 VSS.n9199 VSS.n9192 8.53383
R3153 VSS.n9200 VSS.n9199 8.53383
R3154 VSS.n9200 VSS.n9190 8.53383
R3155 VSS.n9206 VSS.n9190 8.53383
R3156 VSS.n9208 VSS.n9206 8.53383
R3157 VSS.n9209 VSS.n9208 8.53383
R3158 VSS.n9209 VSS.n9188 8.53383
R3159 VSS.n9262 VSS.n9246 8.53383
R3160 VSS.n9262 VSS.n9261 8.53383
R3161 VSS.n9261 VSS.n9259 8.53383
R3162 VSS.n9259 VSS.n9257 8.53383
R3163 VSS.n9257 VSS.n9247 8.53383
R3164 VSS.n9252 VSS.n9247 8.53383
R3165 VSS.n9252 VSS.n9249 8.53383
R3166 VSS.n9249 VSS.n9248 8.53383
R3167 VSS.n7849 VSS.n7847 8.53383
R3168 VSS.n7847 VSS.n7846 8.53383
R3169 VSS.n7846 VSS.n7810 8.53383
R3170 VSS.n8961 VSS.n7810 8.53383
R3171 VSS.n8961 VSS.n7811 8.53383
R3172 VSS.n7821 VSS.n7811 8.53383
R3173 VSS.n7823 VSS.n7821 8.53383
R3174 VSS.n7823 VSS.n7822 8.53383
R3175 VSS.n7854 VSS.n7850 8.53383
R3176 VSS.n8943 VSS.n7854 8.53383
R3177 VSS.n8943 VSS.n7856 8.53383
R3178 VSS.n7869 VSS.n7856 8.53383
R3179 VSS.n7869 VSS.n7868 8.53383
R3180 VSS.n7868 VSS.n7860 8.53383
R3181 VSS.n7861 VSS.n7860 8.53383
R3182 VSS.n7862 VSS.n7861 8.53383
R3183 VSS.n7902 VSS.n7901 8.53383
R3184 VSS.n7902 VSS.n7896 8.53383
R3185 VSS.n7916 VSS.n7896 8.53383
R3186 VSS.n7916 VSS.n7915 8.53383
R3187 VSS.n7915 VSS.n7907 8.53383
R3188 VSS.n7908 VSS.n7907 8.53383
R3189 VSS.n7908 VSS.n7851 8.53383
R3190 VSS.n8955 VSS.n8954 8.53383
R3191 VSS.n7836 VSS.n7833 8.53383
R3192 VSS.n7836 VSS.n7831 8.53383
R3193 VSS.n7841 VSS.n7831 8.53383
R3194 VSS.n7843 VSS.n7841 8.53383
R3195 VSS.n7844 VSS.n7843 8.53383
R3196 VSS.n8955 VSS.n7844 8.53383
R3197 VSS.n7736 VSS.n7640 8.53383
R3198 VSS.n7737 VSS.n7736 8.53383
R3199 VSS.n7737 VSS.n7731 8.53383
R3200 VSS.n7751 VSS.n7731 8.53383
R3201 VSS.n7751 VSS.n7732 8.53383
R3202 VSS.n7741 VSS.n7732 8.53383
R3203 VSS.n7744 VSS.n7741 8.53383
R3204 VSS.n7744 VSS.n7743 8.53383
R3205 VSS.n8983 VSS.n7807 8.53383
R3206 VSS.n8981 VSS.n7807 8.53383
R3207 VSS.n8981 VSS.n8980 8.53383
R3208 VSS.n8980 VSS.n8978 8.53383
R3209 VSS.n8978 VSS.n8970 8.53383
R3210 VSS.n8975 VSS.n8970 8.53383
R3211 VSS.n8975 VSS.n8974 8.53383
R3212 VSS.n8974 VSS.n8971 8.53383
R3213 VSS.n7624 VSS.n7623 8.53383
R3214 VSS.n7623 VSS.n7612 8.53383
R3215 VSS.n8989 VSS.n7612 8.53383
R3216 VSS.n8989 VSS.n8988 8.53383
R3217 VSS.n8988 VSS.n7614 8.53383
R3218 VSS.n7635 VSS.n7614 8.53383
R3219 VSS.n7636 VSS.n7635 8.53383
R3220 VSS.n7804 VSS.n7642 8.53383
R3221 VSS.n7792 VSS.n7787 8.53383
R3222 VSS.n7792 VSS.n7785 8.53383
R3223 VSS.n7795 VSS.n7785 8.53383
R3224 VSS.n7795 VSS.n7783 8.53383
R3225 VSS.n7802 VSS.n7783 8.53383
R3226 VSS.n7802 VSS.n7642 8.53383
R3227 VSS.n7696 VSS.n7675 8.53383
R3228 VSS.n7696 VSS.n7695 8.53383
R3229 VSS.n7695 VSS.n7693 8.53383
R3230 VSS.n7693 VSS.n7677 8.53383
R3231 VSS.n7688 VSS.n7677 8.53383
R3232 VSS.n7688 VSS.n7687 8.53383
R3233 VSS.n7687 VSS.n7680 8.53383
R3234 VSS.n7685 VSS.n7680 8.53383
R3235 VSS.n7773 VSS.n7728 8.53383
R3236 VSS.n7771 VSS.n7728 8.53383
R3237 VSS.n7771 VSS.n7770 8.53383
R3238 VSS.n7770 VSS.n7768 8.53383
R3239 VSS.n7768 VSS.n7760 8.53383
R3240 VSS.n7765 VSS.n7760 8.53383
R3241 VSS.n7765 VSS.n7764 8.53383
R3242 VSS.n7764 VSS.n7761 8.53383
R3243 VSS.n7659 VSS.n7658 8.53383
R3244 VSS.n7658 VSS.n7647 8.53383
R3245 VSS.n7779 VSS.n7647 8.53383
R3246 VSS.n7779 VSS.n7778 8.53383
R3247 VSS.n7778 VSS.n7649 8.53383
R3248 VSS.n7670 VSS.n7649 8.53383
R3249 VSS.n7671 VSS.n7670 8.53383
R3250 VSS.n7725 VSS.n7701 8.53383
R3251 VSS.n7713 VSS.n7708 8.53383
R3252 VSS.n7713 VSS.n7706 8.53383
R3253 VSS.n7716 VSS.n7706 8.53383
R3254 VSS.n7716 VSS.n7704 8.53383
R3255 VSS.n7723 VSS.n7704 8.53383
R3256 VSS.n7723 VSS.n7701 8.53383
R3257 VSS.n7071 VSS.n7070 8.53383
R3258 VSS.n9896 VSS.n7071 8.53383
R3259 VSS.n9896 VSS.n7072 8.53383
R3260 VSS.n7078 VSS.n7072 8.53383
R3261 VSS.n7081 VSS.n7078 8.53383
R3262 VSS.n7083 VSS.n7081 8.53383
R3263 VSS.n7084 VSS.n7083 8.53383
R3264 VSS.n7084 VSS.n7076 8.53383
R3265 VSS.n7126 VSS.n7123 8.53383
R3266 VSS.n7126 VSS.n7121 8.53383
R3267 VSS.n7131 VSS.n7121 8.53383
R3268 VSS.n7132 VSS.n7131 8.53383
R3269 VSS.n7135 VSS.n7132 8.53383
R3270 VSS.n7135 VSS.n7133 8.53383
R3271 VSS.n7133 VSS.n7089 8.53383
R3272 VSS.n7099 VSS.n7088 8.53383
R3273 VSS.n7113 VSS.n7099 8.53383
R3274 VSS.n7113 VSS.n7111 8.53383
R3275 VSS.n7111 VSS.n7110 8.53383
R3276 VSS.n7110 VSS.n7100 8.53383
R3277 VSS.n7105 VSS.n7100 8.53383
R3278 VSS.n7105 VSS.n7104 8.53383
R3279 VSS.n7104 VSS.n7101 8.53383
R3280 VSS.n9876 VSS.n9871 8.53383
R3281 VSS.n9876 VSS.n9869 8.53383
R3282 VSS.n9879 VSS.n9869 8.53383
R3283 VSS.n9879 VSS.n9867 8.53383
R3284 VSS.n9885 VSS.n9867 8.53383
R3285 VSS.n9885 VSS.n7144 8.53383
R3286 VSS.n9887 VSS.n7144 8.53383
R3287 VSS.n7939 VSS.n7893 8.53383
R3288 VSS.n7926 VSS.n7923 8.53383
R3289 VSS.n7926 VSS.n7921 8.53383
R3290 VSS.n7931 VSS.n7921 8.53383
R3291 VSS.n7932 VSS.n7931 8.53383
R3292 VSS.n7935 VSS.n7932 8.53383
R3293 VSS.n7935 VSS.n7893 8.53383
R3294 VSS.n7944 VSS.n7940 8.53383
R3295 VSS.n8918 VSS.n7944 8.53383
R3296 VSS.n8918 VSS.n7946 8.53383
R3297 VSS.n8914 VSS.n7946 8.53383
R3298 VSS.n8914 VSS.n8903 8.53383
R3299 VSS.n8909 VSS.n8903 8.53383
R3300 VSS.n8909 VSS.n8908 8.53383
R3301 VSS.n8908 VSS.n8907 8.53383
R3302 VSS.n7987 VSS.n7980 8.53383
R3303 VSS.n7988 VSS.n7987 8.53383
R3304 VSS.n7989 VSS.n7988 8.53383
R3305 VSS.n7989 VSS.n7977 8.53383
R3306 VSS.n7997 VSS.n7977 8.53383
R3307 VSS.n7997 VSS.n7978 8.53383
R3308 VSS.n7978 VSS.n7941 8.53383
R3309 VSS.n7873 VSS.n7872 8.53383
R3310 VSS.n8936 VSS.n7873 8.53383
R3311 VSS.n8936 VSS.n8935 8.53383
R3312 VSS.n8935 VSS.n7875 8.53383
R3313 VSS.n7885 VSS.n7875 8.53383
R3314 VSS.n7885 VSS.n7884 8.53383
R3315 VSS.n7884 VSS.n7881 8.53383
R3316 VSS.n7882 VSS.n7881 8.53383
R3317 VSS.n6610 VSS.n6609 8.53383
R3318 VSS.n6911 VSS.n6610 8.53383
R3319 VSS.n6911 VSS.n6611 8.53383
R3320 VSS.n6623 VSS.n6611 8.53383
R3321 VSS.n6623 VSS.n6622 8.53383
R3322 VSS.n6622 VSS.n6621 8.53383
R3323 VSS.n6621 VSS.n6616 8.53383
R3324 VSS.n6617 VSS.n6616 8.53383
R3325 VSS.n6643 VSS.n6628 8.53383
R3326 VSS.n6851 VSS.n6643 8.53383
R3327 VSS.n6851 VSS.n6644 8.53383
R3328 VSS.n6654 VSS.n6644 8.53383
R3329 VSS.n6654 VSS.n6653 8.53383
R3330 VSS.n6653 VSS.n6651 8.53383
R3331 VSS.n6651 VSS.n6650 8.53383
R3332 VSS.n6650 VSS.n6648 8.53383
R3333 VSS.n6799 VSS.n6798 8.53383
R3334 VSS.n6802 VSS.n6799 8.53383
R3335 VSS.n6810 VSS.n6802 8.53383
R3336 VSS.n6810 VSS.n6809 8.53383
R3337 VSS.n6809 VSS.n6807 8.53383
R3338 VSS.n6807 VSS.n6806 8.53383
R3339 VSS.n6806 VSS.n6629 8.53383
R3340 VSS.n6891 VSS.n6886 8.53383
R3341 VSS.n6891 VSS.n6884 8.53383
R3342 VSS.n6894 VSS.n6884 8.53383
R3343 VSS.n6894 VSS.n6882 8.53383
R3344 VSS.n6901 VSS.n6882 8.53383
R3345 VSS.n6901 VSS.n6859 8.53383
R3346 VSS.n6903 VSS.n6859 8.53383
R3347 VSS.n6595 VSS.n6580 8.53383
R3348 VSS.n6918 VSS.n6595 8.53383
R3349 VSS.n6918 VSS.n6596 8.53383
R3350 VSS.n6606 VSS.n6596 8.53383
R3351 VSS.n6606 VSS.n6605 8.53383
R3352 VSS.n6605 VSS.n6603 8.53383
R3353 VSS.n6603 VSS.n6602 8.53383
R3354 VSS.n6602 VSS.n6600 8.53383
R3355 VSS.n6867 VSS.n6866 8.53383
R3356 VSS.n6870 VSS.n6867 8.53383
R3357 VSS.n6878 VSS.n6870 8.53383
R3358 VSS.n6878 VSS.n6877 8.53383
R3359 VSS.n6877 VSS.n6875 8.53383
R3360 VSS.n6875 VSS.n6874 8.53383
R3361 VSS.n6874 VSS.n6581 8.53383
R3362 VSS.n6964 VSS.n6959 8.53383
R3363 VSS.n6964 VSS.n6957 8.53383
R3364 VSS.n6967 VSS.n6957 8.53383
R3365 VSS.n6967 VSS.n6955 8.53383
R3366 VSS.n6974 VSS.n6955 8.53383
R3367 VSS.n6974 VSS.n6926 8.53383
R3368 VSS.n6976 VSS.n6926 8.53383
R3369 VSS.n6538 VSS.n6536 8.53383
R3370 VSS.n6536 VSS.n6535 8.53383
R3371 VSS.n6535 VSS.n6512 8.53383
R3372 VSS.n7043 VSS.n6512 8.53383
R3373 VSS.n7043 VSS.n6513 8.53383
R3374 VSS.n6523 VSS.n6513 8.53383
R3375 VSS.n6525 VSS.n6523 8.53383
R3376 VSS.n6525 VSS.n6524 8.53383
R3377 VSS.n6543 VSS.n6539 8.53383
R3378 VSS.n6991 VSS.n6543 8.53383
R3379 VSS.n6991 VSS.n6545 8.53383
R3380 VSS.n6558 VSS.n6545 8.53383
R3381 VSS.n6558 VSS.n6557 8.53383
R3382 VSS.n6557 VSS.n6549 8.53383
R3383 VSS.n6550 VSS.n6549 8.53383
R3384 VSS.n6551 VSS.n6550 8.53383
R3385 VSS.n6937 VSS.n6936 8.53383
R3386 VSS.n6937 VSS.n6931 8.53383
R3387 VSS.n6951 VSS.n6931 8.53383
R3388 VSS.n6951 VSS.n6950 8.53383
R3389 VSS.n6950 VSS.n6942 8.53383
R3390 VSS.n6943 VSS.n6942 8.53383
R3391 VSS.n6943 VSS.n6540 8.53383
R3392 VSS.n7037 VSS.n7036 8.53383
R3393 VSS.n7006 VSS.n7003 8.53383
R3394 VSS.n7007 VSS.n7006 8.53383
R3395 VSS.n7012 VSS.n7007 8.53383
R3396 VSS.n7012 VSS.n7009 8.53383
R3397 VSS.n7009 VSS.n6533 8.53383
R3398 VSS.n7037 VSS.n6533 8.53383
R3399 VSS.n6481 VSS.n6291 8.53383
R3400 VSS.n6293 VSS.n6291 8.53383
R3401 VSS.n6475 VSS.n6293 8.53383
R3402 VSS.n6475 VSS.n6474 8.53383
R3403 VSS.n6474 VSS.n6295 8.53383
R3404 VSS.n6471 VSS.n6295 8.53383
R3405 VSS.n6471 VSS.n6464 8.53383
R3406 VSS.n6464 VSS.n6463 8.53383
R3407 VSS.n6497 VSS.n6482 8.53383
R3408 VSS.n7050 VSS.n6497 8.53383
R3409 VSS.n7050 VSS.n6498 8.53383
R3410 VSS.n6508 VSS.n6498 8.53383
R3411 VSS.n6508 VSS.n6507 8.53383
R3412 VSS.n6507 VSS.n6505 8.53383
R3413 VSS.n6505 VSS.n6504 8.53383
R3414 VSS.n6504 VSS.n6502 8.53383
R3415 VSS.n7020 VSS.n7019 8.53383
R3416 VSS.n7023 VSS.n7020 8.53383
R3417 VSS.n7031 VSS.n7023 8.53383
R3418 VSS.n7031 VSS.n7030 8.53383
R3419 VSS.n7030 VSS.n7028 8.53383
R3420 VSS.n7028 VSS.n7027 8.53383
R3421 VSS.n7027 VSS.n6483 8.53383
R3422 VSS.n7063 VSS.n6271 8.53383
R3423 VSS.n6283 VSS.n6278 8.53383
R3424 VSS.n6284 VSS.n6283 8.53383
R3425 VSS.n6285 VSS.n6284 8.53383
R3426 VSS.n6285 VSS.n6272 8.53383
R3427 VSS.n7064 VSS.n6272 8.53383
R3428 VSS.n7064 VSS.n7063 8.53383
R3429 VSS.n6298 VSS.n6297 8.53383
R3430 VSS.n6458 VSS.n6298 8.53383
R3431 VSS.n6458 VSS.n6299 8.53383
R3432 VSS.n6305 VSS.n6299 8.53383
R3433 VSS.n6308 VSS.n6305 8.53383
R3434 VSS.n6310 VSS.n6308 8.53383
R3435 VSS.n6311 VSS.n6310 8.53383
R3436 VSS.n6311 VSS.n6303 8.53383
R3437 VSS.n6411 VSS.n6408 8.53383
R3438 VSS.n6412 VSS.n6411 8.53383
R3439 VSS.n6415 VSS.n6412 8.53383
R3440 VSS.n6415 VSS.n6331 8.53383
R3441 VSS.n6419 VSS.n6331 8.53383
R3442 VSS.n6419 VSS.n6332 8.53383
R3443 VSS.n6332 VSS.n6316 8.53383
R3444 VSS.n6368 VSS.n6315 8.53383
R3445 VSS.n6369 VSS.n6368 8.53383
R3446 VSS.n6372 VSS.n6369 8.53383
R3447 VSS.n6381 VSS.n6372 8.53383
R3448 VSS.n6381 VSS.n6378 8.53383
R3449 VSS.n6378 VSS.n6377 8.53383
R3450 VSS.n6377 VSS.n6376 8.53383
R3451 VSS.n6376 VSS.n6374 8.53383
R3452 VSS.n6438 VSS.n6433 8.53383
R3453 VSS.n6438 VSS.n6431 8.53383
R3454 VSS.n6441 VSS.n6431 8.53383
R3455 VSS.n6441 VSS.n6429 8.53383
R3456 VSS.n6447 VSS.n6429 8.53383
R3457 VSS.n6447 VSS.n6428 8.53383
R3458 VSS.n6449 VSS.n6428 8.53383
R3459 VSS.n6835 VSS.n6793 8.53383
R3460 VSS.n6824 VSS.n6819 8.53383
R3461 VSS.n6824 VSS.n6817 8.53383
R3462 VSS.n6827 VSS.n6817 8.53383
R3463 VSS.n6827 VSS.n6815 8.53383
R3464 VSS.n6833 VSS.n6815 8.53383
R3465 VSS.n6833 VSS.n6793 8.53383
R3466 VSS.n6689 VSS.n6675 8.53383
R3467 VSS.n6783 VSS.n6689 8.53383
R3468 VSS.n6783 VSS.n6690 8.53383
R3469 VSS.n6779 VSS.n6690 8.53383
R3470 VSS.n6779 VSS.n6776 8.53383
R3471 VSS.n6776 VSS.n6775 8.53383
R3472 VSS.n6775 VSS.n6772 8.53383
R3473 VSS.n6772 VSS.n6771 8.53383
R3474 VSS.n6725 VSS.n6720 8.53383
R3475 VSS.n6726 VSS.n6725 8.53383
R3476 VSS.n6729 VSS.n6726 8.53383
R3477 VSS.n6730 VSS.n6729 8.53383
R3478 VSS.n6735 VSS.n6730 8.53383
R3479 VSS.n6735 VSS.n6732 8.53383
R3480 VSS.n6732 VSS.n6676 8.53383
R3481 VSS.n6658 VSS.n6657 8.53383
R3482 VSS.n6844 VSS.n6658 8.53383
R3483 VSS.n6844 VSS.n6659 8.53383
R3484 VSS.n6671 VSS.n6659 8.53383
R3485 VSS.n6671 VSS.n6670 8.53383
R3486 VSS.n6670 VSS.n6669 8.53383
R3487 VSS.n6669 VSS.n6664 8.53383
R3488 VSS.n6665 VSS.n6664 8.53383
R3489 VSS.n6388 VSS.n6347 8.53383
R3490 VSS.n6388 VSS.n6387 8.53383
R3491 VSS.n6387 VSS.n6350 8.53383
R3492 VSS.n6364 VSS.n6350 8.53383
R3493 VSS.n6364 VSS.n6363 8.53383
R3494 VSS.n6363 VSS.n6355 8.53383
R3495 VSS.n6358 VSS.n6355 8.53383
R3496 VSS.n6358 VSS.n6357 8.53383
R3497 VSS.n6340 VSS.n6339 8.53383
R3498 VSS.n6340 VSS.n6335 8.53383
R3499 VSS.n6403 VSS.n6335 8.53383
R3500 VSS.n6403 VSS.n6402 8.53383
R3501 VSS.n6402 VSS.n6345 8.53383
R3502 VSS.n6396 VSS.n6345 8.53383
R3503 VSS.n6396 VSS.n6395 8.53383
R3504 VSS.n11025 VSS.n3839 8.53383
R3505 VSS.n11015 VSS.n11012 8.53383
R3506 VSS.n11015 VSS.n11010 8.53383
R3507 VSS.n11018 VSS.n11010 8.53383
R3508 VSS.n11020 VSS.n11018 8.53383
R3509 VSS.n11023 VSS.n11020 8.53383
R3510 VSS.n11023 VSS.n3839 8.53383
R3511 VSS.n3854 VSS.n3853 8.53383
R3512 VSS.n10991 VSS.n3854 8.53383
R3513 VSS.n10991 VSS.n10990 8.53383
R3514 VSS.n10990 VSS.n3856 8.53383
R3515 VSS.n3867 VSS.n3856 8.53383
R3516 VSS.n3869 VSS.n3867 8.53383
R3517 VSS.n3870 VSS.n3869 8.53383
R3518 VSS.n3870 VSS.n3864 8.53383
R3519 VSS.n10975 VSS.n10972 8.53383
R3520 VSS.n10975 VSS.n10968 8.53383
R3521 VSS.n10978 VSS.n10968 8.53383
R3522 VSS.n10979 VSS.n10978 8.53383
R3523 VSS.n10982 VSS.n10979 8.53383
R3524 VSS.n10982 VSS.n3879 8.53383
R3525 VSS.n10984 VSS.n3879 8.53383
R3526 VSS.n10950 VSS.n10900 8.53383
R3527 VSS.n10910 VSS.n10903 8.53383
R3528 VSS.n10911 VSS.n10910 8.53383
R3529 VSS.n10912 VSS.n10911 8.53383
R3530 VSS.n10912 VSS.n10901 8.53383
R3531 VSS.n10951 VSS.n10901 8.53383
R3532 VSS.n10951 VSS.n10950 8.53383
R3533 VSS.n7334 VSS.n7293 8.53383
R3534 VSS.n7334 VSS.n7333 8.53383
R3535 VSS.n7333 VSS.n7296 8.53383
R3536 VSS.n7310 VSS.n7296 8.53383
R3537 VSS.n7310 VSS.n7309 8.53383
R3538 VSS.n7309 VSS.n7301 8.53383
R3539 VSS.n7304 VSS.n7301 8.53383
R3540 VSS.n7304 VSS.n7303 8.53383
R3541 VSS.n7286 VSS.n7285 8.53383
R3542 VSS.n7286 VSS.n7281 8.53383
R3543 VSS.n7349 VSS.n7281 8.53383
R3544 VSS.n7349 VSS.n7348 8.53383
R3545 VSS.n7348 VSS.n7291 8.53383
R3546 VSS.n7342 VSS.n7291 8.53383
R3547 VSS.n7342 VSS.n7341 8.53383
R3548 VSS.n10874 VSS.n3907 8.53383
R3549 VSS.n10864 VSS.n10861 8.53383
R3550 VSS.n10864 VSS.n10859 8.53383
R3551 VSS.n10867 VSS.n10859 8.53383
R3552 VSS.n10869 VSS.n10867 8.53383
R3553 VSS.n10872 VSS.n10869 8.53383
R3554 VSS.n10872 VSS.n3907 8.53383
R3555 VSS.n4135 VSS.n4132 8.53383
R3556 VSS.n4445 VSS.n4135 8.53383
R3557 VSS.n4445 VSS.n4137 8.53383
R3558 VSS.n4150 VSS.n4137 8.53383
R3559 VSS.n4150 VSS.n4139 8.53383
R3560 VSS.n4145 VSS.n4139 8.53383
R3561 VSS.n4145 VSS.n4144 8.53383
R3562 VSS.n4144 VSS.n4143 8.53383
R3563 VSS.n4390 VSS.n4387 8.53383
R3564 VSS.n4390 VSS.n4385 8.53383
R3565 VSS.n4395 VSS.n4385 8.53383
R3566 VSS.n4396 VSS.n4395 8.53383
R3567 VSS.n4399 VSS.n4396 8.53383
R3568 VSS.n4399 VSS.n4199 8.53383
R3569 VSS.n4401 VSS.n4199 8.53383
R3570 VSS.n4377 VSS.n4202 8.53383
R3571 VSS.n4375 VSS.n4202 8.53383
R3572 VSS.n4375 VSS.n4374 8.53383
R3573 VSS.n4374 VSS.n4372 8.53383
R3574 VSS.n4372 VSS.n4364 8.53383
R3575 VSS.n4369 VSS.n4364 8.53383
R3576 VSS.n4369 VSS.n4368 8.53383
R3577 VSS.n4368 VSS.n4365 8.53383
R3578 VSS.n4266 VSS.n4265 8.53383
R3579 VSS.n4265 VSS.n4256 8.53383
R3580 VSS.n4341 VSS.n4256 8.53383
R3581 VSS.n4341 VSS.n4340 8.53383
R3582 VSS.n4340 VSS.n4258 8.53383
R3583 VSS.n4337 VSS.n4258 8.53383
R3584 VSS.n4337 VSS.n4336 8.53383
R3585 VSS.n4336 VSS.n4333 8.53383
R3586 VSS.n4263 VSS.n4262 8.53383
R3587 VSS.n4322 VSS.n4263 8.53383
R3588 VSS.n4322 VSS.n4321 8.53383
R3589 VSS.n4321 VSS.n4307 8.53383
R3590 VSS.n4316 VSS.n4307 8.53383
R3591 VSS.n4316 VSS.n4315 8.53383
R3592 VSS.n4315 VSS.n4310 8.53383
R3593 VSS.n4313 VSS.n4310 8.53383
R3594 VSS.n4287 VSS.n4282 8.53383
R3595 VSS.n4287 VSS.n4280 8.53383
R3596 VSS.n4290 VSS.n4280 8.53383
R3597 VSS.n4290 VSS.n4278 8.53383
R3598 VSS.n4296 VSS.n4278 8.53383
R3599 VSS.n4296 VSS.n4273 8.53383
R3600 VSS.n4298 VSS.n4273 8.53383
R3601 VSS.n4347 VSS.n4230 8.53383
R3602 VSS.n4245 VSS.n4240 8.53383
R3603 VSS.n4246 VSS.n4245 8.53383
R3604 VSS.n4247 VSS.n4246 8.53383
R3605 VSS.n4247 VSS.n4231 8.53383
R3606 VSS.n4348 VSS.n4231 8.53383
R3607 VSS.n4348 VSS.n4347 8.53383
R3608 VSS.n4210 VSS.n4201 8.53383
R3609 VSS.n4212 VSS.n4210 8.53383
R3610 VSS.n4213 VSS.n4212 8.53383
R3611 VSS.n4223 VSS.n4213 8.53383
R3612 VSS.n4223 VSS.n4220 8.53383
R3613 VSS.n4220 VSS.n4217 8.53383
R3614 VSS.n4217 VSS.n4216 8.53383
R3615 VSS.n4216 VSS.n4214 8.53383
R3616 VSS.n4177 VSS.n4170 8.53383
R3617 VSS.n4177 VSS.n4176 8.53383
R3618 VSS.n4176 VSS.n4174 8.53383
R3619 VSS.n4174 VSS.n4163 8.53383
R3620 VSS.n4409 VSS.n4163 8.53383
R3621 VSS.n4409 VSS.n4408 8.53383
R3622 VSS.n4408 VSS.n4162 8.53383
R3623 VSS.n4417 VSS.n4131 8.53383
R3624 VSS.n4431 VSS.n4417 8.53383
R3625 VSS.n4431 VSS.n4430 8.53383
R3626 VSS.n4430 VSS.n4428 8.53383
R3627 VSS.n4428 VSS.n4427 8.53383
R3628 VSS.n4427 VSS.n4425 8.53383
R3629 VSS.n4425 VSS.n4422 8.53383
R3630 VSS.n4423 VSS.n4422 8.53383
R3631 VSS.n4124 VSS.n4123 8.53383
R3632 VSS.n4124 VSS.n4109 8.53383
R3633 VSS.n10780 VSS.n4109 8.53383
R3634 VSS.n10780 VSS.n10779 8.53383
R3635 VSS.n10779 VSS.n4111 8.53383
R3636 VSS.n4130 VSS.n4111 8.53383
R3637 VSS.n10773 VSS.n4130 8.53383
R3638 VSS.n10770 VSS.n4134 8.53383
R3639 VSS.n10758 VSS.n10753 8.53383
R3640 VSS.n10758 VSS.n10751 8.53383
R3641 VSS.n10761 VSS.n10751 8.53383
R3642 VSS.n10761 VSS.n10749 8.53383
R3643 VSS.n10768 VSS.n10749 8.53383
R3644 VSS.n10768 VSS.n4134 8.53383
R3645 VSS.n863 VSS.n862 8.53383
R3646 VSS.n1399 VSS.n863 8.53383
R3647 VSS.n1399 VSS.n864 8.53383
R3648 VSS.n870 VSS.n864 8.53383
R3649 VSS.n873 VSS.n870 8.53383
R3650 VSS.n875 VSS.n873 8.53383
R3651 VSS.n876 VSS.n875 8.53383
R3652 VSS.n876 VSS.n868 8.53383
R3653 VSS.n597 VSS.n593 8.53383
R3654 VSS.n598 VSS.n597 8.53383
R3655 VSS.n599 VSS.n598 8.53383
R3656 VSS.n599 VSS.n585 8.53383
R3657 VSS.n14205 VSS.n585 8.53383
R3658 VSS.n14205 VSS.n586 8.53383
R3659 VSS.n586 VSS.n584 8.53383
R3660 VSS.n14214 VSS.n14211 8.53383
R3661 VSS.n14214 VSS.n14209 8.53383
R3662 VSS.n14219 VSS.n14209 8.53383
R3663 VSS.n14220 VSS.n14219 8.53383
R3664 VSS.n14223 VSS.n14220 8.53383
R3665 VSS.n14223 VSS.n581 8.53383
R3666 VSS.n14225 VSS.n581 8.53383
R3667 VSS.n565 VSS.n560 8.53383
R3668 VSS.n566 VSS.n565 8.53383
R3669 VSS.n567 VSS.n566 8.53383
R3670 VSS.n567 VSS.n546 8.53383
R3671 VSS.n14233 VSS.n546 8.53383
R3672 VSS.n14233 VSS.n547 8.53383
R3673 VSS.n547 VSS.n545 8.53383
R3674 VSS.n1147 VSS.n934 8.53383
R3675 VSS.n1147 VSS.n1144 8.53383
R3676 VSS.n1144 VSS.n1143 8.53383
R3677 VSS.n1143 VSS.n1140 8.53383
R3678 VSS.n1140 VSS.n1139 8.53383
R3679 VSS.n1139 VSS.n936 8.53383
R3680 VSS.n1135 VSS.n936 8.53383
R3681 VSS.n911 VSS.n910 8.53383
R3682 VSS.n1155 VSS.n911 8.53383
R3683 VSS.n1155 VSS.n912 8.53383
R3684 VSS.n919 VSS.n912 8.53383
R3685 VSS.n925 VSS.n919 8.53383
R3686 VSS.n925 VSS.n924 8.53383
R3687 VSS.n924 VSS.n921 8.53383
R3688 VSS.n922 VSS.n921 8.53383
R3689 VSS.n14197 VSS.n605 8.53383
R3690 VSS.n14195 VSS.n605 8.53383
R3691 VSS.n14195 VSS.n14194 8.53383
R3692 VSS.n14194 VSS.n14179 8.53383
R3693 VSS.n14189 VSS.n14179 8.53383
R3694 VSS.n14189 VSS.n14188 8.53383
R3695 VSS.n14188 VSS.n14181 8.53383
R3696 VSS.n14184 VSS.n14181 8.53383
R3697 VSS.n12398 VSS.n2480 8.53383
R3698 VSS.n12418 VSS.n12398 8.53383
R3699 VSS.n12418 VSS.n12399 8.53383
R3700 VSS.n12410 VSS.n12399 8.53383
R3701 VSS.n12410 VSS.n12409 8.53383
R3702 VSS.n12409 VSS.n12408 8.53383
R3703 VSS.n12408 VSS.n12401 8.53383
R3704 VSS.n12403 VSS.n12401 8.53383
R3705 VSS.n13035 VSS.n13032 8.53383
R3706 VSS.n13036 VSS.n13035 8.53383
R3707 VSS.n13039 VSS.n13036 8.53383
R3708 VSS.n13039 VSS.n2497 8.53383
R3709 VSS.n13043 VSS.n2497 8.53383
R3710 VSS.n13043 VSS.n2498 8.53383
R3711 VSS.n2498 VSS.n2482 8.53383
R3712 VSS.n2533 VSS.n2481 8.53383
R3713 VSS.n2534 VSS.n2533 8.53383
R3714 VSS.n2537 VSS.n2534 8.53383
R3715 VSS.n2546 VSS.n2537 8.53383
R3716 VSS.n2546 VSS.n2543 8.53383
R3717 VSS.n2543 VSS.n2542 8.53383
R3718 VSS.n2542 VSS.n2541 8.53383
R3719 VSS.n2541 VSS.n2539 8.53383
R3720 VSS.n2473 VSS.n2468 8.53383
R3721 VSS.n2474 VSS.n2473 8.53383
R3722 VSS.n2475 VSS.n2474 8.53383
R3723 VSS.n2475 VSS.n2462 8.53383
R3724 VSS.n13057 VSS.n2462 8.53383
R3725 VSS.n13057 VSS.n2463 8.53383
R3726 VSS.n2463 VSS.n2461 8.53383
R3727 VSS.n2437 VSS.n2436 8.53383
R3728 VSS.n2437 VSS.n2431 8.53383
R3729 VSS.n2444 VSS.n2431 8.53383
R3730 VSS.n2444 VSS.n2394 8.53383
R3731 VSS.n2448 VSS.n2394 8.53383
R3732 VSS.n2449 VSS.n2448 8.53383
R3733 VSS.n2449 VSS.n2392 8.53383
R3734 VSS.n2368 VSS.n2367 8.53383
R3735 VSS.n2368 VSS.n2352 8.53383
R3736 VSS.n13104 VSS.n2352 8.53383
R3737 VSS.n13104 VSS.n2353 8.53383
R3738 VSS.n13099 VSS.n2353 8.53383
R3739 VSS.n13099 VSS.n13098 8.53383
R3740 VSS.n13098 VSS.n13097 8.53383
R3741 VSS.n2391 VSS.n2374 8.53383
R3742 VSS.n2389 VSS.n2374 8.53383
R3743 VSS.n2389 VSS.n2388 8.53383
R3744 VSS.n2388 VSS.n2386 8.53383
R3745 VSS.n2386 VSS.n2376 8.53383
R3746 VSS.n2381 VSS.n2376 8.53383
R3747 VSS.n2381 VSS.n2380 8.53383
R3748 VSS.n2380 VSS.n2377 8.53383
R3749 VSS.n13091 VSS.n2455 8.53383
R3750 VSS.n13089 VSS.n2455 8.53383
R3751 VSS.n13089 VSS.n13088 8.53383
R3752 VSS.n13088 VSS.n13073 8.53383
R3753 VSS.n13083 VSS.n13073 8.53383
R3754 VSS.n13083 VSS.n13082 8.53383
R3755 VSS.n13082 VSS.n13075 8.53383
R3756 VSS.n13078 VSS.n13075 8.53383
R3757 VSS.n1912 VSS.n1911 8.53383
R3758 VSS.n13137 VSS.n1912 8.53383
R3759 VSS.n13137 VSS.n1913 8.53383
R3760 VSS.n1919 VSS.n1913 8.53383
R3761 VSS.n1922 VSS.n1919 8.53383
R3762 VSS.n1924 VSS.n1922 8.53383
R3763 VSS.n1925 VSS.n1924 8.53383
R3764 VSS.n1925 VSS.n1917 8.53383
R3765 VSS.n2338 VSS.n1944 8.53383
R3766 VSS.n2338 VSS.n2335 8.53383
R3767 VSS.n2335 VSS.n2334 8.53383
R3768 VSS.n2334 VSS.n2331 8.53383
R3769 VSS.n2331 VSS.n2330 8.53383
R3770 VSS.n2330 VSS.n1946 8.53383
R3771 VSS.n1946 VSS.n1930 8.53383
R3772 VSS.n2281 VSS.n1929 8.53383
R3773 VSS.n2295 VSS.n2281 8.53383
R3774 VSS.n2295 VSS.n2292 8.53383
R3775 VSS.n2292 VSS.n2291 8.53383
R3776 VSS.n2291 VSS.n2288 8.53383
R3777 VSS.n2288 VSS.n2287 8.53383
R3778 VSS.n2287 VSS.n2282 8.53383
R3779 VSS.n2283 VSS.n2282 8.53383
R3780 VSS.n13117 VSS.n13112 8.53383
R3781 VSS.n13117 VSS.n13110 8.53383
R3782 VSS.n13120 VSS.n13110 8.53383
R3783 VSS.n13120 VSS.n13108 8.53383
R3784 VSS.n13126 VSS.n13108 8.53383
R3785 VSS.n13126 VSS.n2349 8.53383
R3786 VSS.n13128 VSS.n2349 8.53383
R3787 VSS.n14158 VSS.n14157 8.53383
R3788 VSS.n14160 VSS.n14158 8.53383
R3789 VSS.n14161 VSS.n14160 8.53383
R3790 VSS.n14171 VSS.n14161 8.53383
R3791 VSS.n14171 VSS.n14168 8.53383
R3792 VSS.n14168 VSS.n14165 8.53383
R3793 VSS.n14165 VSS.n14164 8.53383
R3794 VSS.n14164 VSS.n14162 8.53383
R3795 VSS.n2404 VSS.n2403 8.53383
R3796 VSS.n2418 VSS.n2404 8.53383
R3797 VSS.n2418 VSS.n2417 8.53383
R3798 VSS.n2417 VSS.n2415 8.53383
R3799 VSS.n2415 VSS.n2414 8.53383
R3800 VSS.n2414 VSS.n2412 8.53383
R3801 VSS.n2412 VSS.n2407 8.53383
R3802 VSS.n2408 VSS.n2407 8.53383
R3803 VSS.n896 VSS.n881 8.53383
R3804 VSS.n1162 VSS.n896 8.53383
R3805 VSS.n1162 VSS.n897 8.53383
R3806 VSS.n907 VSS.n897 8.53383
R3807 VSS.n907 VSS.n906 8.53383
R3808 VSS.n906 VSS.n904 8.53383
R3809 VSS.n904 VSS.n903 8.53383
R3810 VSS.n903 VSS.n901 8.53383
R3811 VSS.n942 VSS.n939 8.53383
R3812 VSS.n945 VSS.n942 8.53383
R3813 VSS.n946 VSS.n945 8.53383
R3814 VSS.n949 VSS.n946 8.53383
R3815 VSS.n953 VSS.n949 8.53383
R3816 VSS.n953 VSS.n950 8.53383
R3817 VSS.n950 VSS.n882 8.53383
R3818 VSS.n1381 VSS.n1374 8.53383
R3819 VSS.n1382 VSS.n1381 8.53383
R3820 VSS.n1382 VSS.n1372 8.53383
R3821 VSS.n1372 VSS.n1370 8.53383
R3822 VSS.n1389 VSS.n1370 8.53383
R3823 VSS.n1389 VSS.n1170 8.53383
R3824 VSS.n1391 VSS.n1170 8.53383
R3825 VSS.n1687 VSS.n1461 8.53383
R3826 VSS.n1687 VSS.n1684 8.53383
R3827 VSS.n1684 VSS.n1674 8.53383
R3828 VSS.n1694 VSS.n1674 8.53383
R3829 VSS.n1694 VSS.n1675 8.53383
R3830 VSS.n1680 VSS.n1675 8.53383
R3831 VSS.n1680 VSS.n1679 8.53383
R3832 VSS.n1679 VSS.n1678 8.53383
R3833 VSS.n629 VSS.n628 8.53383
R3834 VSS.n14119 VSS.n629 8.53383
R3835 VSS.n14119 VSS.n14118 8.53383
R3836 VSS.n14118 VSS.n631 8.53383
R3837 VSS.n646 VSS.n631 8.53383
R3838 VSS.n646 VSS.n645 8.53383
R3839 VSS.n645 VSS.n642 8.53383
R3840 VSS.n643 VSS.n642 8.53383
R3841 VSS.n1448 VSS.n1445 8.53383
R3842 VSS.n1448 VSS.n1442 8.53383
R3843 VSS.n1451 VSS.n1442 8.53383
R3844 VSS.n1454 VSS.n1451 8.53383
R3845 VSS.n1457 VSS.n1454 8.53383
R3846 VSS.n1457 VSS.n652 8.53383
R3847 VSS.n1460 VSS.n652 8.53383
R3848 VSS.n14098 VSS.n14091 8.53383
R3849 VSS.n14099 VSS.n14098 8.53383
R3850 VSS.n14099 VSS.n14089 8.53383
R3851 VSS.n14089 VSS.n14087 8.53383
R3852 VSS.n14106 VSS.n14087 8.53383
R3853 VSS.n14106 VSS.n1463 8.53383
R3854 VSS.n14108 VSS.n1463 8.53383
R3855 VSS.n13694 VSS.n13671 8.53383
R3856 VSS.n13673 VSS.n13671 8.53383
R3857 VSS.n13688 VSS.n13673 8.53383
R3858 VSS.n13688 VSS.n13687 8.53383
R3859 VSS.n13687 VSS.n13675 8.53383
R3860 VSS.n13684 VSS.n13675 8.53383
R3861 VSS.n13684 VSS.n13677 8.53383
R3862 VSS.n13677 VSS.n13676 8.53383
R3863 VSS.n14077 VSS.n1671 8.53383
R3864 VSS.n14075 VSS.n1671 8.53383
R3865 VSS.n14075 VSS.n14074 8.53383
R3866 VSS.n14074 VSS.n14072 8.53383
R3867 VSS.n14072 VSS.n14064 8.53383
R3868 VSS.n14069 VSS.n14064 8.53383
R3869 VSS.n14069 VSS.n14068 8.53383
R3870 VSS.n14068 VSS.n14065 8.53383
R3871 VSS.n1654 VSS.n1653 8.53383
R3872 VSS.n1653 VSS.n1642 8.53383
R3873 VSS.n14083 VSS.n1642 8.53383
R3874 VSS.n14083 VSS.n14082 8.53383
R3875 VSS.n14082 VSS.n1644 8.53383
R3876 VSS.n1665 VSS.n1644 8.53383
R3877 VSS.n1666 VSS.n1665 8.53383
R3878 VSS.n13700 VSS.n13652 8.53383
R3879 VSS.n13662 VSS.n13655 8.53383
R3880 VSS.n13663 VSS.n13662 8.53383
R3881 VSS.n13664 VSS.n13663 8.53383
R3882 VSS.n13664 VSS.n13653 8.53383
R3883 VSS.n13701 VSS.n13653 8.53383
R3884 VSS.n13701 VSS.n13700 8.53383
R3885 VSS.n13205 VSS.n13204 8.53383
R3886 VSS.n13907 VSS.n13205 8.53383
R3887 VSS.n13907 VSS.n13206 8.53383
R3888 VSS.n13212 VSS.n13206 8.53383
R3889 VSS.n13215 VSS.n13212 8.53383
R3890 VSS.n13217 VSS.n13215 8.53383
R3891 VSS.n13218 VSS.n13217 8.53383
R3892 VSS.n13218 VSS.n13210 8.53383
R3893 VSS.n13633 VSS.n13630 8.53383
R3894 VSS.n13634 VSS.n13633 8.53383
R3895 VSS.n13637 VSS.n13634 8.53383
R3896 VSS.n13637 VSS.n13238 8.53383
R3897 VSS.n13641 VSS.n13238 8.53383
R3898 VSS.n13641 VSS.n13239 8.53383
R3899 VSS.n13239 VSS.n13223 8.53383
R3900 VSS.n13532 VSS.n13222 8.53383
R3901 VSS.n13533 VSS.n13532 8.53383
R3902 VSS.n13536 VSS.n13533 8.53383
R3903 VSS.n13545 VSS.n13536 8.53383
R3904 VSS.n13545 VSS.n13542 8.53383
R3905 VSS.n13542 VSS.n13541 8.53383
R3906 VSS.n13541 VSS.n13540 8.53383
R3907 VSS.n13540 VSS.n13538 8.53383
R3908 VSS.n13887 VSS.n13882 8.53383
R3909 VSS.n13887 VSS.n13880 8.53383
R3910 VSS.n13890 VSS.n13880 8.53383
R3911 VSS.n13890 VSS.n13878 8.53383
R3912 VSS.n13896 VSS.n13878 8.53383
R3913 VSS.n13896 VSS.n13650 8.53383
R3914 VSS.n13898 VSS.n13650 8.53383
R3915 VSS.n815 VSS.n813 8.53383
R3916 VSS.n830 VSS.n825 8.53383
R3917 VSS.n831 VSS.n830 8.53383
R3918 VSS.n832 VSS.n831 8.53383
R3919 VSS.n832 VSS.n814 8.53383
R3920 VSS.n1438 VSS.n814 8.53383
R3921 VSS.n1438 VSS.n815 8.53383
R3922 VSS.n844 VSS.n840 8.53383
R3923 VSS.n1406 VSS.n844 8.53383
R3924 VSS.n1406 VSS.n846 8.53383
R3925 VSS.n859 VSS.n846 8.53383
R3926 VSS.n859 VSS.n858 8.53383
R3927 VSS.n858 VSS.n850 8.53383
R3928 VSS.n851 VSS.n850 8.53383
R3929 VSS.n852 VSS.n851 8.53383
R3930 VSS.n1180 VSS.n1176 8.53383
R3931 VSS.n1185 VSS.n1176 8.53383
R3932 VSS.n1186 VSS.n1185 8.53383
R3933 VSS.n1186 VSS.n1173 8.53383
R3934 VSS.n1194 VSS.n1173 8.53383
R3935 VSS.n1194 VSS.n1174 8.53383
R3936 VSS.n1174 VSS.n841 8.53383
R3937 VSS.n1432 VSS.n1416 8.53383
R3938 VSS.n1432 VSS.n1431 8.53383
R3939 VSS.n1431 VSS.n1429 8.53383
R3940 VSS.n1429 VSS.n1427 8.53383
R3941 VSS.n1427 VSS.n1417 8.53383
R3942 VSS.n1422 VSS.n1417 8.53383
R3943 VSS.n1422 VSS.n1419 8.53383
R3944 VSS.n1419 VSS.n1418 8.53383
R3945 VSS.n2208 VSS.n2054 8.53383
R3946 VSS.n2208 VSS.n2207 8.53383
R3947 VSS.n2207 VSS.n2056 8.53383
R3948 VSS.n2203 VSS.n2056 8.53383
R3949 VSS.n2203 VSS.n2190 8.53383
R3950 VSS.n2193 VSS.n2190 8.53383
R3951 VSS.n2196 VSS.n2193 8.53383
R3952 VSS.n2196 VSS.n2195 8.53383
R3953 VSS.n1984 VSS.n1983 8.53383
R3954 VSS.n2249 VSS.n1984 8.53383
R3955 VSS.n2249 VSS.n2248 8.53383
R3956 VSS.n2248 VSS.n1986 8.53383
R3957 VSS.n2001 VSS.n1986 8.53383
R3958 VSS.n2001 VSS.n2000 8.53383
R3959 VSS.n2000 VSS.n1997 8.53383
R3960 VSS.n1998 VSS.n1997 8.53383
R3961 VSS.n2042 VSS.n2039 8.53383
R3962 VSS.n2042 VSS.n2036 8.53383
R3963 VSS.n2045 VSS.n2036 8.53383
R3964 VSS.n2048 VSS.n2045 8.53383
R3965 VSS.n2051 VSS.n2048 8.53383
R3966 VSS.n2051 VSS.n2007 8.53383
R3967 VSS.n2053 VSS.n2007 8.53383
R3968 VSS.n2238 VSS.n2213 8.53383
R3969 VSS.n2226 VSS.n2221 8.53383
R3970 VSS.n2226 VSS.n2219 8.53383
R3971 VSS.n2229 VSS.n2219 8.53383
R3972 VSS.n2229 VSS.n2217 8.53383
R3973 VSS.n2236 VSS.n2217 8.53383
R3974 VSS.n2236 VSS.n2213 8.53383
R3975 VSS.n2124 VSS.n2103 8.53383
R3976 VSS.n2124 VSS.n2123 8.53383
R3977 VSS.n2123 VSS.n2121 8.53383
R3978 VSS.n2121 VSS.n2105 8.53383
R3979 VSS.n2116 VSS.n2105 8.53383
R3980 VSS.n2116 VSS.n2115 8.53383
R3981 VSS.n2115 VSS.n2108 8.53383
R3982 VSS.n2113 VSS.n2108 8.53383
R3983 VSS.n2059 VSS.n2058 8.53383
R3984 VSS.n2184 VSS.n2059 8.53383
R3985 VSS.n2184 VSS.n2183 8.53383
R3986 VSS.n2183 VSS.n2061 8.53383
R3987 VSS.n2076 VSS.n2061 8.53383
R3988 VSS.n2076 VSS.n2075 8.53383
R3989 VSS.n2075 VSS.n2072 8.53383
R3990 VSS.n2073 VSS.n2072 8.53383
R3991 VSS.n2091 VSS.n2088 8.53383
R3992 VSS.n2091 VSS.n2085 8.53383
R3993 VSS.n2094 VSS.n2085 8.53383
R3994 VSS.n2097 VSS.n2094 8.53383
R3995 VSS.n2100 VSS.n2097 8.53383
R3996 VSS.n2100 VSS.n2082 8.53383
R3997 VSS.n2102 VSS.n2082 8.53383
R3998 VSS.n2173 VSS.n2129 8.53383
R3999 VSS.n2161 VSS.n2156 8.53383
R4000 VSS.n2161 VSS.n2154 8.53383
R4001 VSS.n2164 VSS.n2154 8.53383
R4002 VSS.n2164 VSS.n2152 8.53383
R4003 VSS.n2171 VSS.n2152 8.53383
R4004 VSS.n2171 VSS.n2129 8.53383
R4005 VSS.n12651 VSS.n1851 8.53383
R4006 VSS.n12652 VSS.n12651 8.53383
R4007 VSS.n12652 VSS.n12647 8.53383
R4008 VSS.n12666 VSS.n12647 8.53383
R4009 VSS.n12666 VSS.n12648 8.53383
R4010 VSS.n12656 VSS.n12648 8.53383
R4011 VSS.n12659 VSS.n12656 8.53383
R4012 VSS.n12659 VSS.n12658 8.53383
R4013 VSS.n1867 VSS.n1852 8.53383
R4014 VSS.n13185 VSS.n1867 8.53383
R4015 VSS.n13185 VSS.n1868 8.53383
R4016 VSS.n1878 VSS.n1868 8.53383
R4017 VSS.n1878 VSS.n1877 8.53383
R4018 VSS.n1877 VSS.n1875 8.53383
R4019 VSS.n1875 VSS.n1874 8.53383
R4020 VSS.n1874 VSS.n1872 8.53383
R4021 VSS.n2137 VSS.n2136 8.53383
R4022 VSS.n2140 VSS.n2137 8.53383
R4023 VSS.n2148 VSS.n2140 8.53383
R4024 VSS.n2148 VSS.n2147 8.53383
R4025 VSS.n2147 VSS.n2145 8.53383
R4026 VSS.n2145 VSS.n2144 8.53383
R4027 VSS.n2144 VSS.n1853 8.53383
R4028 VSS.n13198 VSS.n1831 8.53383
R4029 VSS.n1843 VSS.n1838 8.53383
R4030 VSS.n1844 VSS.n1843 8.53383
R4031 VSS.n1845 VSS.n1844 8.53383
R4032 VSS.n1845 VSS.n1832 8.53383
R4033 VSS.n13199 VSS.n1832 8.53383
R4034 VSS.n13199 VSS.n13198 8.53383
R4035 VSS.n12670 VSS.n1813 8.53383
R4036 VSS.n12691 VSS.n12670 8.53383
R4037 VSS.n12691 VSS.n12671 8.53383
R4038 VSS.n12682 VSS.n12671 8.53383
R4039 VSS.n12682 VSS.n12681 8.53383
R4040 VSS.n12681 VSS.n12680 8.53383
R4041 VSS.n12680 VSS.n12673 8.53383
R4042 VSS.n12675 VSS.n12673 8.53383
R4043 VSS.n1789 VSS.n1788 8.53383
R4044 VSS.n1789 VSS.n1773 8.53383
R4045 VSS.n13938 VSS.n1773 8.53383
R4046 VSS.n13938 VSS.n1774 8.53383
R4047 VSS.n13933 VSS.n1774 8.53383
R4048 VSS.n13933 VSS.n13932 8.53383
R4049 VSS.n13932 VSS.n13931 8.53383
R4050 VSS.n1812 VSS.n1795 8.53383
R4051 VSS.n1810 VSS.n1795 8.53383
R4052 VSS.n1810 VSS.n1809 8.53383
R4053 VSS.n1809 VSS.n1807 8.53383
R4054 VSS.n1807 VSS.n1797 8.53383
R4055 VSS.n1802 VSS.n1797 8.53383
R4056 VSS.n1802 VSS.n1801 8.53383
R4057 VSS.n1801 VSS.n1798 8.53383
R4058 VSS.n1828 VSS.n1822 8.53383
R4059 VSS.n1828 VSS.n1818 8.53383
R4060 VSS.n13917 VSS.n1818 8.53383
R4061 VSS.n13918 VSS.n13917 8.53383
R4062 VSS.n13919 VSS.n13918 8.53383
R4063 VSS.n13919 VSS.n1815 8.53383
R4064 VSS.n13925 VSS.n1815 8.53383
R4065 VSS.n2012 VSS.n1977 8.53383
R4066 VSS.n2021 VSS.n2014 8.53383
R4067 VSS.n2022 VSS.n2021 8.53383
R4068 VSS.n2023 VSS.n2022 8.53383
R4069 VSS.n2023 VSS.n2011 8.53383
R4070 VSS.n2032 VSS.n2011 8.53383
R4071 VSS.n2032 VSS.n2012 8.53383
R4072 VSS.n2317 VSS.n2279 8.53383
R4073 VSS.n2315 VSS.n2279 8.53383
R4074 VSS.n2315 VSS.n2312 8.53383
R4075 VSS.n2312 VSS.n2311 8.53383
R4076 VSS.n2311 VSS.n2301 8.53383
R4077 VSS.n2306 VSS.n2301 8.53383
R4078 VSS.n2306 VSS.n2303 8.53383
R4079 VSS.n2303 VSS.n2302 8.53383
R4080 VSS.n1962 VSS.n1957 8.53383
R4081 VSS.n1963 VSS.n1962 8.53383
R4082 VSS.n1964 VSS.n1963 8.53383
R4083 VSS.n1964 VSS.n1949 8.53383
R4084 VSS.n2322 VSS.n1949 8.53383
R4085 VSS.n2322 VSS.n1950 8.53383
R4086 VSS.n1950 VSS.n1948 8.53383
R4087 VSS.n2276 VSS.n1981 8.53383
R4088 VSS.n2274 VSS.n1981 8.53383
R4089 VSS.n2274 VSS.n2255 8.53383
R4090 VSS.n2267 VSS.n2255 8.53383
R4091 VSS.n2267 VSS.n2257 8.53383
R4092 VSS.n2264 VSS.n2257 8.53383
R4093 VSS.n2264 VSS.n2259 8.53383
R4094 VSS.n2259 VSS.n2258 8.53383
R4095 VSS.n2700 VSS.n2661 8.53383
R4096 VSS.n2721 VSS.n2700 8.53383
R4097 VSS.n2721 VSS.n2701 8.53383
R4098 VSS.n2712 VSS.n2701 8.53383
R4099 VSS.n2712 VSS.n2711 8.53383
R4100 VSS.n2711 VSS.n2710 8.53383
R4101 VSS.n2710 VSS.n2703 8.53383
R4102 VSS.n2705 VSS.n2703 8.53383
R4103 VSS.n2563 VSS.n2562 8.53383
R4104 VSS.n12989 VSS.n2563 8.53383
R4105 VSS.n12989 VSS.n12988 8.53383
R4106 VSS.n12988 VSS.n2565 8.53383
R4107 VSS.n2580 VSS.n2565 8.53383
R4108 VSS.n2580 VSS.n2579 8.53383
R4109 VSS.n2579 VSS.n2576 8.53383
R4110 VSS.n2577 VSS.n2576 8.53383
R4111 VSS.n2649 VSS.n2646 8.53383
R4112 VSS.n2649 VSS.n2643 8.53383
R4113 VSS.n2652 VSS.n2643 8.53383
R4114 VSS.n2655 VSS.n2652 8.53383
R4115 VSS.n2658 VSS.n2655 8.53383
R4116 VSS.n2658 VSS.n2586 8.53383
R4117 VSS.n2660 VSS.n2586 8.53383
R4118 VSS.n12966 VSS.n12961 8.53383
R4119 VSS.n12966 VSS.n12959 8.53383
R4120 VSS.n12969 VSS.n12959 8.53383
R4121 VSS.n12969 VSS.n12957 8.53383
R4122 VSS.n12976 VSS.n12957 8.53383
R4123 VSS.n12976 VSS.n2663 8.53383
R4124 VSS.n12978 VSS.n2663 8.53383
R4125 VSS.n12947 VSS.n2698 8.53383
R4126 VSS.n12945 VSS.n2698 8.53383
R4127 VSS.n12945 VSS.n12944 8.53383
R4128 VSS.n12944 VSS.n12942 8.53383
R4129 VSS.n12942 VSS.n12934 8.53383
R4130 VSS.n12939 VSS.n12934 8.53383
R4131 VSS.n12939 VSS.n12938 8.53383
R4132 VSS.n12938 VSS.n12935 8.53383
R4133 VSS.n2681 VSS.n2680 8.53383
R4134 VSS.n2680 VSS.n2669 8.53383
R4135 VSS.n12953 VSS.n2669 8.53383
R4136 VSS.n12953 VSS.n12952 8.53383
R4137 VSS.n12952 VSS.n2671 8.53383
R4138 VSS.n2692 VSS.n2671 8.53383
R4139 VSS.n2693 VSS.n2692 8.53383
R4140 VSS.n2780 VSS.n2773 8.53383
R4141 VSS.n2781 VSS.n2780 8.53383
R4142 VSS.n2782 VSS.n2781 8.53383
R4143 VSS.n2782 VSS.n2771 8.53383
R4144 VSS.n2819 VSS.n2771 8.53383
R4145 VSS.n2819 VSS.n2818 8.53383
R4146 VSS.n2818 VSS.n2770 8.53383
R4147 VSS.n2744 VSS.n2743 8.53383
R4148 VSS.n12912 VSS.n2744 8.53383
R4149 VSS.n12912 VSS.n12911 8.53383
R4150 VSS.n12911 VSS.n2746 8.53383
R4151 VSS.n2761 VSS.n2746 8.53383
R4152 VSS.n2761 VSS.n2760 8.53383
R4153 VSS.n2760 VSS.n2757 8.53383
R4154 VSS.n2758 VSS.n2757 8.53383
R4155 VSS.n2830 VSS.n2827 8.53383
R4156 VSS.n2830 VSS.n2824 8.53383
R4157 VSS.n2833 VSS.n2824 8.53383
R4158 VSS.n2836 VSS.n2833 8.53383
R4159 VSS.n2839 VSS.n2836 8.53383
R4160 VSS.n2839 VSS.n2767 8.53383
R4161 VSS.n2841 VSS.n2767 8.53383
R4162 VSS.n12889 VSS.n12884 8.53383
R4163 VSS.n12889 VSS.n12882 8.53383
R4164 VSS.n12892 VSS.n12882 8.53383
R4165 VSS.n12892 VSS.n12880 8.53383
R4166 VSS.n12899 VSS.n12880 8.53383
R4167 VSS.n12899 VSS.n2844 8.53383
R4168 VSS.n12901 VSS.n2844 8.53383
R4169 VSS.n12635 VSS.n3055 8.53383
R4170 VSS.n3057 VSS.n3055 8.53383
R4171 VSS.n12629 VSS.n3057 8.53383
R4172 VSS.n12629 VSS.n12628 8.53383
R4173 VSS.n12628 VSS.n3059 8.53383
R4174 VSS.n12625 VSS.n3059 8.53383
R4175 VSS.n12625 VSS.n12618 8.53383
R4176 VSS.n12618 VSS.n12617 8.53383
R4177 VSS.n12870 VSS.n2878 8.53383
R4178 VSS.n12868 VSS.n2878 8.53383
R4179 VSS.n12868 VSS.n12867 8.53383
R4180 VSS.n12867 VSS.n12865 8.53383
R4181 VSS.n12865 VSS.n12857 8.53383
R4182 VSS.n12862 VSS.n12857 8.53383
R4183 VSS.n12862 VSS.n12861 8.53383
R4184 VSS.n12861 VSS.n12858 8.53383
R4185 VSS.n2861 VSS.n2860 8.53383
R4186 VSS.n2860 VSS.n2849 8.53383
R4187 VSS.n12876 VSS.n2849 8.53383
R4188 VSS.n12876 VSS.n12875 8.53383
R4189 VSS.n12875 VSS.n2851 8.53383
R4190 VSS.n2872 VSS.n2851 8.53383
R4191 VSS.n2873 VSS.n2872 8.53383
R4192 VSS.n12641 VSS.n3036 8.53383
R4193 VSS.n3046 VSS.n3039 8.53383
R4194 VSS.n3047 VSS.n3046 8.53383
R4195 VSS.n3048 VSS.n3047 8.53383
R4196 VSS.n3048 VSS.n3037 8.53383
R4197 VSS.n12642 VSS.n3037 8.53383
R4198 VSS.n12642 VSS.n12641 8.53383
R4199 VSS.n3061 VSS.n3018 8.53383
R4200 VSS.n3082 VSS.n3061 8.53383
R4201 VSS.n3082 VSS.n3062 8.53383
R4202 VSS.n3073 VSS.n3062 8.53383
R4203 VSS.n3073 VSS.n3072 8.53383
R4204 VSS.n3072 VSS.n3071 8.53383
R4205 VSS.n3071 VSS.n3064 8.53383
R4206 VSS.n3066 VSS.n3064 8.53383
R4207 VSS.n2967 VSS.n2966 8.53383
R4208 VSS.n2967 VSS.n2951 8.53383
R4209 VSS.n12733 VSS.n2951 8.53383
R4210 VSS.n12733 VSS.n2952 8.53383
R4211 VSS.n12728 VSS.n2952 8.53383
R4212 VSS.n12728 VSS.n12727 8.53383
R4213 VSS.n12727 VSS.n12726 8.53383
R4214 VSS.n3017 VSS.n2973 8.53383
R4215 VSS.n3015 VSS.n2973 8.53383
R4216 VSS.n3015 VSS.n3014 8.53383
R4217 VSS.n3014 VSS.n3012 8.53383
R4218 VSS.n3012 VSS.n3002 8.53383
R4219 VSS.n3007 VSS.n3002 8.53383
R4220 VSS.n3007 VSS.n3006 8.53383
R4221 VSS.n3006 VSS.n3003 8.53383
R4222 VSS.n3033 VSS.n3027 8.53383
R4223 VSS.n3033 VSS.n3023 8.53383
R4224 VSS.n12712 VSS.n3023 8.53383
R4225 VSS.n12713 VSS.n12712 8.53383
R4226 VSS.n12714 VSS.n12713 8.53383
R4227 VSS.n12714 VSS.n3020 8.53383
R4228 VSS.n12720 VSS.n3020 8.53383
R4229 VSS.n2592 VSS.n2590 8.53383
R4230 VSS.n2601 VSS.n2594 8.53383
R4231 VSS.n2602 VSS.n2601 8.53383
R4232 VSS.n2603 VSS.n2602 8.53383
R4233 VSS.n2603 VSS.n2591 8.53383
R4234 VSS.n2639 VSS.n2591 8.53383
R4235 VSS.n2639 VSS.n2592 8.53383
R4236 VSS.n13022 VSS.n2530 8.53383
R4237 VSS.n13020 VSS.n2530 8.53383
R4238 VSS.n13020 VSS.n13017 8.53383
R4239 VSS.n13017 VSS.n13016 8.53383
R4240 VSS.n13016 VSS.n13006 8.53383
R4241 VSS.n13011 VSS.n13006 8.53383
R4242 VSS.n13011 VSS.n13008 8.53383
R4243 VSS.n13008 VSS.n13007 8.53383
R4244 VSS.n2514 VSS.n2509 8.53383
R4245 VSS.n2515 VSS.n2514 8.53383
R4246 VSS.n2516 VSS.n2515 8.53383
R4247 VSS.n2516 VSS.n2501 8.53383
R4248 VSS.n13027 VSS.n2501 8.53383
R4249 VSS.n13027 VSS.n2502 8.53383
R4250 VSS.n2502 VSS.n2500 8.53383
R4251 VSS.n2631 VSS.n2609 8.53383
R4252 VSS.n2629 VSS.n2609 8.53383
R4253 VSS.n2629 VSS.n2610 8.53383
R4254 VSS.n2622 VSS.n2610 8.53383
R4255 VSS.n2622 VSS.n2612 8.53383
R4256 VSS.n2619 VSS.n2612 8.53383
R4257 VSS.n2619 VSS.n2614 8.53383
R4258 VSS.n2614 VSS.n2613 8.53383
R4259 VSS.n2976 VSS.n2943 8.53383
R4260 VSS.n2996 VSS.n2976 8.53383
R4261 VSS.n2996 VSS.n2995 8.53383
R4262 VSS.n2995 VSS.n2981 8.53383
R4263 VSS.n2990 VSS.n2981 8.53383
R4264 VSS.n2990 VSS.n2989 8.53383
R4265 VSS.n2989 VSS.n2984 8.53383
R4266 VSS.n2987 VSS.n2984 8.53383
R4267 VSS.n12742 VSS.n12741 8.53383
R4268 VSS.n12742 VSS.n12737 8.53383
R4269 VSS.n12748 VSS.n12737 8.53383
R4270 VSS.n12748 VSS.n2948 8.53383
R4271 VSS.n12752 VSS.n2948 8.53383
R4272 VSS.n12752 VSS.n2946 8.53383
R4273 VSS.n2946 VSS.n2944 8.53383
R4274 VSS.n12779 VSS.n12761 8.53383
R4275 VSS.n12769 VSS.n12766 8.53383
R4276 VSS.n12769 VSS.n12764 8.53383
R4277 VSS.n12772 VSS.n12764 8.53383
R4278 VSS.n12774 VSS.n12772 8.53383
R4279 VSS.n12777 VSS.n12774 8.53383
R4280 VSS.n12777 VSS.n12761 8.53383
R4281 VSS.n1760 VSS.n1759 8.53383
R4282 VSS.n13987 VSS.n1760 8.53383
R4283 VSS.n13987 VSS.n13986 8.53383
R4284 VSS.n13986 VSS.n13972 8.53383
R4285 VSS.n13981 VSS.n13972 8.53383
R4286 VSS.n13981 VSS.n13980 8.53383
R4287 VSS.n13980 VSS.n13975 8.53383
R4288 VSS.n13978 VSS.n13975 8.53383
R4289 VSS.n13952 VSS.n13947 8.53383
R4290 VSS.n13952 VSS.n13945 8.53383
R4291 VSS.n13955 VSS.n13945 8.53383
R4292 VSS.n13955 VSS.n13943 8.53383
R4293 VSS.n13961 VSS.n13943 8.53383
R4294 VSS.n13961 VSS.n1770 8.53383
R4295 VSS.n13963 VSS.n1770 8.53383
R4296 VSS.n14019 VSS.n1716 8.53383
R4297 VSS.n1731 VSS.n1726 8.53383
R4298 VSS.n1732 VSS.n1731 8.53383
R4299 VSS.n1733 VSS.n1732 8.53383
R4300 VSS.n1733 VSS.n1717 8.53383
R4301 VSS.n14020 VSS.n1717 8.53383
R4302 VSS.n14020 VSS.n14019 8.53383
R4303 VSS.n13553 VSS.n13510 8.53383
R4304 VSS.n13553 VSS.n13552 8.53383
R4305 VSS.n13552 VSS.n13514 8.53383
R4306 VSS.n13528 VSS.n13514 8.53383
R4307 VSS.n13528 VSS.n13527 8.53383
R4308 VSS.n13527 VSS.n13519 8.53383
R4309 VSS.n13522 VSS.n13519 8.53383
R4310 VSS.n13522 VSS.n13521 8.53383
R4311 VSS.n13569 VSS.n13563 8.53383
R4312 VSS.n13569 VSS.n13559 8.53383
R4313 VSS.n13572 VSS.n13559 8.53383
R4314 VSS.n13573 VSS.n13572 8.53383
R4315 VSS.n13575 VSS.n13573 8.53383
R4316 VSS.n13575 VSS.n13557 8.53383
R4317 VSS.n13557 VSS.n13511 8.53383
R4318 VSS.n13606 VSS.n13481 8.53383
R4319 VSS.n13496 VSS.n13491 8.53383
R4320 VSS.n13497 VSS.n13496 8.53383
R4321 VSS.n13498 VSS.n13497 8.53383
R4322 VSS.n13498 VSS.n13482 8.53383
R4323 VSS.n13607 VSS.n13482 8.53383
R4324 VSS.n13607 VSS.n13606 8.53383
R4325 VSS.n11420 VSS.n11414 8.28285
R4326 VSS.n8494 VSS.n8493 8.0005
R4327 VSS.n8373 VSS.n8372 8.0005
R4328 VSS.n8393 VSS.n8392 8.0005
R4329 VSS.n8251 VSS.n8250 8.0005
R4330 VSS.n6759 VSS.n6716 8.0005
R4331 VSS.n9956 VSS.n9955 8.0005
R4332 VSS.n8026 VSS.n8025 8.0005
R4333 VSS.n8112 VSS.n8096 8.0005
R4334 VSS.n8891 VSS.n7973 8.0005
R4335 VSS.n8854 VSS.n8852 8.0005
R4336 VSS.n8269 VSS.n8268 8.0005
R4337 VSS.n9584 VSS.n9580 8.0005
R4338 VSS.n9275 VSS.n9273 8.0005
R4339 VSS.n9496 VSS.n9492 8.0005
R4340 VSS.n9472 VSS.n9470 8.0005
R4341 VSS.n9814 VSS.n9813 8.0005
R4342 VSS.n7354 VSS.n7353 8.0005
R4343 VSS.n7201 VSS.n7198 8.0005
R4344 VSS.n9173 VSS.n9172 8.0005
R4345 VSS.n9196 VSS.n9192 8.0005
R4346 VSS.n7901 VSS.n7898 8.0005
R4347 VSS.n7833 VSS.n7832 8.0005
R4348 VSS.n7625 VSS.n7624 8.0005
R4349 VSS.n7787 VSS.n7786 8.0005
R4350 VSS.n7660 VSS.n7659 8.0005
R4351 VSS.n7708 VSS.n7707 8.0005
R4352 VSS.n7123 VSS.n7122 8.0005
R4353 VSS.n9871 VSS.n9870 8.0005
R4354 VSS.n7923 VSS.n7922 8.0005
R4355 VSS.n7985 VSS.n7980 8.0005
R4356 VSS.n6798 VSS.n6796 8.0005
R4357 VSS.n6886 VSS.n6885 8.0005
R4358 VSS.n6866 VSS.n6864 8.0005
R4359 VSS.n6959 VSS.n6958 8.0005
R4360 VSS.n6936 VSS.n6933 8.0005
R4361 VSS.n7003 VSS.n7002 8.0005
R4362 VSS.n7019 VSS.n7017 8.0005
R4363 VSS.n6279 VSS.n6278 8.0005
R4364 VSS.n6408 VSS.n6407 8.0005
R4365 VSS.n6433 VSS.n6432 8.0005
R4366 VSS.n6819 VSS.n6818 8.0005
R4367 VSS.n6723 VSS.n6720 8.0005
R4368 VSS.n6339 VSS.n6338 8.0005
R4369 VSS.n11012 VSS.n11011 8.0005
R4370 VSS.n10972 VSS.n10971 8.0005
R4371 VSS.n10905 VSS.n10903 8.0005
R4372 VSS.n7285 VSS.n7284 8.0005
R4373 VSS.n10861 VSS.n10860 8.0005
R4374 VSS.n4387 VSS.n4386 8.0005
R4375 VSS.n4282 VSS.n4281 8.0005
R4376 VSS.n4241 VSS.n4240 8.0005
R4377 VSS.n4179 VSS.n4170 8.0005
R4378 VSS.n4123 VSS.n4122 8.0005
R4379 VSS.n10753 VSS.n10752 8.0005
R4380 VSS.n594 VSS.n593 8.0005
R4381 VSS.n14211 VSS.n14210 8.0005
R4382 VSS.n563 VSS.n560 8.0005
R4383 VSS.n1149 VSS.n934 8.0005
R4384 VSS.n13032 VSS.n13031 8.0005
R4385 VSS.n2471 VSS.n2468 8.0005
R4386 VSS.n2436 VSS.n2433 8.0005
R4387 VSS.n2367 VSS.n2366 8.0005
R4388 VSS.n2340 VSS.n1944 8.0005
R4389 VSS.n13112 VSS.n13111 8.0005
R4390 VSS.n940 VSS.n939 8.0005
R4391 VSS.n1378 VSS.n1374 8.0005
R4392 VSS.n1445 VSS.n1443 8.0005
R4393 VSS.n14095 VSS.n14091 8.0005
R4394 VSS.n1655 VSS.n1654 8.0005
R4395 VSS.n13657 VSS.n13655 8.0005
R4396 VSS.n13630 VSS.n13629 8.0005
R4397 VSS.n13882 VSS.n13881 8.0005
R4398 VSS.n826 VSS.n825 8.0005
R4399 VSS.n1180 VSS.n1179 8.0005
R4400 VSS.n2039 VSS.n2037 8.0005
R4401 VSS.n2221 VSS.n2220 8.0005
R4402 VSS.n2088 VSS.n2086 8.0005
R4403 VSS.n2156 VSS.n2155 8.0005
R4404 VSS.n2136 VSS.n2134 8.0005
R4405 VSS.n1839 VSS.n1838 8.0005
R4406 VSS.n1788 VSS.n1787 8.0005
R4407 VSS.n1822 VSS.n1821 8.0005
R4408 VSS.n2016 VSS.n2014 8.0005
R4409 VSS.n1960 VSS.n1957 8.0005
R4410 VSS.n2646 VSS.n2644 8.0005
R4411 VSS.n12961 VSS.n12960 8.0005
R4412 VSS.n2682 VSS.n2681 8.0005
R4413 VSS.n2778 VSS.n2773 8.0005
R4414 VSS.n2827 VSS.n2825 8.0005
R4415 VSS.n12884 VSS.n12883 8.0005
R4416 VSS.n2862 VSS.n2861 8.0005
R4417 VSS.n3041 VSS.n3039 8.0005
R4418 VSS.n2966 VSS.n2965 8.0005
R4419 VSS.n3027 VSS.n3026 8.0005
R4420 VSS.n2596 VSS.n2594 8.0005
R4421 VSS.n2512 VSS.n2509 8.0005
R4422 VSS.n12741 VSS.n12740 8.0005
R4423 VSS.n12766 VSS.n12765 8.0005
R4424 VSS.n13947 VSS.n13946 8.0005
R4425 VSS.n1727 VSS.n1726 8.0005
R4426 VSS.n13563 VSS.n13562 8.0005
R4427 VSS.n13492 VSS.n13491 8.0005
R4428 VSS VSS.n11252 6.77697
R4429 VSS.n3656 VSS 6.77697
R4430 VSS.n3666 VSS 6.77697
R4431 VSS.n11242 VSS 6.77697
R4432 VSS.n11485 VSS.n11476 6.32234
R4433 VSS.n11422 VSS.n11421 5.57294
R4434 VSS.n11413 VSS 4.68305
R4435 VSS.n3675 VSS 4.67264
R4436 VSS.n11232 VSS 4.67264
R4437 VSS.n11411 VSS.n3688 4.6505
R4438 VSS.n11392 VSS.n3689 4.6505
R4439 VSS.n11391 VSS.n3690 4.6505
R4440 VSS.n11374 VSS.n3691 4.6505
R4441 VSS.n11373 VSS.n3692 4.6505
R4442 VSS.n11358 VSS.n11357 4.6505
R4443 VSS.n11355 VSS.n3694 4.6505
R4444 VSS.n11354 VSS.n3695 4.6505
R4445 VSS.n11410 VSS.n11409 4.6505
R4446 VSS.n11408 VSS.n11407 4.6505
R4447 VSS.n11406 VSS.n11405 4.6505
R4448 VSS.n11404 VSS.n11403 4.6505
R4449 VSS.n11402 VSS.n11401 4.6505
R4450 VSS.n11400 VSS.n11399 4.6505
R4451 VSS.n11398 VSS.n11397 4.6505
R4452 VSS.n11396 VSS.n11395 4.6505
R4453 VSS.n11394 VSS.n11393 4.6505
R4454 VSS.n11390 VSS.n11389 4.6505
R4455 VSS.n11388 VSS.n11387 4.6505
R4456 VSS.n11386 VSS.n11385 4.6505
R4457 VSS.n11384 VSS.n11383 4.6505
R4458 VSS.n11382 VSS.n11381 4.6505
R4459 VSS.n11380 VSS.n11379 4.6505
R4460 VSS.n11378 VSS.n11377 4.6505
R4461 VSS.n11376 VSS.n11375 4.6505
R4462 VSS.n11372 VSS.n11371 4.6505
R4463 VSS.n11370 VSS.n11369 4.6505
R4464 VSS.n11368 VSS.n11367 4.6505
R4465 VSS.n11366 VSS.n11365 4.6505
R4466 VSS.n11364 VSS.n11363 4.6505
R4467 VSS.n11362 VSS.n11361 4.6505
R4468 VSS.n11360 VSS.n11359 4.6505
R4469 VSS.n11356 VSS.n3693 4.6505
R4470 VSS.n11353 VSS.n11352 4.6505
R4471 VSS.n11351 VSS.n11350 4.6505
R4472 VSS.n11412 VSS.n3686 4.6505
R4473 VSS.n11349 VSS.n11344 4.6505
R4474 VSS.n3664 VSS.n3642 4.6505
R4475 VSS.n3661 VSS.n3643 4.6505
R4476 VSS.n3655 VSS.n3654 4.6505
R4477 VSS.n3651 VSS.n3645 4.6505
R4478 VSS.n3674 VSS.n3640 4.6505
R4479 VSS.n3673 VSS.n3672 4.6505
R4480 VSS.n3671 VSS.n3670 4.6505
R4481 VSS.n3669 VSS.n3641 4.6505
R4482 VSS.n3668 VSS.n3667 4.6505
R4483 VSS.n3666 VSS.n3665 4.6505
R4484 VSS.n3663 VSS.n3662 4.6505
R4485 VSS.n3660 VSS.n3659 4.6505
R4486 VSS.n3658 VSS.n3644 4.6505
R4487 VSS.n3657 VSS.n3656 4.6505
R4488 VSS.n3653 VSS.n3652 4.6505
R4489 VSS.n3650 VSS.n3649 4.6505
R4490 VSS.n3648 VSS.n3647 4.6505
R4491 VSS.n3646 VSS.n3639 4.6505
R4492 VSS.n11246 VSS.n11245 4.6505
R4493 VSS.n11247 VSS.n11217 4.6505
R4494 VSS.n11253 VSS.n11215 4.6505
R4495 VSS.n11256 VSS.n11255 4.6505
R4496 VSS.n11249 VSS.n11248 4.6505
R4497 VSS.n11250 VSS.n11216 4.6505
R4498 VSS.n11252 VSS.n11251 4.6505
R4499 VSS.n11254 VSS.n11214 4.6505
R4500 VSS.n11257 VSS.n11213 4.6505
R4501 VSS.n11259 VSS.n11258 4.6505
R4502 VSS.n11260 VSS.n11212 4.6505
R4503 VSS.n11244 VSS.n11218 4.6505
R4504 VSS.n11239 VSS.n11238 4.6505
R4505 VSS.n11241 VSS.n11240 4.6505
R4506 VSS.n11243 VSS.n11242 4.6505
R4507 VSS.n11234 VSS.n11233 4.6505
R4508 VSS.n11235 VSS.n11219 4.6505
R4509 VSS.n11237 VSS.n11236 4.6505
R4510 VSS.n3628 VSS.n3627 4.61383
R4511 VSS.n3627 VSS.n3626 4.61383
R4512 VSS.n11322 VSS.n11321 4.61383
R4513 VSS.n11323 VSS.n11322 4.61383
R4514 VSS.n11283 VSS.n11280 4.4948
R4515 VSS.n11307 VSS.n11306 4.4948
R4516 VSS.n11425 VSS.n3676 4.47386
R4517 VSS.n12550 VSS.n3373 4.4066
R4518 VSS.n5394 VSS.n4706 4.4066
R4519 VSS.n6133 VSS 4.4066
R4520 VSS.n6117 VSS 4.4066
R4521 VSS.n5951 VSS 4.4066
R4522 VSS.n5935 VSS 4.4066
R4523 VSS.n5770 VSS 4.4066
R4524 VSS.n5754 VSS 4.4066
R4525 VSS.n5590 VSS 4.4066
R4526 VSS.n5574 VSS 4.4066
R4527 VSS.n5410 VSS 4.4066
R4528 VSS.n5230 VSS 4.4066
R4529 VSS.n5214 VSS 4.4066
R4530 VSS.n10117 VSS 4.4066
R4531 VSS VSS.n10162 4.4066
R4532 VSS.n11160 VSS 4.4066
R4533 VSS.n11176 VSS 4.4066
R4534 VSS VSS.n12296 4.4066
R4535 VSS.n12319 VSS 4.4066
R4536 VSS VSS.n12478 4.4066
R4537 VSS.n12176 VSS 4.4066
R4538 VSS.n12194 VSS 4.4066
R4539 VSS.n14488 VSS 4.4066
R4540 VSS VSS.n14485 4.4066
R4541 VSS VSS.n3318 4.4066
R4542 VSS.n12559 VSS 4.4066
R4543 VSS.n3410 VSS 4.4066
R4544 VSS VSS.n3585 4.4066
R4545 VSS.n11895 VSS 4.4066
R4546 VSS.n12009 VSS 4.4066
R4547 VSS.n12026 VSS 4.4066
R4548 VSS.n11560 VSS 4.39702
R4549 VSS.n14032 VSS.n14028 4.11196
R4550 VSS.n13999 VSS.n1751 4.11196
R4551 VSS.n12833 VSS.n12829 4.11196
R4552 VSS.n12999 VSS.n12998 4.11196
R4553 VSS.n2733 VSS.n2728 4.11196
R4554 VSS.n12921 VSS.n2736 4.11196
R4555 VSS.n2913 VSS.n2908 4.11196
R4556 VSS.n12844 VSS.n2916 4.11196
R4557 VSS.n13157 VSS.n1898 4.11196
R4558 VSS.n13166 VSS.n1894 4.11196
R4559 VSS.n13173 VSS.n1888 4.11196
R4560 VSS.n13177 VSS.n1886 4.11196
R4561 VSS.n14132 VSS.n14128 4.11196
R4562 VSS.n14050 VSS.n14045 4.11196
R4563 VSS.n14054 VSS.n14043 4.11196
R4564 VSS.n10959 VSS.n3888 4.11196
R4565 VSS.n11003 VSS.n3845 4.11196
R4566 VSS.n11118 VSS.n3820 4.11196
R4567 VSS.n9997 VSS.n4654 4.11196
R4568 VSS.n10006 VSS.n4650 4.11196
R4569 VSS.n10015 VSS.n4646 4.11196
R4570 VSS.n10024 VSS.n4642 4.11196
R4571 VSS.n10031 VSS.n4636 4.11196
R4572 VSS.n9935 VSS.n9934 4.11196
R4573 VSS.n9929 VSS.n9926 4.11196
R4574 VSS.n9921 VSS.n9918 4.11196
R4575 VSS.n9913 VSS.n9910 4.11196
R4576 VSS.n9533 VSS.n9529 4.11196
R4577 VSS.n7606 VSS.n7603 4.11196
R4578 VSS.n9854 VSS.n7150 4.11196
R4579 VSS.n4355 VSS.n4205 4.11196
R4580 VSS.n9988 VSS.n4658 4.11196
R4581 VSS.n9947 VSS.n9946 4.11196
R4582 VSS.n9941 VSS.n9940 4.11196
R4583 VSS.n8837 VSS.n8012 4.11196
R4584 VSS.n8842 VSS.n8841 4.11196
R4585 VSS.n9539 VSS.n7595 4.11196
R4586 VSS.n9860 VSS.n9858 4.11196
R4587 VSS.n9907 VSS.n9905 4.11196
R4588 VSS.n10037 VSS.n10035 4.11196
R4589 VSS.n4438 VSS.n4157 4.11196
R4590 VSS.n12428 VSS.n12427 4.11196
R4591 VSS.n13064 VSS.n13063 4.11196
R4592 VSS.n13148 VSS.n1902 4.11196
R4593 VSS.n2426 VSS.n2425 4.11196
R4594 VSS.n14147 VSS.n14146 4.11196
R4595 VSS.n14141 VSS.n14138 4.11196
R4596 VSS.n14040 VSS.n14038 4.11196
R4597 VSS.n12704 VSS.n12702 4.11196
R4598 VSS.n12841 VSS.n12839 4.11196
R4599 VSS.n8516 VSS.n8515 3.89651
R4600 VSS.n9988 VSS.n9987 3.89651
R4601 VSS.n9946 VSS.n6235 3.89651
R4602 VSS.n9940 VSS.n6240 3.89651
R4603 VSS.n8837 VSS.n8836 3.89651
R4604 VSS.n8841 VSS.n8839 3.89651
R4605 VSS.n9541 VSS.n9539 3.89651
R4606 VSS.n9858 VSS.n9857 3.89651
R4607 VSS.n9854 VSS.n9853 3.89651
R4608 VSS.n7603 VSS.n7602 3.89651
R4609 VSS.n9529 VSS.n7598 3.89651
R4610 VSS.n9905 VSS.n9904 3.89651
R4611 VSS.n9910 VSS.n6264 3.89651
R4612 VSS.n9918 VSS.n6259 3.89651
R4613 VSS.n9926 VSS.n6254 3.89651
R4614 VSS.n9934 VSS.n6247 3.89651
R4615 VSS.n10035 VSS.n10034 3.89651
R4616 VSS.n10031 VSS.n10030 3.89651
R4617 VSS.n10024 VSS.n10023 3.89651
R4618 VSS.n10015 VSS.n10014 3.89651
R4619 VSS.n10006 VSS.n10005 3.89651
R4620 VSS.n9997 VSS.n9996 3.89651
R4621 VSS.n11120 VSS.n11118 3.89651
R4622 VSS.n11003 VSS.n11002 3.89651
R4623 VSS.n10961 VSS.n10959 3.89651
R4624 VSS.n10849 VSS.n10848 3.89651
R4625 VSS.n4356 VSS.n4355 3.89651
R4626 VSS.n4438 VSS.n4437 3.89651
R4627 VSS.n14243 VSS.n14242 3.89651
R4628 VSS.n12427 VSS.n12424 3.89651
R4629 VSS.n13065 VSS.n13064 3.89651
R4630 VSS.n13148 VSS.n13147 3.89651
R4631 VSS.n2425 VSS.n2424 3.89651
R4632 VSS.n14146 VSS.n612 3.89651
R4633 VSS.n14138 VSS.n618 3.89651
R4634 VSS.n14038 VSS.n1707 3.89651
R4635 VSS.n14043 VSS.n1701 3.89651
R4636 VSS.n14050 VSS.n14049 3.89651
R4637 VSS.n14128 VSS.n621 3.89651
R4638 VSS.n12702 VSS.n12701 3.89651
R4639 VSS.n1886 VSS.n1885 3.89651
R4640 VSS.n13173 VSS.n13172 3.89651
R4641 VSS.n13166 VSS.n13165 3.89651
R4642 VSS.n13157 VSS.n13156 3.89651
R4643 VSS.n12839 VSS.n2922 3.89651
R4644 VSS.n12846 VSS.n12844 3.89651
R4645 VSS.n2913 VSS.n2912 3.89651
R4646 VSS.n12923 VSS.n12921 3.89651
R4647 VSS.n2733 VSS.n2732 3.89651
R4648 VSS.n12998 VSS.n2553 3.89651
R4649 VSS.n12829 VSS.n2925 3.89651
R4650 VSS.n13999 VSS.n13998 3.89651
R4651 VSS.n14028 VSS.n1710 3.89651
R4652 VSS.n13621 VSS.n13614 3.89651
R4653 VSS.n4331 VSS.n4329 3.71869
R4654 VSS.n6099 VSS.n4663 3.59425
R4655 VSS.n12363 VSS.n12362 3.59425
R4656 VSS VSS.n3605 3.33963
R4657 VSS.n11231 VSS.n11230 3.3223
R4658 VSS.n14375 VSS 3.31776
R4659 VSS.n3282 VSS.n3281 3.12488
R4660 VSS.n980 VSS 2.84776
R4661 VSS.n11500 VSS.n3637 2.52171
R4662 VSS.n1238 VSS 2.37788
R4663 VSS.n5110 VSS 2.37087
R4664 VSS.n5112 VSS 2.37087
R4665 VSS.n5119 VSS 2.37087
R4666 VSS.n5117 VSS 2.37087
R4667 VSS.n5138 VSS 2.37087
R4668 VSS.n4735 VSS 2.37087
R4669 VSS.n5145 VSS 2.37087
R4670 VSS.n4732 VSS 2.37087
R4671 VSS.n5152 VSS 2.37087
R4672 VSS.n5159 VSS 2.37087
R4673 VSS VSS.n5180 2.37087
R4674 VSS.n5179 VSS 2.37087
R4675 VSS.n10163 VSS 2.37087
R4676 VSS.n10169 VSS 2.37087
R4677 VSS.n10173 VSS 2.37087
R4678 VSS.n12297 VSS 2.37087
R4679 VSS VSS.n12308 2.37087
R4680 VSS.n12479 VSS 2.37087
R4681 VSS VSS.n3590 2.37087
R4682 VSS.n12514 VSS 2.37087
R4683 VSS VSS.n14487 2.37087
R4684 VSS.n14486 VSS 2.37087
R4685 VSS.n3319 VSS 2.37087
R4686 VSS VSS.n12552 2.37087
R4687 VSS VSS.n3374 2.37087
R4688 VSS.n12527 VSS 2.37087
R4689 VSS.n12525 VSS 2.37087
R4690 VSS.n12523 VSS 2.37087
R4691 VSS.n12521 VSS 2.37087
R4692 VSS.n11276 VSS 2.00407
R4693 VSS.n8745 VSS.n8744 1.921
R4694 VSS.n9559 VSS.n9558 1.921
R4695 VSS.n8553 VSS.n8552 1.921
R4696 VSS.n7395 VSS.n7394 1.921
R4697 VSS.n3928 VSS.n3927 1.921
R4698 VSS.n9442 VSS.n9441 1.921
R4699 VSS.n9510 VSS.n9316 1.921
R4700 VSS.n9832 VSS.n7185 1.921
R4701 VSS.n9245 VSS.n9244 1.921
R4702 VSS.n8952 VSS.n8951 1.921
R4703 VSS.n7805 VSS.n7641 1.921
R4704 VSS.n7726 VSS.n7700 1.921
R4705 VSS.n8927 VSS.n8926 1.921
R4706 VSS.n6905 VSS.n6904 1.921
R4707 VSS.n6978 VSS.n6977 1.921
R4708 VSS.n7000 VSS.n6999 1.921
R4709 VSS.n7059 VSS.n7058 1.921
R4710 VSS.n6838 VSS.n6791 1.921
R4711 VSS.n5886 VSS.n5885 1.921
R4712 VSS.n5705 VSS.n5704 1.921
R4713 VSS.n5525 VSS.n5524 1.921
R4714 VSS.n5345 VSS.n5344 1.921
R4715 VSS.n10079 VSS.n10078 1.921
R4716 VSS.n6077 VSS.n6076 1.921
R4717 VSS.n4383 VSS.n4197 1.921
R4718 VSS.n1338 VSS.n1337 1.921
R4719 VSS.n582 VSS.n579 1.921
R4720 VSS.n1393 VSS.n1392 1.921
R4721 VSS.n957 VSS.n956 1.921
R4722 VSS.n13715 VSS.n13714 1.921
R4723 VSS.n13255 VSS.n13254 1.921
R4724 VSS.n1609 VSS.n1608 1.921
R4725 VSS.n14109 VSS.n1462 1.921
R4726 VSS.n13696 VSS.n13695 1.921
R4727 VSS.n1415 VSS.n1414 1.921
R4728 VSS.n2239 VSS.n2212 1.921
R4729 VSS.n2174 VSS.n2128 1.921
R4730 VSS.n13194 VSS.n13193 1.921
R4731 VSS.n2277 VSS.n1978 1.921
R4732 VSS.n12979 VSS.n2662 1.921
R4733 VSS.n2813 VSS.n2812 1.921
R4734 VSS.n12902 VSS.n2843 1.921
R4735 VSS.n12637 VSS.n12636 1.921
R4736 VSS.n2633 VSS.n2632 1.921
R4737 VSS.n12247 VSS.n12246 1.921
R4738 VSS.n12140 VSS.n12139 1.921
R4739 VSS.n11972 VSS.n11971 1.921
R4740 VSS.n3544 VSS.n3543 1.921
R4741 VSS.n12596 VSS.n12595 1.921
R4742 VSS.n11627 VSS.n11626 1.921
R4743 VSS.n9023 VSS.n9022 1.9205
R4744 VSS.n7524 VSS.n7523 1.9205
R4745 VSS.n8781 VSS.n8780 1.9205
R4746 VSS.n6742 VSS.n6740 1.9205
R4747 VSS.n8118 VSS.n8117 1.9205
R4748 VSS.n8874 VSS.n8872 1.9205
R4749 VSS.n8819 VSS.n8818 1.9205
R4750 VSS.n7371 VSS.n7370 1.9205
R4751 VSS.n7141 VSS.n7140 1.9205
R4752 VSS.n6425 VSS.n6424 1.9205
R4753 VSS.n3757 VSS.n3756 1.9205
R4754 VSS.n11071 VSS.n11070 1.9205
R4755 VSS.n11028 VSS.n3838 1.9205
R4756 VSS.n10919 VSS.n10917 1.9205
R4757 VSS.n10877 VSS.n3906 1.9205
R4758 VSS.n4054 VSS.n4053 1.9205
R4759 VSS.n4270 VSS.n4269 1.9205
R4760 VSS.n10771 VSS.n4133 1.9205
R4761 VSS.n656 VSS.n655 1.9205
R4762 VSS.n512 VSS.n511 1.9205
R4763 VSS.n1132 VSS.n604 1.9205
R4764 VSS.n13049 VSS.n13048 1.9205
R4765 VSS.n13096 VSS.n13095 1.9205
R4766 VSS.n2346 VSS.n2345 1.9205
R4767 VSS.n13647 VSS.n13646 1.9205
R4768 VSS.n13930 VSS.n13929 1.9205
R4769 VSS.n12725 VSS.n12724 1.9205
R4770 VSS.n3220 VSS.n3219 1.9205
R4771 VSS.n12782 VSS.n12760 1.9205
R4772 VSS.n1767 VSS.n1766 1.9205
R4773 VSS.n13586 VSS.n13585 1.9205
R4774 VSS.n13451 VSS.n13450 1.9205
R4775 VSS.n700 VSS 1.90776
R4776 VSS.n12807 VSS.n12806 1.87823
R4777 VSS.n11487 VSS 1.85727
R4778 VSS.n9663 VSS.n9662 1.84989
R4779 VSS.n8675 VSS.n8674 1.84989
R4780 VSS.n8783 VSS.n8782 1.84989
R4781 VSS.n9975 VSS.n6231 1.84989
R4782 VSS.n8149 VSS.n8148 1.84989
R4783 VSS.n8871 VSS.n8002 1.84989
R4784 VSS.n8821 VSS.n8820 1.84989
R4785 VSS.n7373 VSS.n7372 1.84989
R4786 VSS.n9890 VSS.n7142 1.84989
R4787 VSS.n6452 VSS.n6426 1.84989
R4788 VSS.n4606 VSS.n4605 1.84989
R4789 VSS.n3718 VSS.n3717 1.84989
R4790 VSS.n6394 VSS.n6393 1.84989
R4791 VSS.n3880 VSS.n3877 1.84989
R4792 VSS.n7340 VSS.n7339 1.84989
R4793 VSS.n4015 VSS.n4014 1.84989
R4794 VSS.n4301 VSS.n4271 1.84989
R4795 VSS.n10772 VSS.n4128 1.84989
R4796 VSS.n1268 VSS.n1267 1.84989
R4797 VSS.n10694 VSS.n10693 1.84989
R4798 VSS.n14199 VSS.n14198 1.84989
R4799 VSS.n13051 VSS.n13050 1.84989
R4800 VSS.n13092 VSS.n2454 1.84989
R4801 VSS.n13131 VSS.n2347 1.84989
R4802 VSS.n13901 VSS.n13648 1.84989
R4803 VSS.n13926 VSS.n1814 1.84989
R4804 VSS.n12721 VSS.n3019 1.84989
R4805 VSS.n3140 VSS.n3139 1.84989
R4806 VSS.n12759 VSS.n12758 1.84989
R4807 VSS.n13966 VSS.n1768 1.84989
R4808 VSS.n13582 VSS.n13581 1.84989
R4809 VSS.n13298 VSS.n13297 1.84989
R4810 VSS.n3282 VSS.n3279 1.84939
R4811 VSS.n8568 VSS.n8567 1.84939
R4812 VSS.n9557 VSS.n9556 1.84939
R4813 VSS.n8460 VSS.n8459 1.84939
R4814 VSS.n9368 VSS.n9367 1.84939
R4815 VSS.n7424 VSS.n7423 1.84939
R4816 VSS.n9061 VSS.n9060 1.84939
R4817 VSS.n9512 VSS.n9511 1.84939
R4818 VSS.n9834 VSS.n9833 1.84939
R4819 VSS.n9243 VSS.n9242 1.84939
R4820 VSS.n8950 VSS.n8949 1.84939
R4821 VSS.n7806 VSS.n7639 1.84939
R4822 VSS.n7727 VSS.n7674 1.84939
R4823 VSS.n8925 VSS.n8924 1.84939
R4824 VSS.n6858 VSS.n6857 1.84939
R4825 VSS.n6925 VSS.n6924 1.84939
R4826 VSS.n6998 VSS.n6997 1.84939
R4827 VSS.n7057 VSS.n7056 1.84939
R4828 VSS.n6790 VSS.n6789 1.84939
R4829 VSS.n5995 VSS.n5994 1.84939
R4830 VSS.n5796 VSS.n5795 1.84939
R4831 VSS.n5615 VSS.n5614 1.84939
R4832 VSS.n5436 VSS.n5435 1.84939
R4833 VSS.n5255 VSS.n5254 1.84939
R4834 VSS.n6181 VSS.n6180 1.84939
R4835 VSS.n4382 VSS.n4381 1.84939
R4836 VSS.n1000 VSS.n999 1.84939
R4837 VSS.n2400 VSS.n2398 1.84939
R4838 VSS.n1169 VSS.n1168 1.84939
R4839 VSS.n14304 VSS.n14303 1.84939
R4840 VSS.n1521 VSS.n1520 1.84939
R4841 VSS.n13761 VSS.n13760 1.84939
R4842 VSS.n715 VSS.n714 1.84939
R4843 VSS.n14111 VSS.n14110 1.84939
R4844 VSS.n1670 VSS.n1669 1.84939
R4845 VSS.n1413 VSS.n1412 1.84939
R4846 VSS.n2241 VSS.n2240 1.84939
R4847 VSS.n2176 VSS.n2175 1.84939
R4848 VSS.n13192 VSS.n13191 1.84939
R4849 VSS.n2278 VSS.n1976 1.84939
R4850 VSS.n12981 VSS.n12980 1.84939
R4851 VSS.n2697 VSS.n2696 1.84939
R4852 VSS.n12904 VSS.n12903 1.84939
R4853 VSS.n2877 VSS.n2876 1.84939
R4854 VSS.n2529 VSS.n2528 1.84939
R4855 VSS.n11574 VSS.n11573 1.84939
R4856 VSS.n11697 VSS.n11696 1.84939
R4857 VSS.n12050 VSS.n12049 1.84939
R4858 VSS.n11829 VSS.n11828 1.84939
R4859 VSS.n3454 VSS.n3453 1.84939
R4860 VSS.n12386 VSS.n12385 1.84939
R4861 VSS VSS 1.84247
R4862 VSS.n3629 VSS.n3628 1.79444
R4863 VSS.n11313 VSS.n11303 1.74595
R4864 VSS VSS 1.57079
R4865 VSS.n11287 VSS.n11284 1.45505
R4866 VSS.n1501 VSS 1.43788
R4867 VSS.n3628 VSS.n3625 1.35808
R4868 VSS VSS 1.29911
R4869 VSS VSS.n10631 1.11354
R4870 VSS.n10630 VSS 1.11354
R4871 VSS VSS 1.02744
R4872 VSS.n5111 VSS.n5110 0.976535
R4873 VSS.n5113 VSS.n5112 0.976535
R4874 VSS.n5119 VSS.n5118 0.976535
R4875 VSS.n5117 VSS.n4738 0.976535
R4876 VSS.n5139 VSS.n5138 0.976535
R4877 VSS.n5140 VSS.n4735 0.976535
R4878 VSS.n5146 VSS.n5145 0.976535
R4879 VSS.n5147 VSS.n4732 0.976535
R4880 VSS.n5153 VSS.n5152 0.976535
R4881 VSS.n5159 VSS.n5158 0.976535
R4882 VSS.n5180 VSS.n4718 0.976535
R4883 VSS.n5179 VSS.n5178 0.976535
R4884 VSS.n10163 VSS.n4563 0.976535
R4885 VSS.n10170 VSS.n10169 0.976535
R4886 VSS.n10173 VSS.n10172 0.976535
R4887 VSS.n12297 VSS.n3594 0.976535
R4888 VSS.n12308 VSS.n12298 0.976535
R4889 VSS.n12480 VSS.n12479 0.976535
R4890 VSS.n12516 VSS.n3590 0.976535
R4891 VSS.n12515 VSS.n12514 0.976535
R4892 VSS.n14487 VSS.n20 0.976535
R4893 VSS.n14486 VSS.n21 0.976535
R4894 VSS.n10541 VSS.n3319 0.976535
R4895 VSS.n12552 VSS.n12551 0.976535
R4896 VSS.n12529 VSS.n3374 0.976535
R4897 VSS.n12528 VSS.n12527 0.976535
R4898 VSS.n12526 VSS.n12525 0.976535
R4899 VSS.n12524 VSS.n12523 0.976535
R4900 VSS.n12522 VSS.n12521 0.976535
R4901 VSS.n13750 VSS 0.967877
R4902 VSS.n10802 VSS.n10801 0.95507
R4903 VSS.n11319 VSS.n11318 0.921712
R4904 VSS.n11500 VSS.n11493 0.921712
R4905 VSS.n11323 VSS.n11319 0.824742
R4906 VSS VSS 0.75576
R4907 VSS VSS.n11343 0.741385
R4908 VSS.n11193 VSS.n11192 0.614203
R4909 VSS.n11514 VSS.n11513 0.542292
R4910 VSS.n13288 VSS 0.497878
R4911 VSS VSS 0.484084
R4912 VSS.n6100 VSS 0.426857
R4913 VSS.n5918 VSS 0.426857
R4914 VSS.n11488 VSS 0.424356
R4915 VSS.n5197 VSS 0.39425
R4916 VSS.n10145 VSS 0.389562
R4917 VSS.n5737 VSS 0.383312
R4918 VSS.n3299 VSS 0.380708
R4919 VSS.n5 VSS 0.380708
R4920 VSS.n5377 VSS 0.380187
R4921 VSS.n11814 VSS 0.379146
R4922 VSS.n8340 VSS 0.3755
R4923 VSS.n8322 VSS 0.3755
R4924 VSS.n7517 VSS 0.3755
R4925 VSS.n9726 VSS 0.3755
R4926 VSS.n5557 VSS 0.369771
R4927 VSS.n3957 VSS 0.368208
R4928 VSS.n11797 VSS 0.361958
R4929 VSS.n10808 VSS.n10804 0.352765
R4930 VSS.n691 VSS 0.352583
R4931 VSS.n3331 VSS 0.346333
R4932 VSS.n9355 VSS 0.341646
R4933 VSS.n10787 VSS.n10786 0.340206
R4934 VSS.n10744 VSS.n10742 0.339716
R4935 VSS.n12274 VSS 0.339563
R4936 VSS.n3385 VSS 0.336958
R4937 VSS.n10725 VSS.n10724 0.334553
R4938 VSS.n12361 VSS 0.330188
R4939 VSS.n9738 VSS.n9737 0.329265
R4940 VSS.n994 VSS 0.3255
R4941 VSS.n9754 VSS.n9753 0.324095
R4942 VSS.n13426 VSS 0.322896
R4943 VSS.n1515 VSS 0.322896
R4944 VSS.n13756 VSS 0.322896
R4945 VSS.n13293 VSS 0.322896
R4946 VSS.n10744 VSS 0.318729
R4947 VSS.n1245 VSS 0.317167
R4948 VSS.n8420 VSS.n8417 0.315283
R4949 VSS.n8646 VSS.n8645 0.315283
R4950 VSS.n8719 VSS.n8715 0.315283
R4951 VSS.n9721 VSS.n9720 0.315283
R4952 VSS.n7482 VSS 0.313
R4953 VSS.n9765 VSS.n9761 0.310818
R4954 VSS.n14370 VSS 0.304667
R4955 VSS.n11284 VSS.n11279 0.291409
R4956 VSS.n11303 VSS.n11302 0.291409
R4957 VSS.n10786 VSS 0.284875
R4958 VSS.n11277 VSS 0.278917
R4959 VSS.n11186 VSS 0.278625
R4960 VSS.n12339 VSS 0.265604
R4961 VSS.n4332 VSS.n4331 0.252499
R4962 VSS.n11082 VSS.n11081 0.25175
R4963 VSS.n12815 VSS.n12814 0.25175
R4964 VSS.n11325 VSS.n11324 0.247667
R4965 VSS.n11143 VSS 0.247375
R4966 VSS.n11503 VSS.n11502 0.24733
R4967 VSS.n12042 VSS 0.246854
R4968 VSS.n1324 VSS 0.242435
R4969 VSS.n9116 VSS 0.235396
R4970 VSS.n10100 VSS 0.234354
R4971 VSS.n12206 VSS 0.234354
R4972 VSS.n6155 VSS.n6154 0.232887
R4973 VSS.n4325 VSS.n4324 0.232887
R4974 VSS.n12459 VSS.n12458 0.232887
R4975 VSS.n5605 VSS 0.228104
R4976 VSS.n4028 VSS 0.226021
R4977 VSS.n12579 VSS 0.226021
R4978 VSS.n3212 VSS 0.226021
R4979 VSS.n12463 VSS 0.221854
R4980 VSS.n10715 VSS 0.221854
R4981 VSS VSS 0.212408
R4982 VSS.n3444 VSS 0.210917
R4983 VSS.n5245 VSS 0.209875
R4984 VSS.n8429 VSS 0.207271
R4985 VSS.n8625 VSS 0.207271
R4986 VSS.n8711 VSS 0.207271
R4987 VSS.n9700 VSS 0.207271
R4988 VSS.n11929 VSS 0.204146
R4989 VSS.n1074 VSS 0.203203
R4990 VSS.n5425 VSS 0.201542
R4991 VSS.n6150 VSS 0.186437
R4992 VSS.n5967 VSS 0.186437
R4993 VSS.n5786 VSS 0.185396
R4994 VSS.n9424 VSS 0.183833
R4995 VSS.n14360 VSS 0.181229
R4996 VSS.n9770 VSS 0.180188
R4997 VSS.n463 VSS 0.178625
R4998 VSS.n13371 VSS 0.178625
R4999 VSS.n13836 VSS 0.178625
R5000 VSS.n1596 VSS 0.178625
R5001 VSS.n5400 VSS.n5399 0.174048
R5002 VSS.n10612 VSS.n10611 0.17393
R5003 VSS.n6123 VSS.n6122 0.17393
R5004 VSS.n5941 VSS.n5940 0.17393
R5005 VSS.n11166 VSS.n11165 0.17393
R5006 VSS.n12016 VSS.n12015 0.17393
R5007 VSS.n5760 VSS.n5759 0.173813
R5008 VSS.n5580 VSS.n5579 0.173813
R5009 VSS.n5220 VSS.n5219 0.173813
R5010 VSS.n10123 VSS.n10122 0.173813
R5011 VSS.n12184 VSS.n12183 0.173813
R5012 VSS.n1596 VSS 0.172914
R5013 VSS.n463 VSS 0.172914
R5014 VSS.n13836 VSS 0.172914
R5015 VSS.n13371 VSS 0.172914
R5016 VSS.n1074 VSS 0.171854
R5017 VSS.n4089 VSS.n4032 0.169915
R5018 VSS.n8488 VSS.n8487 0.168417
R5019 VSS.n9984 VSS.n9983 0.168417
R5020 VSS.n8125 VSS.n8124 0.168417
R5021 VSS.n8833 VSS.n8832 0.168417
R5022 VSS.n4360 VSS.n4359 0.168417
R5023 VSS.n4434 VSS.n4433 0.168417
R5024 VSS.n10697 VSS.n10696 0.168417
R5025 VSS.n12421 VSS.n12420 0.168417
R5026 VSS.n13069 VSS.n13068 0.168417
R5027 VSS.n2421 VSS.n2420 0.168417
R5028 VSS.n8433 VSS.n8432 0.167667
R5029 VSS.n10783 VSS.n4106 0.167667
R5030 VSS.n10747 VSS.n10746 0.167667
R5031 VSS.n10712 VSS.n10710 0.167667
R5032 VSS.n13429 VSS.n13428 0.167667
R5033 VSS.n13479 VSS.n13478 0.167667
R5034 VSS.n13591 VSS.n1714 0.167667
R5035 VSS.n14004 VSS.n14003 0.167667
R5036 VSS.n12803 VSS.n12802 0.167667
R5037 VSS.n4058 VSS.n3908 0.167667
R5038 VSS.n10898 VSS.n10897 0.167667
R5039 VSS.n10921 VSS.n3840 0.167667
R5040 VSS.n11049 VSS.n11048 0.167667
R5041 VSS.n4443 VSS.n4442 0.167667
R5042 VSS.n4228 VSS.n4225 0.167667
R5043 VSS.n9770 VSS 0.167167
R5044 VSS.n4328 VSS.n4327 0.167167
R5045 VSS.n1324 VSS 0.165604
R5046 VSS.n4325 VSS.n4260 0.16503
R5047 VSS.n14360 VSS 0.163543
R5048 VSS.n9424 VSS 0.155139
R5049 VSS.n13597 VSS.n13592 0.154349
R5050 VSS.n14010 VSS.n14005 0.154349
R5051 VSS.n12791 VSS.n12790 0.154349
R5052 VSS.n2620 VSS.n2613 0.154349
R5053 VSS.n2885 VSS.n2884 0.154349
R5054 VSS.n2802 VSS.n2794 0.154349
R5055 VSS.n2265 VSS.n2258 0.154349
R5056 VSS.n1423 VSS.n1418 0.154349
R5057 VSS.n10886 VSS.n10885 0.154349
R5058 VSS.n10931 VSS.n10930 0.154349
R5059 VSS.n11037 VSS.n11036 0.154349
R5060 VSS.n6666 VSS.n6665 0.154349
R5061 VSS.n6570 VSS.n6569 0.154349
R5062 VSS.n7883 VSS.n7882 0.154349
R5063 VSS.n9253 VSS.n9248 0.154349
R5064 VSS.n9572 VSS.n7562 0.154349
R5065 VSS.n8172 VSS.n8171 0.154349
R5066 VSS.n8204 VSS.n8203 0.154349
R5067 VSS.n8229 VSS.n8228 0.154349
R5068 VSS.n6225 VSS.n6219 0.154349
R5069 VSS.n6705 VSS.n6704 0.154349
R5070 VSS.n8134 VSS.n8133 0.154349
R5071 VSS.n8077 VSS.n8076 0.154349
R5072 VSS.n8056 VSS.n8055 0.154349
R5073 VSS.n7962 VSS.n7961 0.154349
R5074 VSS.n8801 VSS.n8796 0.154349
R5075 VSS.n7579 VSS.n7574 0.154349
R5076 VSS.n9304 VSS.n9297 0.154349
R5077 VSS.n9010 VSS.n9009 0.154349
R5078 VSS.n7230 VSS.n7217 0.154349
R5079 VSS.n7174 VSS.n7173 0.154349
R5080 VSS.n7251 VSS.n7243 0.154349
R5081 VSS.n7320 VSS.n7313 0.154349
R5082 VSS.n9223 VSS.n9218 0.154349
R5083 VSS.n7822 VSS.n7809 0.154349
R5084 VSS.n7862 VSS.n7857 0.154349
R5085 VSS.n7743 VSS.n7730 0.154349
R5086 VSS.n8976 VSS.n8971 0.154349
R5087 VSS.n7686 VSS.n7685 0.154349
R5088 VSS.n7766 VSS.n7761 0.154349
R5089 VSS.n7082 VSS.n7076 0.154349
R5090 VSS.n7106 VSS.n7101 0.154349
R5091 VSS.n8907 VSS.n8902 0.154349
R5092 VSS.n6618 VSS.n6617 0.154349
R5093 VSS.n6648 VSS.n6645 0.154349
R5094 VSS.n6600 VSS.n6597 0.154349
R5095 VSS.n6524 VSS.n6511 0.154349
R5096 VSS.n6551 VSS.n6546 0.154349
R5097 VSS.n6472 VSS.n6463 0.154349
R5098 VSS.n6502 VSS.n6499 0.154349
R5099 VSS.n6309 VSS.n6303 0.154349
R5100 VSS.n6374 VSS.n6367 0.154349
R5101 VSS.n6771 VSS.n6770 0.154349
R5102 VSS.n6357 VSS.n6351 0.154349
R5103 VSS.n3868 VSS.n3864 0.154349
R5104 VSS.n7303 VSS.n7297 0.154349
R5105 VSS.n4143 VSS.n4138 0.154349
R5106 VSS.n4370 VSS.n4365 0.154349
R5107 VSS.n4338 VSS.n4333 0.154349
R5108 VSS.n4314 VSS.n4313 0.154349
R5109 VSS.n4214 VSS.n4209 0.154349
R5110 VSS.n4424 VSS.n4423 0.154349
R5111 VSS.n874 VSS.n868 0.154349
R5112 VSS.n2409 VSS.n2408 0.154349
R5113 VSS.n14184 VSS.n14183 0.154349
R5114 VSS.n923 VSS.n922 0.154349
R5115 VSS.n12403 VSS.n12402 0.154349
R5116 VSS.n2539 VSS.n2532 0.154349
R5117 VSS.n13078 VSS.n13077 0.154349
R5118 VSS.n2382 VSS.n2377 0.154349
R5119 VSS.n1923 VSS.n1917 0.154349
R5120 VSS.n2284 VSS.n2283 0.154349
R5121 VSS.n14162 VSS.n14155 0.154349
R5122 VSS.n901 VSS.n898 0.154349
R5123 VSS.n1678 VSS.n1673 0.154349
R5124 VSS.n644 VSS.n643 0.154349
R5125 VSS.n13685 VSS.n13676 0.154349
R5126 VSS.n14070 VSS.n14065 0.154349
R5127 VSS.n13216 VSS.n13210 0.154349
R5128 VSS.n13538 VSS.n13531 0.154349
R5129 VSS.n852 VSS.n847 0.154349
R5130 VSS.n2195 VSS.n2189 0.154349
R5131 VSS.n1999 VSS.n1998 0.154349
R5132 VSS.n2114 VSS.n2113 0.154349
R5133 VSS.n2074 VSS.n2073 0.154349
R5134 VSS.n12658 VSS.n12646 0.154349
R5135 VSS.n1872 VSS.n1869 0.154349
R5136 VSS.n12675 VSS.n12674 0.154349
R5137 VSS.n1803 VSS.n1798 0.154349
R5138 VSS.n2307 VSS.n2302 0.154349
R5139 VSS.n2705 VSS.n2704 0.154349
R5140 VSS.n2578 VSS.n2577 0.154349
R5141 VSS.n12940 VSS.n12935 0.154349
R5142 VSS.n2759 VSS.n2758 0.154349
R5143 VSS.n12626 VSS.n12617 0.154349
R5144 VSS.n12863 VSS.n12858 0.154349
R5145 VSS.n3066 VSS.n3065 0.154349
R5146 VSS.n3008 VSS.n3003 0.154349
R5147 VSS.n13012 VSS.n13007 0.154349
R5148 VSS.n2988 VSS.n2987 0.154349
R5149 VSS.n13979 VSS.n13978 0.154349
R5150 VSS.n13521 VSS.n13515 0.154349
R5151 VSS.n13493 VSS.n13480 0.154346
R5152 VSS.n13571 VSS.n13570 0.154346
R5153 VSS.n13598 VSS.n13597 0.154346
R5154 VSS.n1728 VSS.n1715 0.154346
R5155 VSS.n13954 VSS.n13953 0.154346
R5156 VSS.n14011 VSS.n14010 0.154346
R5157 VSS.n12771 VSS.n12770 0.154346
R5158 VSS.n12749 VSS.n12736 0.154346
R5159 VSS.n12791 VSS.n2929 0.154346
R5160 VSS.n2621 VSS.n2620 0.154346
R5161 VSS.n3040 VSS.n3035 0.154346
R5162 VSS.n12891 VSS.n12890 0.154346
R5163 VSS.n2884 VSS.n2879 0.154346
R5164 VSS.n2779 VSS.n2769 0.154346
R5165 VSS.n2803 VSS.n2802 0.154346
R5166 VSS.n2266 VSS.n2265 0.154346
R5167 VSS.n1840 VSS.n1830 0.154346
R5168 VSS.n2163 VSS.n2162 0.154346
R5169 VSS.n1424 VSS.n1423 0.154346
R5170 VSS.n13656 VSS.n13651 0.154346
R5171 VSS.n10866 VSS.n10865 0.154346
R5172 VSS.n7350 VSS.n7280 0.154346
R5173 VSS.n10886 VSS.n3892 0.154346
R5174 VSS.n10904 VSS.n10899 0.154346
R5175 VSS.n10977 VSS.n10976 0.154346
R5176 VSS.n10931 VSS.n10928 0.154346
R5177 VSS.n11017 VSS.n11016 0.154346
R5178 VSS.n6404 VSS.n6334 0.154346
R5179 VSS.n11037 VSS.n3824 0.154346
R5180 VSS.n6666 VSS.n6656 0.154346
R5181 VSS.n6280 VSS.n6270 0.154346
R5182 VSS.n7013 VSS.n7001 0.154346
R5183 VSS.n6966 VSS.n6965 0.154346
R5184 VSS.n6570 VSS.n6560 0.154346
R5185 VSS.n7883 VSS.n7871 0.154346
R5186 VSS.n7715 VSS.n7714 0.154346
R5187 VSS.n7794 VSS.n7793 0.154346
R5188 VSS.n9254 VSS.n9253 0.154346
R5189 VSS.n9821 VSS.n9820 0.154346
R5190 VSS.n9572 VSS.n9571 0.154346
R5191 VSS.n7986 VSS.n7976 0.154346
R5192 VSS.n8172 VSS.n8161 0.154346
R5193 VSS.n8495 VSS.n8491 0.154346
R5194 VSS.n8371 VSS.n8365 0.154346
R5195 VSS.n8204 VSS.n8193 0.154346
R5196 VSS.n8394 VSS.n8390 0.154346
R5197 VSS.n8267 VSS.n8261 0.154346
R5198 VSS.n8260 VSS.n8246 0.154346
R5199 VSS.n8229 VSS.n8223 0.154346
R5200 VSS.n8855 VSS.n8850 0.154346
R5201 VSS.n6724 VSS.n6719 0.154346
R5202 VSS.n9963 VSS.n9962 0.154346
R5203 VSS.n6225 VSS.n6212 0.154346
R5204 VSS.n6758 VSS.n6717 0.154346
R5205 VSS.n6705 VSS.n6691 0.154346
R5206 VSS.n8133 VSS.n8132 0.154346
R5207 VSS.n8027 VSS.n8015 0.154346
R5208 VSS.n8111 VSS.n8097 0.154346
R5209 VSS.n8086 VSS.n8076 0.154346
R5210 VSS.n8055 VSS.n8050 0.154346
R5211 VSS.n8890 VSS.n7974 0.154346
R5212 VSS.n7962 VSS.n7947 0.154346
R5213 VSS.n8809 VSS.n8796 0.154346
R5214 VSS.n7587 VSS.n7574 0.154346
R5215 VSS.n9585 VSS.n7550 0.154346
R5216 VSS.n9198 VSS.n9197 0.154346
R5217 VSS.n9305 VSS.n9304 0.154346
R5218 VSS.n9280 VSS.n9279 0.154346
R5219 VSS.n9010 VSS.n8993 0.154346
R5220 VSS.n9498 VSS.n9497 0.154346
R5221 VSS.n9485 VSS.n9469 0.154346
R5222 VSS.n7239 VSS.n7217 0.154346
R5223 VSS.n7174 VSS.n7157 0.154346
R5224 VSS.n7202 VSS.n7189 0.154346
R5225 VSS.n7252 VSS.n7251 0.154346
R5226 VSS.n7362 VSS.n7352 0.154346
R5227 VSS.n7328 VSS.n7313 0.154346
R5228 VSS.n9174 VSS.n9159 0.154346
R5229 VSS.n9231 VSS.n9218 0.154346
R5230 VSS.n7838 VSS.n7837 0.154346
R5231 VSS.n7917 VSS.n7895 0.154346
R5232 VSS.n8962 VSS.n7809 0.154346
R5233 VSS.n7870 VSS.n7857 0.154346
R5234 VSS.n8990 VSS.n7611 0.154346
R5235 VSS.n7752 VSS.n7730 0.154346
R5236 VSS.n8977 VSS.n8976 0.154346
R5237 VSS.n7780 VSS.n7646 0.154346
R5238 VSS.n7686 VSS.n7681 0.154346
R5239 VSS.n7767 VSS.n7766 0.154346
R5240 VSS.n9878 VSS.n9877 0.154346
R5241 VSS.n7082 VSS.n7069 0.154346
R5242 VSS.n7128 VSS.n7127 0.154346
R5243 VSS.n7107 VSS.n7106 0.154346
R5244 VSS.n7928 VSS.n7927 0.154346
R5245 VSS.n8915 VSS.n8902 0.154346
R5246 VSS.n6893 VSS.n6892 0.154346
R5247 VSS.n6618 VSS.n6608 0.154346
R5248 VSS.n6811 VSS.n6795 0.154346
R5249 VSS.n6655 VSS.n6645 0.154346
R5250 VSS.n6879 VSS.n6863 0.154346
R5251 VSS.n6607 VSS.n6597 0.154346
R5252 VSS.n6952 VSS.n6930 0.154346
R5253 VSS.n7044 VSS.n6511 0.154346
R5254 VSS.n6559 VSS.n6546 0.154346
R5255 VSS.n7032 VSS.n7016 0.154346
R5256 VSS.n6473 VSS.n6472 0.154346
R5257 VSS.n6509 VSS.n6499 0.154346
R5258 VSS.n6440 VSS.n6439 0.154346
R5259 VSS.n6309 VSS.n6296 0.154346
R5260 VSS.n6416 VSS.n6406 0.154346
R5261 VSS.n6382 VSS.n6367 0.154346
R5262 VSS.n6826 VSS.n6825 0.154346
R5263 VSS.n6780 VSS.n6770 0.154346
R5264 VSS.n6365 VSS.n6351 0.154346
R5265 VSS.n3868 VSS.n3852 0.154346
R5266 VSS.n7311 VSS.n7297 0.154346
R5267 VSS.n10760 VSS.n10759 0.154346
R5268 VSS.n10781 VSS.n4108 0.154346
R5269 VSS.n4178 VSS.n4161 0.154346
R5270 VSS.n4242 VSS.n4229 0.154346
R5271 VSS.n4151 VSS.n4138 0.154346
R5272 VSS.n4392 VSS.n4391 0.154346
R5273 VSS.n4371 VSS.n4370 0.154346
R5274 VSS.n4289 VSS.n4288 0.154346
R5275 VSS.n4339 VSS.n4338 0.154346
R5276 VSS.n4314 VSS.n4261 0.154346
R5277 VSS.n4224 VSS.n4209 0.154346
R5278 VSS.n4424 VSS.n4414 0.154346
R5279 VSS.n874 VSS.n861 0.154346
R5280 VSS.n941 VSS.n937 0.154346
R5281 VSS.n1961 VSS.n1947 0.154346
R5282 VSS.n2409 VSS.n2397 0.154346
R5283 VSS.n14183 VSS.n14182 0.154346
R5284 VSS.n564 VSS.n544 0.154346
R5285 VSS.n14216 VSS.n14215 0.154346
R5286 VSS.n595 VSS.n583 0.154346
R5287 VSS.n1148 VSS.n935 0.154346
R5288 VSS.n923 VSS.n909 0.154346
R5289 VSS.n13119 VSS.n13118 0.154346
R5290 VSS.n2513 VSS.n2499 0.154346
R5291 VSS.n2472 VSS.n2460 0.154346
R5292 VSS.n12402 VSS.n12397 0.154346
R5293 VSS.n13040 VSS.n13030 0.154346
R5294 VSS.n2547 VSS.n2532 0.154346
R5295 VSS.n13077 VSS.n13076 0.154346
R5296 VSS.n2445 VSS.n2430 0.154346
R5297 VSS.n13105 VSS.n2351 0.154346
R5298 VSS.n2383 VSS.n2382 0.154346
R5299 VSS.n1923 VSS.n1910 0.154346
R5300 VSS.n2339 VSS.n1945 0.154346
R5301 VSS.n2284 VSS.n2280 0.154346
R5302 VSS.n14172 VSS.n14155 0.154346
R5303 VSS.n908 VSS.n898 0.154346
R5304 VSS.n1380 VSS.n1379 0.154346
R5305 VSS.n1178 VSS.n1172 0.154346
R5306 VSS.n1695 VSS.n1673 0.154346
R5307 VSS.n1450 VSS.n1449 0.154346
R5308 VSS.n644 VSS.n627 0.154346
R5309 VSS.n14097 VSS.n14096 0.154346
R5310 VSS.n14084 VSS.n1641 0.154346
R5311 VSS.n13686 VSS.n13685 0.154346
R5312 VSS.n14071 VSS.n14070 0.154346
R5313 VSS.n13889 VSS.n13888 0.154346
R5314 VSS.n13216 VSS.n13203 0.154346
R5315 VSS.n13638 VSS.n13628 0.154346
R5316 VSS.n13546 VSS.n13531 0.154346
R5317 VSS.n827 VSS.n812 0.154346
R5318 VSS.n860 VSS.n847 0.154346
R5319 VSS.n2228 VSS.n2227 0.154346
R5320 VSS.n2044 VSS.n2043 0.154346
R5321 VSS.n2204 VSS.n2189 0.154346
R5322 VSS.n1999 VSS.n1982 0.154346
R5323 VSS.n2093 VSS.n2092 0.154346
R5324 VSS.n2114 VSS.n2109 0.154346
R5325 VSS.n2074 VSS.n2057 0.154346
R5326 VSS.n2149 VSS.n2133 0.154346
R5327 VSS.n12667 VSS.n12646 0.154346
R5328 VSS.n1879 VSS.n1869 0.154346
R5329 VSS.n13916 VSS.n1829 0.154346
R5330 VSS.n12674 VSS.n12669 0.154346
R5331 VSS.n13939 VSS.n1772 0.154346
R5332 VSS.n1804 VSS.n1803 0.154346
R5333 VSS.n2015 VSS.n2010 0.154346
R5334 VSS.n2308 VSS.n2307 0.154346
R5335 VSS.n12968 VSS.n12967 0.154346
R5336 VSS.n2704 VSS.n2699 0.154346
R5337 VSS.n2651 VSS.n2650 0.154346
R5338 VSS.n2578 VSS.n2561 0.154346
R5339 VSS.n12954 VSS.n2668 0.154346
R5340 VSS.n12941 VSS.n12940 0.154346
R5341 VSS.n2832 VSS.n2831 0.154346
R5342 VSS.n2759 VSS.n2742 0.154346
R5343 VSS.n12877 VSS.n2848 0.154346
R5344 VSS.n12627 VSS.n12626 0.154346
R5345 VSS.n12864 VSS.n12863 0.154346
R5346 VSS.n12711 VSS.n3034 0.154346
R5347 VSS.n3065 VSS.n3060 0.154346
R5348 VSS.n12734 VSS.n2950 0.154346
R5349 VSS.n3009 VSS.n3008 0.154346
R5350 VSS.n2595 VSS.n2589 0.154346
R5351 VSS.n13013 VSS.n13012 0.154346
R5352 VSS.n2988 VSS.n2975 0.154346
R5353 VSS.n13979 VSS.n1758 0.154346
R5354 VSS.n13529 VSS.n13515 0.154346
R5355 VSS.n5786 VSS 0.1505
R5356 VSS.n13493 VSS.n13492 0.149542
R5357 VSS.n13570 VSS.n13562 0.149542
R5358 VSS.n1728 VSS.n1727 0.149542
R5359 VSS.n13953 VSS.n13946 0.149542
R5360 VSS.n12770 VSS.n12765 0.149542
R5361 VSS.n12740 VSS.n12736 0.149542
R5362 VSS.n3041 VSS.n3040 0.149542
R5363 VSS.n12890 VSS.n12883 0.149542
R5364 VSS.n2779 VSS.n2778 0.149542
R5365 VSS.n1840 VSS.n1839 0.149542
R5366 VSS.n2162 VSS.n2155 0.149542
R5367 VSS.n13657 VSS.n13656 0.149542
R5368 VSS.n10865 VSS.n10860 0.149542
R5369 VSS.n7284 VSS.n7280 0.149542
R5370 VSS.n10905 VSS.n10904 0.149542
R5371 VSS.n10976 VSS.n10971 0.149542
R5372 VSS.n11016 VSS.n11011 0.149542
R5373 VSS.n6338 VSS.n6334 0.149542
R5374 VSS.n6280 VSS.n6279 0.149542
R5375 VSS.n7002 VSS.n7001 0.149542
R5376 VSS.n6965 VSS.n6958 0.149542
R5377 VSS.n7714 VSS.n7707 0.149542
R5378 VSS.n7793 VSS.n7786 0.149542
R5379 VSS.n9820 VSS.n9813 0.149542
R5380 VSS.n7986 VSS.n7985 0.149542
R5381 VSS.n8495 VSS.n8494 0.149542
R5382 VSS.n8372 VSS.n8371 0.149542
R5383 VSS.n8394 VSS.n8393 0.149542
R5384 VSS.n8268 VSS.n8267 0.149542
R5385 VSS.n8250 VSS.n8246 0.149542
R5386 VSS.n8855 VSS.n8854 0.149542
R5387 VSS.n6724 VSS.n6723 0.149542
R5388 VSS.n9962 VSS.n9955 0.149542
R5389 VSS.n6759 VSS.n6758 0.149542
R5390 VSS.n8027 VSS.n8026 0.149542
R5391 VSS.n8112 VSS.n8111 0.149542
R5392 VSS.n8891 VSS.n8890 0.149542
R5393 VSS.n9585 VSS.n9584 0.149542
R5394 VSS.n9198 VSS.n9196 0.149542
R5395 VSS.n9279 VSS.n9273 0.149542
R5396 VSS.n9498 VSS.n9496 0.149542
R5397 VSS.n9470 VSS.n9469 0.149542
R5398 VSS.n7202 VSS.n7201 0.149542
R5399 VSS.n7353 VSS.n7352 0.149542
R5400 VSS.n9174 VSS.n9173 0.149542
R5401 VSS.n7837 VSS.n7832 0.149542
R5402 VSS.n7898 VSS.n7895 0.149542
R5403 VSS.n7625 VSS.n7611 0.149542
R5404 VSS.n7660 VSS.n7646 0.149542
R5405 VSS.n9877 VSS.n9870 0.149542
R5406 VSS.n7127 VSS.n7122 0.149542
R5407 VSS.n7927 VSS.n7922 0.149542
R5408 VSS.n6892 VSS.n6885 0.149542
R5409 VSS.n6796 VSS.n6795 0.149542
R5410 VSS.n6864 VSS.n6863 0.149542
R5411 VSS.n6933 VSS.n6930 0.149542
R5412 VSS.n7017 VSS.n7016 0.149542
R5413 VSS.n6439 VSS.n6432 0.149542
R5414 VSS.n6407 VSS.n6406 0.149542
R5415 VSS.n6825 VSS.n6818 0.149542
R5416 VSS.n10759 VSS.n10752 0.149542
R5417 VSS.n4122 VSS.n4108 0.149542
R5418 VSS.n4179 VSS.n4178 0.149542
R5419 VSS.n4242 VSS.n4241 0.149542
R5420 VSS.n4391 VSS.n4386 0.149542
R5421 VSS.n4288 VSS.n4281 0.149542
R5422 VSS.n941 VSS.n940 0.149542
R5423 VSS.n1961 VSS.n1960 0.149542
R5424 VSS.n564 VSS.n563 0.149542
R5425 VSS.n14215 VSS.n14210 0.149542
R5426 VSS.n595 VSS.n594 0.149542
R5427 VSS.n1149 VSS.n1148 0.149542
R5428 VSS.n13118 VSS.n13111 0.149542
R5429 VSS.n2513 VSS.n2512 0.149542
R5430 VSS.n2472 VSS.n2471 0.149542
R5431 VSS.n13031 VSS.n13030 0.149542
R5432 VSS.n2433 VSS.n2430 0.149542
R5433 VSS.n2366 VSS.n2351 0.149542
R5434 VSS.n2340 VSS.n2339 0.149542
R5435 VSS.n1380 VSS.n1378 0.149542
R5436 VSS.n1179 VSS.n1178 0.149542
R5437 VSS.n1449 VSS.n1443 0.149542
R5438 VSS.n14097 VSS.n14095 0.149542
R5439 VSS.n1655 VSS.n1641 0.149542
R5440 VSS.n13888 VSS.n13881 0.149542
R5441 VSS.n13629 VSS.n13628 0.149542
R5442 VSS.n827 VSS.n826 0.149542
R5443 VSS.n2227 VSS.n2220 0.149542
R5444 VSS.n2043 VSS.n2037 0.149542
R5445 VSS.n2092 VSS.n2086 0.149542
R5446 VSS.n2134 VSS.n2133 0.149542
R5447 VSS.n1829 VSS.n1821 0.149542
R5448 VSS.n1787 VSS.n1772 0.149542
R5449 VSS.n2016 VSS.n2015 0.149542
R5450 VSS.n12967 VSS.n12960 0.149542
R5451 VSS.n2650 VSS.n2644 0.149542
R5452 VSS.n2682 VSS.n2668 0.149542
R5453 VSS.n2831 VSS.n2825 0.149542
R5454 VSS.n2862 VSS.n2848 0.149542
R5455 VSS.n3034 VSS.n3026 0.149542
R5456 VSS.n2965 VSS.n2950 0.149542
R5457 VSS.n2596 VSS.n2595 0.149542
R5458 VSS.n6150 VSS 0.147559
R5459 VSS.n5967 VSS 0.147559
R5460 VSS.n8510 VSS 0.146833
R5461 VSS.n6209 VSS 0.146833
R5462 VSS VSS.n9950 0.146833
R5463 VSS.n8158 VSS 0.146833
R5464 VSS VSS.n8433 0.146833
R5465 VSS.n11114 VSS 0.146833
R5466 VSS VSS.n11007 0.146833
R5467 VSS.n10955 VSS 0.146833
R5468 VSS VSS.n10856 0.146833
R5469 VSS.n4089 VSS 0.146833
R5470 VSS.n10783 VSS 0.146833
R5471 VSS VSS.n4153 0.146833
R5472 VSS VSS.n4276 0.146833
R5473 VSS.n4351 VSS 0.146833
R5474 VSS.n4412 VSS 0.146833
R5475 VSS VSS.n10747 0.146833
R5476 VSS.n14236 VSS 0.146833
R5477 VSS.n10710 VSS 0.146833
R5478 VSS VSS.n12431 0.146833
R5479 VSS.n13060 VSS 0.146833
R5480 VSS VSS.n2429 0.146833
R5481 VSS.n12825 VSS 0.146833
R5482 VSS VSS.n1747 0.146833
R5483 VSS.n14024 VSS 0.146833
R5484 VSS.n13610 VSS 0.146833
R5485 VSS VSS.n13429 0.146833
R5486 VSS.n5916 VSS.n4677 0.142792
R5487 VSS.n6098 VSS.n4668 0.142557
R5488 VSS.n10525 VSS.n20 0.140359
R5489 VSS.n10538 VSS.n21 0.140359
R5490 VSS.n10172 VSS.n10171 0.140147
R5491 VSS.n10170 VSS.n4561 0.140147
R5492 VSS.n4563 VSS.n4562 0.140147
R5493 VSS.n5178 VSS.n5177 0.140147
R5494 VSS.n5175 VSS.n4718 0.140147
R5495 VSS.n5158 VSS.n5157 0.140147
R5496 VSS.n5153 VSS.n4731 0.140147
R5497 VSS.n5148 VSS.n5147 0.140147
R5498 VSS.n5146 VSS.n4734 0.140147
R5499 VSS.n5141 VSS.n5140 0.140147
R5500 VSS.n5139 VSS.n4737 0.140147
R5501 VSS.n5134 VSS.n4738 0.140147
R5502 VSS.n5118 VSS.n5116 0.140147
R5503 VSS.n5114 VSS.n5113 0.140147
R5504 VSS.n5111 VSS.n4745 0.140147
R5505 VSS.n3594 VSS.n3593 0.140147
R5506 VSS.n12304 VSS.n12298 0.140147
R5507 VSS.n12480 VSS.n3604 0.140147
R5508 VSS.n12517 VSS.n12516 0.140147
R5509 VSS.n12515 VSS.n3592 0.140147
R5510 VSS.n10541 VSS.n10540 0.140147
R5511 VSS.n12551 VSS.n3320 0.140147
R5512 VSS.n12530 VSS.n12529 0.140147
R5513 VSS.n12528 VSS.n3380 0.140147
R5514 VSS.n12526 VSS.n3586 0.140147
R5515 VSS.n12524 VSS.n3588 0.140147
R5516 VSS.n12522 VSS.n3589 0.140147
R5517 VSS.n8511 VSS.n8510 0.14005
R5518 VSS.n9950 VSS.n9949 0.14005
R5519 VSS.n6210 VSS.n6209 0.14005
R5520 VSS.n8159 VSS.n8158 0.14005
R5521 VSS.n4276 VSS.n4275 0.14005
R5522 VSS.n4412 VSS.n4160 0.14005
R5523 VSS.n14237 VSS.n14236 0.14005
R5524 VSS.n13061 VSS.n13060 0.14005
R5525 VSS.n12431 VSS.n12430 0.14005
R5526 VSS.n2429 VSS.n2428 0.14005
R5527 VSS.n10631 VSS.n4545 0.139843
R5528 VSS.n12303 VSS.n3605 0.139843
R5529 VSS.n10630 VSS.n10629 0.139843
R5530 VSS.n9985 VSS.n9984 0.13959
R5531 VSS.n8124 VSS.n8123 0.13959
R5532 VSS.n8834 VSS.n8833 0.13959
R5533 VSS.n4435 VSS.n4434 0.13959
R5534 VSS.n4359 VSS.n4358 0.13959
R5535 VSS.n12422 VSS.n12421 0.13959
R5536 VSS.n13068 VSS.n13067 0.13959
R5537 VSS.n2422 VSS.n2421 0.13959
R5538 VSS.n4534 VSS 0.137248
R5539 VSS.n1515 VSS.n1513 0.136775
R5540 VSS.n8429 VSS.n8428 0.136775
R5541 VSS.n8625 VSS.n8624 0.136775
R5542 VSS.n8712 VSS.n8711 0.136775
R5543 VSS.n9700 VSS.n9699 0.136775
R5544 VSS.n9116 VSS.n9057 0.136775
R5545 VSS.n7483 VSS.n7482 0.136775
R5546 VSS.n4029 VSS.n4028 0.136775
R5547 VSS.n9770 VSS.n9768 0.136775
R5548 VSS.n9424 VSS.n9422 0.136775
R5549 VSS.n10716 VSS.n10715 0.136775
R5550 VSS.n994 VSS.n992 0.136775
R5551 VSS.n14360 VSS.n14358 0.136775
R5552 VSS.n14371 VSS.n14370 0.136775
R5553 VSS.n1074 VSS.n1072 0.136775
R5554 VSS.n1245 VSS.n1243 0.136775
R5555 VSS.n1324 VSS.n1322 0.136775
R5556 VSS.n464 VSS.n463 0.136775
R5557 VSS.n13756 VSS.n13754 0.136775
R5558 VSS.n13293 VSS.n13292 0.136775
R5559 VSS.n13371 VSS.n13369 0.136775
R5560 VSS.n13836 VSS.n13834 0.136775
R5561 VSS.n1596 VSS.n1594 0.136775
R5562 VSS.n13426 VSS.n13424 0.136775
R5563 VSS.n11276 VSS 0.129576
R5564 VSS.n5375 VSS.n4709 0.128457
R5565 VSS.n8639 VSS.n8638 0.127988
R5566 VSS.n8723 VSS.n8722 0.127988
R5567 VSS.n9714 VSS.n9713 0.127988
R5568 VSS.n5555 VSS.n4697 0.127988
R5569 VSS.n5195 VSS.n5183 0.126108
R5570 VSS.n9747 VSS.n9746 0.125637
R5571 VSS.n13427 VSS 0.1255
R5572 VSS.n13401 VSS 0.1255
R5573 VSS.n1713 VSS 0.1255
R5574 VSS.n1746 VSS 0.1255
R5575 VSS.n2928 VSS 0.1255
R5576 VSS.n1516 VSS 0.1255
R5577 VSS.n3909 VSS 0.1255
R5578 VSS.n3891 VSS 0.1255
R5579 VSS.n3842 VSS 0.1255
R5580 VSS.n3823 VSS 0.1255
R5581 VSS.n9359 VSS 0.1255
R5582 VSS.n8489 VSS 0.1255
R5583 VSS.n4660 VSS 0.1255
R5584 VSS.n8121 VSS 0.1255
R5585 VSS.n8014 VSS 0.1255
R5586 VSS.n8342 VSS 0.1255
R5587 VSS.n8728 VSS 0.1255
R5588 VSS.n7519 VSS 0.1255
R5589 VSS.n7497 VSS 0.1255
R5590 VSS.n7419 VSS 0.1255
R5591 VSS.n10817 VSS 0.1255
R5592 VSS.n4670 VSS 0.1255
R5593 VSS.n4679 VSS 0.1255
R5594 VSS.n4688 VSS 0.1255
R5595 VSS.n4699 VSS 0.1255
R5596 VSS.n4711 VSS 0.1255
R5597 VSS.n5185 VSS 0.1255
R5598 VSS.n10132 VSS 0.1255
R5599 VSS.n11080 VSS 0.1255
R5600 VSS.n10745 VSS 0.1255
R5601 VSS.n4152 VSS 0.1255
R5602 VSS.n4203 VSS 0.1255
R5603 VSS.n4330 VSS 0.1255
R5604 VSS.n4329 VSS.n4260 0.1255
R5605 VSS.n4227 VSS 0.1255
R5606 VSS.n4159 VSS 0.1255
R5607 VSS.n543 VSS 0.1255
R5608 VSS.n12396 VSS 0.1255
R5609 VSS.n2458 VSS 0.1255
R5610 VSS.n2396 VSS 0.1255
R5611 VSS.n14368 VSS 0.1255
R5612 VSS.n995 VSS 0.1255
R5613 VSS.n1246 VSS 0.1255
R5614 VSS.n707 VSS 0.1255
R5615 VSS.n13757 VSS 0.1255
R5616 VSS.n13294 VSS 0.1255
R5617 VSS.n12344 VSS 0.1255
R5618 VSS.n11691 VSS 0.1255
R5619 VSS.n11777 VSS 0.1255
R5620 VSS.n11824 VSS 0.1255
R5621 VSS.n3395 VSS 0.1255
R5622 VSS.n3355 VSS 0.1255
R5623 VSS.n3186 VSS 0.1255
R5624 VSS.n12813 VSS 0.1255
R5625 VSS.n5735 VSS.n4686 0.12505
R5626 VSS.n14480 VSS.t0 0.124605
R5627 VSS.n4525 VSS 0.1227
R5628 VSS.n10812 VSS.n10811 0.122113
R5629 VSS.n10143 VSS.n10130 0.122113
R5630 VSS.n9731 VSS.n9730 0.121642
R5631 VSS.n11412 VSS.n11411 0.120292
R5632 VSS.n11411 VSS.n11410 0.120292
R5633 VSS.n11410 VSS.n11408 0.120292
R5634 VSS.n11408 VSS.n11406 0.120292
R5635 VSS.n11406 VSS.n11404 0.120292
R5636 VSS.n11404 VSS.n11402 0.120292
R5637 VSS.n11402 VSS.n11400 0.120292
R5638 VSS.n11400 VSS.n11398 0.120292
R5639 VSS.n11398 VSS.n11396 0.120292
R5640 VSS.n11393 VSS.n11392 0.120292
R5641 VSS.n11392 VSS.n11391 0.120292
R5642 VSS.n11391 VSS.n11390 0.120292
R5643 VSS.n11390 VSS.n11388 0.120292
R5644 VSS.n11388 VSS.n11386 0.120292
R5645 VSS.n11386 VSS.n11384 0.120292
R5646 VSS.n11384 VSS.n11382 0.120292
R5647 VSS.n11382 VSS.n11380 0.120292
R5648 VSS.n11380 VSS.n11378 0.120292
R5649 VSS.n11375 VSS.n11374 0.120292
R5650 VSS.n11374 VSS.n11373 0.120292
R5651 VSS.n11373 VSS.n11372 0.120292
R5652 VSS.n11372 VSS.n11370 0.120292
R5653 VSS.n11370 VSS.n11368 0.120292
R5654 VSS.n11368 VSS.n11366 0.120292
R5655 VSS.n11366 VSS.n11364 0.120292
R5656 VSS.n11364 VSS.n11362 0.120292
R5657 VSS.n11362 VSS.n11360 0.120292
R5658 VSS.n11356 VSS.n11355 0.120292
R5659 VSS.n11353 VSS.n11351 0.120292
R5660 VSS.n3674 VSS.n3673 0.120292
R5661 VSS.n3669 VSS.n3668 0.120292
R5662 VSS.n3664 VSS.n3663 0.120292
R5663 VSS.n3663 VSS.n3643 0.120292
R5664 VSS.n3659 VSS.n3643 0.120292
R5665 VSS.n3659 VSS.n3658 0.120292
R5666 VSS.n3654 VSS.n3653 0.120292
R5667 VSS.n3653 VSS.n3651 0.120292
R5668 VSS.n3651 VSS.n3650 0.120292
R5669 VSS.n3650 VSS.n3648 0.120292
R5670 VSS.n11235 VSS.n11234 0.120292
R5671 VSS.n11240 VSS.n11239 0.120292
R5672 VSS.n11245 VSS.n11244 0.120292
R5673 VSS.n11245 VSS.n11217 0.120292
R5674 VSS.n11249 VSS.n11217 0.120292
R5675 VSS.n11250 VSS.n11249 0.120292
R5676 VSS.n11215 VSS.n11214 0.120292
R5677 VSS.n11256 VSS.n11214 0.120292
R5678 VSS.n11257 VSS.n11256 0.120292
R5679 VSS.n11258 VSS.n11257 0.120292
R5680 VSS.n9758 VSS.n9757 0.119998
R5681 VSS.n11332 VSS.n11331 0.119058
R5682 VSS.n11334 VSS.n3622 0.119058
R5683 VSS.n11186 VSS.n11185 0.118209
R5684 VSS.n4535 VSS.n4534 0.112194
R5685 VSS.n4525 VSS.n4100 0.112194
R5686 VSS.n13609 VSS.n13480 0.106269
R5687 VSS.n13571 VSS.n13240 0.106269
R5688 VSS.n13598 VSS.n13591 0.106269
R5689 VSS.n14022 VSS.n1715 0.106269
R5690 VSS.n13954 VSS.n13942 0.106269
R5691 VSS.n14011 VSS.n14004 0.106269
R5692 VSS.n12771 VSS.n12762 0.106269
R5693 VSS.n12750 VSS.n12749 0.106269
R5694 VSS.n12802 VSS.n2929 0.106269
R5695 VSS.n2621 VSS.n2560 0.106269
R5696 VSS.n12644 VSS.n3035 0.106269
R5697 VSS.n12891 VSS.n12879 0.106269
R5698 VSS.n2903 VSS.n2879 0.106269
R5699 VSS.n2821 VSS.n2769 0.106269
R5700 VSS.n2803 VSS.n2741 0.106269
R5701 VSS.n2266 VSS.n2254 0.106269
R5702 VSS.n13201 VSS.n1830 0.106269
R5703 VSS.n2163 VSS.n2151 0.106269
R5704 VSS.n1424 VSS.n626 0.106269
R5705 VSS.n13703 VSS.n13651 0.106269
R5706 VSS.n10866 VSS.n10857 0.106269
R5707 VSS.n7351 VSS.n7350 0.106269
R5708 VSS.n10897 VSS.n3892 0.106269
R5709 VSS.n10953 VSS.n10899 0.106269
R5710 VSS.n10977 VSS.n10967 0.106269
R5711 VSS.n10928 VSS.n10921 0.106269
R5712 VSS.n11017 VSS.n11008 0.106269
R5713 VSS.n6405 VSS.n6404 0.106269
R5714 VSS.n11048 VSS.n3824 0.106269
R5715 VSS.n6846 VSS.n6656 0.106269
R5716 VSS.n7066 VSS.n6270 0.106269
R5717 VSS.n7034 VSS.n7013 0.106269
R5718 VSS.n6966 VSS.n6954 0.106269
R5719 VSS.n6986 VSS.n6560 0.106269
R5720 VSS.n8938 VSS.n7871 0.106269
R5721 VSS.n7715 VSS.n7145 0.106269
R5722 VSS.n7794 VSS.n7782 0.106269
R5723 VSS.n9254 VSS.n8992 0.106269
R5724 VSS.n9821 VSS.n9809 0.106269
R5725 VSS.n9571 VSS.n7565 0.106269
R5726 VSS.n7999 VSS.n7976 0.106269
R5727 VSS.n8832 VSS.n8161 0.106269
R5728 VSS.n8509 VSS.n8491 0.106269
R5729 VSS.n8389 VSS.n8365 0.106269
R5730 VSS.n8794 VSS.n8193 0.106269
R5731 VSS.n8408 VSS.n8390 0.106269
R5732 VSS.n8285 VSS.n8261 0.106269
R5733 VSS.n8771 VSS.n8260 0.106269
R5734 VSS.n8223 VSS.n7588 0.106269
R5735 VSS.n8850 VSS.n8849 0.106269
R5736 VSS.n6737 VSS.n6719 0.106269
R5737 VSS.n9963 VSS.n9951 0.106269
R5738 VSS.n9983 VSS.n6212 0.106269
R5739 VSS.n6739 VSS.n6717 0.106269
R5740 VSS.n6767 VSS.n6691 0.106269
R5741 VSS.n8132 VSS.n8125 0.106269
R5742 VSS.n8157 VSS.n8015 0.106269
R5743 VSS.n8097 VSS.n8007 0.106269
R5744 VSS.n8087 VSS.n8086 0.106269
R5745 VSS.n8074 VSS.n8050 0.106269
R5746 VSS.n8000 VSS.n7974 0.106269
R5747 VSS.n8899 VSS.n7947 0.106269
R5748 VSS.n8810 VSS.n8809 0.106269
R5749 VSS.n9548 VSS.n7587 0.106269
R5750 VSS.n9596 VSS.n7550 0.106269
R5751 VSS.n9197 VSS.n7549 0.106269
R5752 VSS.n9305 VSS.n7156 0.106269
R5753 VSS.n9280 VSS.n9271 0.106269
R5754 VSS.n9522 VSS.n8993 0.106269
R5755 VSS.n9497 VSS.n9487 0.106269
R5756 VSS.n9486 VSS.n9485 0.106269
R5757 VSS.n7240 VSS.n7239 0.106269
R5758 VSS.n9844 VSS.n7157 0.106269
R5759 VSS.n7380 VSS.n7189 0.106269
R5760 VSS.n7252 VSS.n7242 0.106269
R5761 VSS.n7363 VSS.n7362 0.106269
R5762 VSS.n7329 VSS.n7328 0.106269
R5763 VSS.n9270 VSS.n9159 0.106269
R5764 VSS.n9234 VSS.n9231 0.106269
R5765 VSS.n7838 VSS.n7609 0.106269
R5766 VSS.n7918 VSS.n7917 0.106269
R5767 VSS.n8963 VSS.n8962 0.106269
R5768 VSS.n8941 VSS.n7870 0.106269
R5769 VSS.n8991 VSS.n8990 0.106269
R5770 VSS.n7753 VSS.n7752 0.106269
R5771 VSS.n8977 VSS.n8966 0.106269
R5772 VSS.n7781 VSS.n7780 0.106269
R5773 VSS.n7681 VSS.n7068 0.106269
R5774 VSS.n7767 VSS.n7756 0.106269
R5775 VSS.n9878 VSS.n9866 0.106269
R5776 VSS.n9898 VSS.n7069 0.106269
R5777 VSS.n7128 VSS.n3881 0.106269
R5778 VSS.n7107 VSS.n3851 0.106269
R5779 VSS.n7928 VSS.n7920 0.106269
R5780 VSS.n8916 VSS.n8915 0.106269
R5781 VSS.n6893 VSS.n6881 0.106269
R5782 VSS.n6913 VSS.n6608 0.106269
R5783 VSS.n6812 VSS.n6811 0.106269
R5784 VSS.n6849 VSS.n6655 0.106269
R5785 VSS.n6880 VSS.n6879 0.106269
R5786 VSS.n6916 VSS.n6607 0.106269
R5787 VSS.n6953 VSS.n6952 0.106269
R5788 VSS.n7045 VSS.n7044 0.106269
R5789 VSS.n6989 VSS.n6559 0.106269
R5790 VSS.n7033 VSS.n7032 0.106269
R5791 VSS.n6473 VSS.n6462 0.106269
R5792 VSS.n7048 VSS.n6509 0.106269
R5793 VSS.n6440 VSS.n6269 0.106269
R5794 VSS.n6460 VSS.n6296 0.106269
R5795 VSS.n6417 VSS.n6416 0.106269
R5796 VSS.n6383 VSS.n6382 0.106269
R5797 VSS.n6826 VSS.n6814 0.106269
R5798 VSS.n6781 VSS.n6780 0.106269
R5799 VSS.n6385 VSS.n6365 0.106269
R5800 VSS.n10993 VSS.n3852 0.106269
R5801 VSS.n7331 VSS.n7311 0.106269
R5802 VSS.n10760 VSS.n10748 0.106269
R5803 VSS.n10782 VSS.n10781 0.106269
R5804 VSS.n4411 VSS.n4161 0.106269
R5805 VSS.n4350 VSS.n4229 0.106269
R5806 VSS.n4443 VSS.n4151 0.106269
R5807 VSS.n4392 VSS.n4384 0.106269
R5808 VSS.n4371 VSS.n4360 0.106269
R5809 VSS.n4289 VSS.n4277 0.106269
R5810 VSS.n4339 VSS.n4332 0.106269
R5811 VSS.n4324 VSS.n4261 0.106269
R5812 VSS.n4225 VSS.n4224 0.106269
R5813 VSS.n4433 VSS.n4414 0.106269
R5814 VSS.n1401 VSS.n861 0.106269
R5815 VSS.n955 VSS.n937 0.106269
R5816 VSS.n2324 VSS.n1947 0.106269
R5817 VSS.n2420 VSS.n2397 0.106269
R5818 VSS.n14182 VSS.n14175 0.106269
R5819 VSS.n14235 VSS.n544 0.106269
R5820 VSS.n14216 VSS.n14208 0.106269
R5821 VSS.n14207 VSS.n583 0.106269
R5822 VSS.n1130 VSS.n935 0.106269
R5823 VSS.n1157 VSS.n909 0.106269
R5824 VSS.n13119 VSS.n13107 0.106269
R5825 VSS.n13029 VSS.n2499 0.106269
R5826 VSS.n13059 VSS.n2460 0.106269
R5827 VSS.n12420 VSS.n12397 0.106269
R5828 VSS.n13041 VSS.n13040 0.106269
R5829 VSS.n2548 VSS.n2547 0.106269
R5830 VSS.n13076 VSS.n13069 0.106269
R5831 VSS.n2446 VSS.n2445 0.106269
R5832 VSS.n13106 VSS.n13105 0.106269
R5833 VSS.n2383 VSS.n1909 0.106269
R5834 VSS.n13139 VSS.n1910 0.106269
R5835 VSS.n2326 VSS.n1945 0.106269
R5836 VSS.n2297 VSS.n2280 0.106269
R5837 VSS.n14173 VSS.n14172 0.106269
R5838 VSS.n1160 VSS.n908 0.106269
R5839 VSS.n1379 VSS.n1369 0.106269
R5840 VSS.n1196 VSS.n1172 0.106269
R5841 VSS.n1696 VSS.n1695 0.106269
R5842 VSS.n1450 VSS.n1441 0.106269
R5843 VSS.n14121 VSS.n627 0.106269
R5844 VSS.n14096 VSS.n14086 0.106269
R5845 VSS.n14085 VSS.n14084 0.106269
R5846 VSS.n13686 VSS.n13202 0.106269
R5847 VSS.n14071 VSS.n14060 0.106269
R5848 VSS.n13889 VSS.n13877 0.106269
R5849 VSS.n13909 VSS.n13203 0.106269
R5850 VSS.n13639 VSS.n13638 0.106269
R5851 VSS.n13547 VSS.n13546 0.106269
R5852 VSS.n1440 VSS.n812 0.106269
R5853 VSS.n1404 VSS.n860 0.106269
R5854 VSS.n2228 VSS.n2216 0.106269
R5855 VSS.n2044 VSS.n2035 0.106269
R5856 VSS.n2205 VSS.n2204 0.106269
R5857 VSS.n2251 VSS.n1982 0.106269
R5858 VSS.n2093 VSS.n2084 0.106269
R5859 VSS.n2109 VSS.n1880 0.106269
R5860 VSS.n2186 VSS.n2057 0.106269
R5861 VSS.n2150 VSS.n2149 0.106269
R5862 VSS.n12668 VSS.n12667 0.106269
R5863 VSS.n13183 VSS.n1879 0.106269
R5864 VSS.n13916 VSS.n13915 0.106269
R5865 VSS.n12693 VSS.n12669 0.106269
R5866 VSS.n13940 VSS.n13939 0.106269
R5867 VSS.n1804 VSS.n1757 0.106269
R5868 VSS.n2034 VSS.n2010 0.106269
R5869 VSS.n2308 VSS.n2300 0.106269
R5870 VSS.n12968 VSS.n12956 0.106269
R5871 VSS.n2723 VSS.n2699 0.106269
R5872 VSS.n2651 VSS.n2642 0.106269
R5873 VSS.n12991 VSS.n2561 0.106269
R5874 VSS.n12955 VSS.n12954 0.106269
R5875 VSS.n12941 VSS.n12930 0.106269
R5876 VSS.n2832 VSS.n2823 0.106269
R5877 VSS.n12914 VSS.n2742 0.106269
R5878 VSS.n12878 VSS.n12877 0.106269
R5879 VSS.n12627 VSS.n12616 0.106269
R5880 VSS.n12864 VSS.n12853 0.106269
R5881 VSS.n12711 VSS.n12710 0.106269
R5882 VSS.n3084 VSS.n3060 0.106269
R5883 VSS.n12735 VSS.n12734 0.106269
R5884 VSS.n3009 VSS.n3000 0.106269
R5885 VSS.n2641 VSS.n2589 0.106269
R5886 VSS.n13013 VSS.n13005 0.106269
R5887 VSS.n2998 VSS.n2975 0.106269
R5888 VSS.n13989 VSS.n1758 0.106269
R5889 VSS.n13550 VSS.n13529 0.106269
R5890 VSS.n8489 VSS.n8488 0.105167
R5891 VSS.n9984 VSS.n4660 0.105167
R5892 VSS.n8124 VSS.n8121 0.105167
R5893 VSS.n8833 VSS.n8014 0.105167
R5894 VSS.n4359 VSS.n4203 0.105167
R5895 VSS.n4434 VSS.n4159 0.105167
R5896 VSS.n10696 VSS.n543 0.105167
R5897 VSS.n12421 VSS.n12396 0.105167
R5898 VSS.n13068 VSS.n2458 0.105167
R5899 VSS.n2421 VSS.n2396 0.105167
R5900 VSS.n13611 VSS.n13479 0.105167
R5901 VSS.n13611 VSS.n13610 0.105167
R5902 VSS.n14025 VSS.n1714 0.105167
R5903 VSS.n1714 VSS.n1713 0.105167
R5904 VSS.n14025 VSS.n14024 0.105167
R5905 VSS.n14003 VSS.n14002 0.105167
R5906 VSS.n14003 VSS.n1746 0.105167
R5907 VSS.n14002 VSS.n1747 0.105167
R5908 VSS.n12826 VSS.n12803 0.105167
R5909 VSS.n12803 VSS.n2928 0.105167
R5910 VSS.n12826 VSS.n12825 0.105167
R5911 VSS.n10855 VSS.n3908 0.105167
R5912 VSS.n10856 VSS.n10855 0.105167
R5913 VSS.n10956 VSS.n10898 0.105167
R5914 VSS.n10898 VSS.n3891 0.105167
R5915 VSS.n10956 VSS.n10955 0.105167
R5916 VSS.n11006 VSS.n3840 0.105167
R5917 VSS.n3842 VSS.n3840 0.105167
R5918 VSS.n11007 VSS.n11006 0.105167
R5919 VSS.n11115 VSS.n11049 0.105167
R5920 VSS.n11049 VSS.n3823 0.105167
R5921 VSS.n11115 VSS.n11114 0.105167
R5922 VSS.n8510 VSS 0.105167
R5923 VSS.n6209 VSS 0.105167
R5924 VSS.n9950 VSS 0.105167
R5925 VSS.n8158 VSS 0.105167
R5926 VSS.n8433 VSS 0.105167
R5927 VSS.n11114 VSS 0.105167
R5928 VSS.n11007 VSS 0.105167
R5929 VSS.n10955 VSS 0.105167
R5930 VSS.n10856 VSS 0.105167
R5931 VSS VSS.n4089 0.105167
R5932 VSS VSS.n10783 0.105167
R5933 VSS.n4352 VSS.n4228 0.105167
R5934 VSS.n4352 VSS.n4351 0.105167
R5935 VSS.n4441 VSS.n4153 0.105167
R5936 VSS.n4442 VSS.n4441 0.105167
R5937 VSS.n4442 VSS.n4152 0.105167
R5938 VSS VSS.n4153 0.105167
R5939 VSS.n4276 VSS 0.105167
R5940 VSS.n4351 VSS 0.105167
R5941 VSS.n4228 VSS.n4227 0.105167
R5942 VSS VSS.n4412 0.105167
R5943 VSS.n10747 VSS 0.105167
R5944 VSS.n14236 VSS 0.105167
R5945 VSS VSS.n10710 0.105167
R5946 VSS.n12431 VSS 0.105167
R5947 VSS.n13060 VSS 0.105167
R5948 VSS.n2429 VSS 0.105167
R5949 VSS.n12825 VSS 0.105167
R5950 VSS VSS.n1747 0.105167
R5951 VSS.n14024 VSS 0.105167
R5952 VSS.n13610 VSS 0.105167
R5953 VSS.n13429 VSS 0.105167
R5954 VSS.n12462 VSS.n12460 0.104667
R5955 VSS.n6153 VSS.n6152 0.104667
R5956 VSS.n8633 VSS.n8342 0.104667
R5957 VSS VSS.n8627 0.104667
R5958 VSS.n8729 VSS.n8728 0.104667
R5959 VSS.n8710 VSS 0.104667
R5960 VSS.n9708 VSS.n7519 0.104667
R5961 VSS VSS.n9702 0.104667
R5962 VSS.n7499 VSS.n7497 0.104667
R5963 VSS.n10818 VSS.n10817 0.104667
R5964 VSS.n4027 VSS 0.104667
R5965 VSS.n9771 VSS 0.104667
R5966 VSS VSS.n9426 0.104667
R5967 VSS.n6089 VSS.n4670 0.104667
R5968 VSS VSS.n5969 0.104667
R5969 VSS.n5907 VSS.n4679 0.104667
R5970 VSS VSS.n5788 0.104667
R5971 VSS.n5726 VSS.n4688 0.104667
R5972 VSS VSS.n5607 0.104667
R5973 VSS.n5546 VSS.n4699 0.104667
R5974 VSS VSS.n5427 0.104667
R5975 VSS.n5366 VSS.n4711 0.104667
R5976 VSS VSS.n5247 0.104667
R5977 VSS.n5186 VSS.n5185 0.104667
R5978 VSS.n10134 VSS.n10132 0.104667
R5979 VSS.n4327 VSS.n4326 0.104667
R5980 VSS VSS.n14362 0.104667
R5981 VSS VSS.n1076 0.104667
R5982 VSS VSS.n1326 0.104667
R5983 VSS.n769 VSS 0.104667
R5984 VSS VSS.n13373 0.104667
R5985 VSS VSS.n13838 0.104667
R5986 VSS VSS.n1598 0.104667
R5987 VSS.n11992 VSS.n11824 0.104667
R5988 VSS VSS.n11931 0.104667
R5989 VSS VSS.n3446 0.104667
R5990 VSS VSS.n12581 0.104667
R5991 VSS.n3291 VSS.n3186 0.104667
R5992 VSS VSS.n3214 0.104667
R5993 VSS.n11778 VSS.n11777 0.104146
R5994 VSS.n12814 VSS.n12812 0.103865
R5995 VSS.n8432 VSS.n8431 0.103365
R5996 VSS.n8632 VSS.n8631 0.103365
R5997 VSS.n8731 VSS.n8730 0.103365
R5998 VSS.n9707 VSS.n9706 0.103365
R5999 VSS.n9118 VSS.n9117 0.103365
R6000 VSS.n9363 VSS.n9362 0.103365
R6001 VSS.n9773 VSS.n9772 0.103365
R6002 VSS.n10820 VSS.n10819 0.103365
R6003 VSS.n6088 VSS.n6087 0.103365
R6004 VSS.n5906 VSS.n5905 0.103365
R6005 VSS.n5725 VSS.n5724 0.103365
R6006 VSS.n5545 VSS.n5544 0.103365
R6007 VSS.n5365 VSS.n5364 0.103365
R6008 VSS.n10098 VSS.n4574 0.103365
R6009 VSS.n10133 VSS.n3716 0.103365
R6010 VSS.n10713 VSS.n10712 0.103365
R6011 VSS.n771 VSS.n710 0.103365
R6012 VSS.n771 VSS.n770 0.103365
R6013 VSS.n12266 VSS.n12265 0.103365
R6014 VSS.n12159 VSS.n12158 0.103365
R6015 VSS.n11991 VSS.n11990 0.103365
R6016 VSS.n3563 VSS.n3562 0.103365
R6017 VSS.n12584 VSS.n3116 0.103365
R6018 VSS.n3290 VSS.n3289 0.103365
R6019 VSS.n3199 VSS 0.103162
R6020 VSS.n3346 VSS 0.103162
R6021 VSS.n11791 VSS 0.103162
R6022 VSS.n11540 VSS 0.103162
R6023 VSS.n3621 VSS 0.103162
R6024 VSS.n11909 VSS 0.103002
R6025 VSS.n11765 VSS 0.103002
R6026 VSS.n3424 VSS 0.102841
R6027 VSS.n5968 VSS.n4671 0.102547
R6028 VSS.n5787 VSS.n4680 0.102547
R6029 VSS.n5606 VSS.n4689 0.102547
R6030 VSS.n5426 VSS.n4700 0.102547
R6031 VSS.n5246 VSS.n4712 0.102547
R6032 VSS.n4575 VSS.n4572 0.102547
R6033 VSS.n3715 VSS.n3714 0.102547
R6034 VSS.n11684 VSS.n11569 0.102547
R6035 VSS.n11753 VSS.n11693 0.102547
R6036 VSS.n11782 VSS.n11779 0.102547
R6037 VSS.n11930 VSS.n11825 0.102547
R6038 VSS.n3445 VSS.n3397 0.102547
R6039 VSS.n12580 VSS.n3117 0.102547
R6040 VSS.n3213 VSS.n3187 0.102547
R6041 VSS.n10100 VSS 0.0999792
R6042 VSS VSS.n12206 0.0999792
R6043 VSS VSS.n11356 0.0994583
R6044 VSS.n9116 VSS 0.0989375
R6045 VSS VSS.n3674 0.0981562
R6046 VSS VSS.n3669 0.0981562
R6047 VSS.n11234 VSS 0.0981562
R6048 VSS.n11239 VSS 0.0981562
R6049 VSS.n11313 VSS.n11200 0.0974697
R6050 VSS VSS.n3664 0.0968542
R6051 VSS.n3654 VSS 0.0968542
R6052 VSS.n11244 VSS 0.0968542
R6053 VSS VSS.n11215 0.0968542
R6054 VSS.n11324 VSS.n11323 0.0963763
R6055 VSS.n6090 VSS 0.095417
R6056 VSS.n5908 VSS 0.095417
R6057 VSS.n4091 VSS.n4090 0.0949964
R6058 VSS.n708 VSS.n707 0.0947708
R6059 VSS.n10786 VSS.n4105 0.0895625
R6060 VSS.n3356 VSS.n3355 0.0885208
R6061 VSS VSS.n12042 0.0874792
R6062 VSS.n5187 VSS 0.0871183
R6063 VSS.n11143 VSS 0.0869583
R6064 VSS.n10135 VSS 0.0855622
R6065 VSS.n8049 VSS.n6238 0.0843334
R6066 VSS.n8011 VSS.n8008 0.0843334
R6067 VSS.n9546 VSS.n7589 0.0843334
R6068 VSS.n8527 VSS.n8364 0.0843334
R6069 VSS.n9148 VSS.n9144 0.0843334
R6070 VSS.n9232 VSS.n7596 0.0843334
R6071 VSS.n8939 VSS.n6252 0.0843334
R6072 VSS.n8900 VSS.n6245 0.0843334
R6073 VSS.n6847 VSS.n4653 0.0843334
R6074 VSS.n6914 VSS.n4649 0.0843334
R6075 VSS.n6987 VSS.n4645 0.0843334
R6076 VSS.n7046 VSS.n4640 0.0843334
R6077 VSS.n6768 VSS.n4657 0.0843334
R6078 VSS.n14251 VSS.n536 0.0843334
R6079 VSS.n13141 VSS.n1906 0.0843334
R6080 VSS.n1158 VSS.n616 0.0843334
R6081 VSS.n1119 VSS.n1115 0.0843334
R6082 VSS.n801 VSS.n797 0.0843334
R6083 VSS.n1402 VSS.n619 0.0843334
R6084 VSS.n2252 VSS.n1897 0.0843334
R6085 VSS.n2187 VSS.n1892 0.0843334
R6086 VSS.n2298 VSS.n1901 0.0843334
R6087 VSS.n12993 VSS.n2558 0.0843334
R6088 VSS.n12928 VSS.n2724 0.0843334
R6089 VSS.n12916 VSS.n2739 0.0843334
R6090 VSS.n12851 VSS.n2904 0.0843334
R6091 VSS.n12614 VSS.n2918 0.0843334
R6092 VSS.n8760 VSS.n8756 0.0843334
R6093 VSS.n9610 VSS.n7548 0.0843334
R6094 VSS.n9457 VSS.n9453 0.0843334
R6095 VSS.n9800 VSS.n9794 0.0843334
R6096 VSS.n9524 VSS.n7601 0.0843334
R6097 VSS.n9846 VSS.n7153 0.0843334
R6098 VSS.n9862 VSS.n7146 0.0843334
R6099 VSS.n8964 VSS.n6257 0.0843334
R6100 VSS.n7754 VSS.n6262 0.0843334
R6101 VSS.n9900 VSS.n6266 0.0843334
R6102 VSS.n10039 VSS.n4632 0.0843334
R6103 VSS.n11122 VSS.n3814 0.0843334
R6104 VSS.n10995 VSS.n3848 0.0843334
R6105 VSS.n10963 VSS.n3882 0.0843334
R6106 VSS.n10841 VSS.n3915 0.0843334
R6107 VSS.n14153 VSS.n607 0.0843334
R6108 VSS.n1360 VSS.n1354 0.0843334
R6109 VSS.n1637 VSS.n1636 0.0843334
R6110 VSS.n13868 VSS.n13862 0.0843334
R6111 VSS.n14123 VSS.n624 0.0843334
R6112 VSS.n14058 VSS.n1697 0.0843334
R6113 VSS.n13911 VSS.n1703 0.0843334
R6114 VSS.n13181 VSS.n1881 0.0843334
R6115 VSS.n12706 VSS.n12695 0.0843334
R6116 VSS.n13003 VSS.n2549 0.0843334
R6117 VSS.n2974 VSS.n2924 0.0843334
R6118 VSS.n13991 VSS.n1754 0.0843334
R6119 VSS.n13548 VSS.n1709 0.0843334
R6120 VSS.n10844 VSS.n3914 0.0842037
R6121 VSS.n13616 VSS.n13398 0.0842037
R6122 VSS.n9945 VSS.n6236 0.0842037
R6123 VSS.n8838 VSS.n8009 0.0842037
R6124 VSS.n7593 VSS.n7591 0.0842037
R6125 VSS.n9603 VSS.n9598 0.0842037
R6126 VSS.n8759 VSS.n8757 0.0842037
R6127 VSS.n8517 VSS.n8410 0.0842037
R6128 VSS.n9799 VSS.n9795 0.0842037
R6129 VSS.n9456 VSS.n9454 0.0842037
R6130 VSS.n9147 VSS.n9145 0.0842037
R6131 VSS.n9855 VSS.n7147 0.0842037
R6132 VSS.n7154 VSS.n7152 0.0842037
R6133 VSS.n9528 VSS.n7599 0.0842037
R6134 VSS.n9538 VSS.n9537 0.0842037
R6135 VSS.n9909 VSS.n6265 0.0842037
R6136 VSS.n9917 VSS.n6260 0.0842037
R6137 VSS.n9925 VSS.n6255 0.0842037
R6138 VSS.n9933 VSS.n6250 0.0842037
R6139 VSS.n9939 VSS.n6243 0.0842037
R6140 VSS.n10032 VSS.n4633 0.0842037
R6141 VSS.n10026 VSS.n10025 0.0842037
R6142 VSS.n10017 VSS.n10016 0.0842037
R6143 VSS.n10008 VSS.n10007 0.0842037
R6144 VSS.n9999 VSS.n9998 0.0842037
R6145 VSS.n9990 VSS.n9989 0.0842037
R6146 VSS.n3818 VSS.n3815 0.0842037
R6147 VSS.n3849 VSS.n3847 0.0842037
R6148 VSS.n3886 VSS.n3883 0.0842037
R6149 VSS.n14244 VSS.n538 0.0842037
R6150 VSS.n1907 VSS.n1905 0.0842037
R6151 VSS.n611 VSS.n609 0.0842037
R6152 VSS.n14145 VSS.n614 0.0842037
R6153 VSS.n1359 VSS.n1355 0.0842037
R6154 VSS.n1118 VSS.n1116 0.0842037
R6155 VSS.n13867 VSS.n13863 0.0842037
R6156 VSS.n1635 VSS.n1634 0.0842037
R6157 VSS.n800 VSS.n798 0.0842037
R6158 VSS.n14042 VSS.n1702 0.0842037
R6159 VSS.n14051 VSS.n1699 0.0842037
R6160 VSS.n14127 VSS.n622 0.0842037
R6161 VSS.n14137 VSS.n14136 0.0842037
R6162 VSS.n12699 VSS.n12696 0.0842037
R6163 VSS.n13174 VSS.n1883 0.0842037
R6164 VSS.n13168 VSS.n13167 0.0842037
R6165 VSS.n13159 VSS.n13158 0.0842037
R6166 VSS.n13150 VSS.n13149 0.0842037
R6167 VSS.n12843 VSS.n2917 0.0842037
R6168 VSS.n2914 VSS.n2906 0.0842037
R6169 VSS.n12920 VSS.n2737 0.0842037
R6170 VSS.n2734 VSS.n2726 0.0842037
R6171 VSS.n12997 VSS.n2556 0.0842037
R6172 VSS.n12426 VSS.n2551 0.0842037
R6173 VSS.n12838 VSS.n12837 0.0842037
R6174 VSS.n1755 VSS.n1753 0.0842037
R6175 VSS.n14037 VSS.n14036 0.0842037
R6176 VSS.n9360 VSS.n9359 0.0838333
R6177 VSS.n5727 VSS 0.0834875
R6178 VSS.n3292 VSS 0.0826231
R6179 VSS.n12810 VSS 0.0826231
R6180 VSS.n5367 VSS 0.0824502
R6181 VSS.n11993 VSS 0.0821044
R6182 VSS.n10739 VSS.n10734 0.0819275
R6183 VSS.n11692 VSS.n11691 0.08175
R6184 VSS.n8634 VSS 0.0810055
R6185 VSS.n8727 VSS 0.0810055
R6186 VSS.n9709 VSS 0.0810055
R6187 VSS.n7500 VSS 0.0810055
R6188 VSS.n9943 VSS.n9942 0.0808942
R6189 VSS.n8846 VSS.n8010 0.0808942
R6190 VSS.n9544 VSS.n7592 0.0808942
R6191 VSS.n9608 VSS.n9607 0.0808942
R6192 VSS.n8768 VSS.n8767 0.0808942
R6193 VSS.n8525 VSS.n8524 0.0808942
R6194 VSS.n9806 VSS.n9805 0.0808942
R6195 VSS.n9465 VSS.n9464 0.0808942
R6196 VSS.n9156 VSS.n9155 0.0808942
R6197 VSS.n9863 VSS.n7149 0.0808942
R6198 VSS.n9848 VSS.n7151 0.0808942
R6199 VSS.n7608 VSS.n7607 0.0808942
R6200 VSS.n9535 VSS.n9534 0.0808942
R6201 VSS.n9903 VSS.n9902 0.0808942
R6202 VSS.n9915 VSS.n9914 0.0808942
R6203 VSS.n9923 VSS.n9922 0.0808942
R6204 VSS.n9931 VSS.n9930 0.0808942
R6205 VSS.n9937 VSS.n9936 0.0808942
R6206 VSS.n10040 VSS.n4635 0.0808942
R6207 VSS.n10029 VSS.n10028 0.0808942
R6208 VSS.n10020 VSS.n10019 0.0808942
R6209 VSS.n10011 VSS.n10010 0.0808942
R6210 VSS.n10002 VSS.n10001 0.0808942
R6211 VSS.n9993 VSS.n9992 0.0808942
R6212 VSS.n11123 VSS.n3817 0.0808942
R6213 VSS.n10997 VSS.n3846 0.0808942
R6214 VSS.n10964 VSS.n3885 0.0808942
R6215 VSS.n10842 VSS.n3912 0.0808942
R6216 VSS.n14249 VSS.n541 0.0808942
R6217 VSS.n13143 VSS.n1904 0.0808942
R6218 VSS.n14151 VSS.n610 0.0808942
R6219 VSS.n14143 VSS.n14142 0.0808942
R6220 VSS.n1366 VSS.n1365 0.0808942
R6221 VSS.n1127 VSS.n1126 0.0808942
R6222 VSS.n13874 VSS.n13873 0.0808942
R6223 VSS.n1628 VSS.n1625 0.0808942
R6224 VSS.n809 VSS.n808 0.0808942
R6225 VSS.n13912 VSS.n1706 0.0808942
R6226 VSS.n14056 VSS.n14055 0.0808942
R6227 VSS.n14048 VSS.n625 0.0808942
R6228 VSS.n14134 VSS.n14133 0.0808942
R6229 VSS.n12707 VSS.n12698 0.0808942
R6230 VSS.n13179 VSS.n13178 0.0808942
R6231 VSS.n13171 VSS.n13170 0.0808942
R6232 VSS.n13162 VSS.n13161 0.0808942
R6233 VSS.n13153 VSS.n13152 0.0808942
R6234 VSS.n12612 VSS.n2921 0.0808942
R6235 VSS.n12849 VSS.n2907 0.0808942
R6236 VSS.n2909 VSS.n2740 0.0808942
R6237 VSS.n12926 VSS.n2727 0.0808942
R6238 VSS.n2729 VSS.n2559 0.0808942
R6239 VSS.n13001 VSS.n13000 0.0808942
R6240 VSS.n12835 VSS.n12834 0.0808942
R6241 VSS.n13993 VSS.n1752 0.0808942
R6242 VSS.n14034 VSS.n14033 0.0808942
R6243 VSS.n13625 VSS.n13624 0.0808942
R6244 VSS.n12464 VSS 0.0794216
R6245 VSS VSS.n6149 0.0794216
R6246 VSS VSS.n5966 0.0794216
R6247 VSS VSS.n5785 0.0794216
R6248 VSS VSS.n5604 0.0794216
R6249 VSS VSS.n5424 0.0794216
R6250 VSS VSS.n5244 0.0794216
R6251 VSS.n10101 VSS 0.0794216
R6252 VSS.n11144 VSS 0.0794216
R6253 VSS VSS.n12338 0.0794216
R6254 VSS VSS.n12205 0.0794216
R6255 VSS VSS.n12041 0.0794216
R6256 VSS VSS.n11928 0.0794216
R6257 VSS VSS.n3443 0.0794216
R6258 VSS VSS.n12578 0.0794216
R6259 VSS VSS.n3211 0.0794216
R6260 VSS.n3396 VSS.n3395 0.0791458
R6261 VSS.n5547 VSS 0.0789924
R6262 VSS.n10816 VSS 0.0785817
R6263 VSS.n10729 VSS.n10728 0.07852
R6264 VSS.n11778 VSS 0.076399
R6265 VSS VSS.n11125 0.0761666
R6266 VSS VSS.n3850 0.0761666
R6267 VSS VSS.n10966 0.0761666
R6268 VSS VSS.n3916 0.0761666
R6269 VSS VSS.n2550 0.0761666
R6270 VSS VSS.n3273 0.0761666
R6271 VSS VSS.n1756 0.0761666
R6272 VSS VSS.n13941 0.0761666
R6273 VSS VSS.n13627 0.0761666
R6274 VSS.n5154 VSS.n4706 0.0757941
R6275 VSS.n12550 VSS.n12549 0.0757941
R6276 VSS.n8075 VSS.n8049 0.0746667
R6277 VSS.n8795 VSS.n8008 0.0746667
R6278 VSS.n9547 VSS.n9546 0.0746667
R6279 VSS.n8528 VSS.n8527 0.0746667
R6280 VSS.n9144 VSS.n9143 0.0746667
R6281 VSS.n9233 VSS.n9232 0.0746667
R6282 VSS.n8940 VSS.n8939 0.0746667
R6283 VSS.n8901 VSS.n8900 0.0746667
R6284 VSS.n6848 VSS.n6847 0.0746667
R6285 VSS.n6915 VSS.n6914 0.0746667
R6286 VSS.n6988 VSS.n6987 0.0746667
R6287 VSS.n7047 VSS.n7046 0.0746667
R6288 VSS.n6769 VSS.n6768 0.0746667
R6289 VSS.n14252 VSS.n14251 0.0746667
R6290 VSS.n13141 VSS.n13140 0.0746667
R6291 VSS.n1159 VSS.n1158 0.0746667
R6292 VSS.n1115 VSS.n1114 0.0746667
R6293 VSS.n797 VSS.n796 0.0746667
R6294 VSS.n1403 VSS.n1402 0.0746667
R6295 VSS.n2253 VSS.n2252 0.0746667
R6296 VSS.n2188 VSS.n2187 0.0746667
R6297 VSS.n2299 VSS.n2298 0.0746667
R6298 VSS.n12993 VSS.n12992 0.0746667
R6299 VSS.n12929 VSS.n12928 0.0746667
R6300 VSS.n12916 VSS.n12915 0.0746667
R6301 VSS.n12852 VSS.n12851 0.0746667
R6302 VSS.n12615 VSS.n12614 0.0746667
R6303 VSS.n8756 VSS.n8755 0.0739167
R6304 VSS VSS.n8770 0.0739167
R6305 VSS VSS.n6738 0.0739167
R6306 VSS VSS.n8848 0.0739167
R6307 VSS VSS.n7590 0.0739167
R6308 VSS.n9611 VSS.n9610 0.0739167
R6309 VSS.n9597 VSS 0.0739167
R6310 VSS.n8409 VSS 0.0739167
R6311 VSS.n9453 VSS.n9452 0.0739167
R6312 VSS VSS.n9467 0.0739167
R6313 VSS.n9794 VSS.n9793 0.0739167
R6314 VSS VSS.n9808 0.0739167
R6315 VSS VSS.n9158 0.0739167
R6316 VSS.n9524 VSS.n9523 0.0739167
R6317 VSS.n9526 VSS 0.0739167
R6318 VSS.n9846 VSS.n9845 0.0739167
R6319 VSS VSS.n7155 0.0739167
R6320 VSS.n7241 VSS.n7146 0.0739167
R6321 VSS VSS.n9865 0.0739167
R6322 VSS VSS.n7919 0.0739167
R6323 VSS VSS.n6861 0.0739167
R6324 VSS.n8965 VSS.n8964 0.0739167
R6325 VSS VSS.n6928 0.0739167
R6326 VSS.n7755 VSS.n7754 0.0739167
R6327 VSS VSS.n7014 0.0739167
R6328 VSS.n9900 VSS.n9899 0.0739167
R6329 VSS.n7067 VSS 0.0739167
R6330 VSS VSS.n6813 0.0739167
R6331 VSS VSS.n5792 0.0739167
R6332 VSS VSS.n5611 0.0739167
R6333 VSS VSS.n5431 0.0739167
R6334 VSS VSS.n5251 0.0739167
R6335 VSS.n6461 VSS.n4632 0.0739167
R6336 VSS VSS.n10042 0.0739167
R6337 VSS VSS.n6048 0.0739167
R6338 VSS.n6384 VSS.n3814 0.0739167
R6339 VSS.n10995 VSS.n10994 0.0739167
R6340 VSS.n7330 VSS.n3882 0.0739167
R6341 VSS.n10841 VSS.n10840 0.0739167
R6342 VSS VSS.n537 0.0739167
R6343 VSS VSS.n1908 0.0739167
R6344 VSS.n14174 VSS.n14153 0.0739167
R6345 VSS VSS.n608 0.0739167
R6346 VSS VSS.n2325 0.0739167
R6347 VSS.n1354 VSS.n1353 0.0739167
R6348 VSS VSS.n1368 0.0739167
R6349 VSS VSS.n1129 0.0739167
R6350 VSS.n1637 VSS.n1624 0.0739167
R6351 VSS VSS.n1639 0.0739167
R6352 VSS.n13862 VSS.n13861 0.0739167
R6353 VSS VSS.n13876 0.0739167
R6354 VSS VSS.n811 0.0739167
R6355 VSS.n14123 VSS.n14122 0.0739167
R6356 VSS.n14125 VSS 0.0739167
R6357 VSS.n14059 VSS.n14058 0.0739167
R6358 VSS VSS.n1698 0.0739167
R6359 VSS.n13911 VSS.n13910 0.0739167
R6360 VSS VSS.n13914 0.0739167
R6361 VSS VSS.n2009 0.0739167
R6362 VSS VSS.n2666 0.0739167
R6363 VSS VSS.n2822 0.0739167
R6364 VSS.n13182 VSS.n13181 0.0739167
R6365 VSS VSS.n1882 0.0739167
R6366 VSS.n12695 VSS.n12694 0.0739167
R6367 VSS VSS.n12709 0.0739167
R6368 VSS VSS.n2588 0.0739167
R6369 VSS.n12995 VSS 0.0739167
R6370 VSS VSS.n2725 0.0739167
R6371 VSS.n12918 VSS 0.0739167
R6372 VSS VSS.n2905 0.0739167
R6373 VSS.n12611 VSS 0.0739167
R6374 VSS.n13004 VSS.n13003 0.0739167
R6375 VSS.n2999 VSS.n2974 0.0739167
R6376 VSS.n13991 VSS.n13990 0.0739167
R6377 VSS.n13549 VSS.n13548 0.0739167
R6378 VSS.n13397 VSS.n13396 0.0739167
R6379 VSS.n708 VSS 0.0734889
R6380 VSS.n12345 VSS.n12344 0.072375
R6381 VSS.n3356 VSS 0.0712123
R6382 VSS.n12339 VSS.n11683 0.0702917
R6383 VSS.n9360 VSS 0.0697521
R6384 VSS.n11692 VSS 0.0689647
R6385 VSS VSS.n12339 0.0687292
R6386 VSS.n3396 VSS 0.0681003
R6387 VSS.n995 VSS.n994 0.0676875
R6388 VSS.n12362 VSS.n12361 0.066646
R6389 VSS.n12345 VSS 0.0658527
R6390 VSS.n11921 VSS.n11916 0.0652425
R6391 VSS.n3206 VSS.n3184 0.065125
R6392 VSS.n13427 VSS.n13426 0.0650833
R6393 VSS.n1516 VSS.n1515 0.0650833
R6394 VSS.n13757 VSS.n13756 0.0650833
R6395 VSS.n13294 VSS.n13293 0.0650833
R6396 VSS.n11916 VSS.n11823 0.0647725
R6397 VSS.n1326 VSS.n1324 0.0645625
R6398 VSS.n3434 VSS.n3431 0.0635975
R6399 VSS.n12364 VSS 0.063
R6400 VSS.n8416 VSS 0.063
R6401 VSS.n8414 VSS 0.063
R6402 VSS.n8622 VSS 0.063
R6403 VSS.n8652 VSS 0.063
R6404 VSS.n9697 VSS 0.063
R6405 VSS.n9055 VSS 0.063
R6406 VSS.n3969 VSS 0.063
R6407 VSS.n6153 VSS 0.063
R6408 VSS.n4691 VSS 0.063
R6409 VSS.n4702 VSS 0.063
R6410 VSS.n4714 VSS 0.063
R6411 VSS.n4571 VSS 0.063
R6412 VSS.n3713 VSS 0.063
R6413 VSS.n11080 VSS 0.063
R6414 VSS.n4105 VSS 0.063
R6415 VSS.n10784 VSS 0.063
R6416 VSS.n4328 VSS 0.063
R6417 VSS.n4330 VSS 0.063
R6418 VSS.n4326 VSS 0.063
R6419 VSS.n10745 VSS 0.063
R6420 VSS.n10652 VSS 0.063
R6421 VSS.n10711 VSS 0.063
R6422 VSS.n12460 VSS 0.063
R6423 VSS.n11683 VSS 0.063
R6424 VSS.n11752 VSS 0.063
R6425 VSS.n11781 VSS 0.063
R6426 VSS.n11884 VSS 0.063
R6427 VSS.n3399 VSS 0.063
R6428 VSS.n3173 VSS 0.063
R6429 VSS.n12813 VSS 0.063
R6430 VSS.n3191 VSS 0.063
R6431 VSS.n13427 VSS 0.063
R6432 VSS.n10745 VSS.n10744 0.0609167
R6433 VSS VSS.n11806 0.0607775
R6434 VSS VSS.n11412 0.0603958
R6435 VSS.n11393 VSS 0.0603958
R6436 VSS.n11375 VSS 0.0603958
R6437 VSS.n11357 VSS 0.0603958
R6438 VSS VSS.n11354 0.0603958
R6439 VSS VSS.n11353 0.0603958
R6440 VSS.n11344 VSS 0.0603958
R6441 VSS.n3673 VSS 0.0603958
R6442 VSS.n3670 VSS 0.0603958
R6443 VSS.n3668 VSS 0.0603958
R6444 VSS.n3665 VSS 0.0603958
R6445 VSS.n3658 VSS 0.0603958
R6446 VSS VSS.n3657 0.0603958
R6447 VSS.n3648 VSS 0.0603958
R6448 VSS VSS.n3646 0.0603958
R6449 VSS VSS.n11235 0.0603958
R6450 VSS.n11236 VSS 0.0603958
R6451 VSS.n11240 VSS 0.0603958
R6452 VSS.n11243 VSS 0.0603958
R6453 VSS VSS.n11250 0.0603958
R6454 VSS.n11251 VSS 0.0603958
R6455 VSS.n11258 VSS 0.0603958
R6456 VSS VSS.n11212 0.0603958
R6457 VSS.n3353 VSS.n3175 0.0603075
R6458 VSS.n3207 VSS.n3206 0.0603075
R6459 VSS.n11182 VSS.n11181 0.0600725
R6460 VSS.n3385 VSS.n3384 0.0598752
R6461 VSS.n1246 VSS.n1245 0.0593542
R6462 VSS VSS.n12463 0.0593235
R6463 VSS.n1515 VSS 0.0593235
R6464 VSS.n6150 VSS 0.0593235
R6465 VSS.n8429 VSS 0.0593235
R6466 VSS.n8625 VSS 0.0593235
R6467 VSS.n8711 VSS 0.0593235
R6468 VSS.n9700 VSS 0.0593235
R6469 VSS.n9116 VSS 0.0593235
R6470 VSS.n7482 VSS 0.0593235
R6471 VSS.n4028 VSS 0.0593235
R6472 VSS.n9770 VSS 0.0593235
R6473 VSS.n9424 VSS 0.0593235
R6474 VSS.n5967 VSS 0.0593235
R6475 VSS.n5786 VSS 0.0593235
R6476 VSS.n5605 VSS 0.0593235
R6477 VSS.n5425 VSS 0.0593235
R6478 VSS.n5245 VSS 0.0593235
R6479 VSS VSS.n10100 0.0593235
R6480 VSS VSS.n11143 0.0593235
R6481 VSS.n10786 VSS 0.0593235
R6482 VSS.n10744 VSS 0.0593235
R6483 VSS.n10715 VSS 0.0593235
R6484 VSS.n994 VSS 0.0593235
R6485 VSS.n14360 VSS 0.0593235
R6486 VSS.n14370 VSS 0.0593235
R6487 VSS.n1074 VSS 0.0593235
R6488 VSS.n1245 VSS 0.0593235
R6489 VSS.n1324 VSS 0.0593235
R6490 VSS.n463 VSS 0.0593235
R6491 VSS.n13756 VSS 0.0593235
R6492 VSS.n13293 VSS 0.0593235
R6493 VSS.n13371 VSS 0.0593235
R6494 VSS.n13836 VSS 0.0593235
R6495 VSS.n1596 VSS 0.0593235
R6496 VSS.n12339 VSS 0.0593235
R6497 VSS.n12206 VSS 0.0593235
R6498 VSS.n12042 VSS 0.0593235
R6499 VSS.n11929 VSS 0.0593235
R6500 VSS.n3444 VSS 0.0593235
R6501 VSS.n12579 VSS 0.0593235
R6502 VSS.n3212 VSS 0.0593235
R6503 VSS.n13426 VSS 0.0593235
R6504 VSS.n11774 VSS.n11772 0.0584275
R6505 VSS.n1076 VSS.n1074 0.0583125
R6506 VSS.n3354 VSS.n3353 0.05737
R6507 VSS.n12274 VSS.n12273 0.057271
R6508 VSS.n6090 VSS.n6089 0.0572708
R6509 VSS.n5908 VSS.n5907 0.0572708
R6510 VSS.n11118 VSS.n11117 0.0564896
R6511 VSS.n11004 VSS.n11003 0.0564896
R6512 VSS.n10959 VSS.n10958 0.0564896
R6513 VSS.n4355 VSS.n4354 0.0564896
R6514 VSS.n4439 VSS.n4438 0.0564896
R6515 VSS.n12829 VSS.n12828 0.0564896
R6516 VSS.n14000 VSS.n13999 0.0564896
R6517 VSS.n14028 VSS.n14027 0.0564896
R6518 VSS.n13574 VSS.n13511 0.0560583
R6519 VSS.n13963 VSS.n13962 0.0560583
R6520 VSS.n12751 VSS.n2944 0.0560583
R6521 VSS.n7341 VSS.n7279 0.0560583
R6522 VSS.n10984 VSS.n10983 0.0560583
R6523 VSS.n6395 VSS.n6333 0.0560583
R6524 VSS.n7998 VSS.n7941 0.0560583
R6525 VSS.n8508 VSS.n8185 0.0560583
R6526 VSS.n8407 VSS.n8217 0.0560583
R6527 VSS.n8284 VSS.n7568 0.0560583
R6528 VSS.n6736 VSS.n6676 0.0560583
R6529 VSS.n9972 VSS.n9971 0.0560583
R6530 VSS.n8156 VSS.n8016 0.0560583
R6531 VSS.n8870 VSS.n8004 0.0560583
R6532 VSS.n9207 VSS.n9188 0.0560583
R6533 VSS.n9290 VSS.n9288 0.0560583
R6534 VSS.n9468 VSS.n7183 0.0560583
R6535 VSS.n7379 VSS.n7190 0.0560583
R6536 VSS.n7894 VSS.n7851 0.0560583
R6537 VSS.n7636 VSS.n7610 0.0560583
R6538 VSS.n7671 VSS.n7645 0.0560583
R6539 VSS.n9887 VSS.n9886 0.0560583
R6540 VSS.n6794 VSS.n6629 0.0560583
R6541 VSS.n6862 VSS.n6581 0.0560583
R6542 VSS.n6929 VSS.n6540 0.0560583
R6543 VSS.n7015 VSS.n6483 0.0560583
R6544 VSS.n6449 VSS.n6448 0.0560583
R6545 VSS.n10773 VSS.n4107 0.0560583
R6546 VSS.n4298 VSS.n4297 0.0560583
R6547 VSS.n4410 VSS.n4162 0.0560583
R6548 VSS.n954 VSS.n882 0.0560583
R6549 VSS.n2323 VSS.n1948 0.0560583
R6550 VSS.n14234 VSS.n545 0.0560583
R6551 VSS.n14206 VSS.n584 0.0560583
R6552 VSS.n13028 VSS.n2500 0.0560583
R6553 VSS.n13058 VSS.n2461 0.0560583
R6554 VSS.n2447 VSS.n2392 0.0560583
R6555 VSS.n13128 VSS.n13127 0.0560583
R6556 VSS.n1195 VSS.n841 0.0560583
R6557 VSS.n1460 VSS.n1458 0.0560583
R6558 VSS.n1666 VSS.n1640 0.0560583
R6559 VSS.n13898 VSS.n13897 0.0560583
R6560 VSS.n2053 VSS.n2052 0.0560583
R6561 VSS.n2102 VSS.n2101 0.0560583
R6562 VSS.n2132 VSS.n1853 0.0560583
R6563 VSS.n13925 VSS.n1816 0.0560583
R6564 VSS.n2660 VSS.n2659 0.0560583
R6565 VSS.n2693 VSS.n2667 0.0560583
R6566 VSS.n2841 VSS.n2840 0.0560583
R6567 VSS.n2873 VSS.n2847 0.0560583
R6568 VSS.n12720 VSS.n3021 0.0560583
R6569 VSS.n11772 VSS.n11689 0.0558425
R6570 VSS.n11807 VSS 0.055725
R6571 VSS.n3431 VSS.n3394 0.0553725
R6572 VSS.n9355 VSS.n9354 0.0551877
R6573 VSS.n13590 VSS.n13589 0.0545568
R6574 VSS.n1763 VSS.n1745 0.0545568
R6575 VSS.n12801 VSS.n2930 0.0545568
R6576 VSS.n2902 VSS.n2842 0.0545568
R6577 VSS.n2811 VSS.n2789 0.0545568
R6578 VSS.n10896 VSS.n3893 0.0545568
R6579 VSS.n10942 VSS.n10941 0.0545568
R6580 VSS.n11047 VSS.n3825 0.0545568
R6581 VSS.n6985 VSS.n6561 0.0545568
R6582 VSS.n9563 VSS.n9562 0.0545568
R6583 VSS.n8388 VSS.n8187 0.0545568
R6584 VSS.n8772 VSS.n8219 0.0545568
R6585 VSS.n8237 VSS.n8218 0.0545568
R6586 VSS.n8793 VSS.n8194 0.0545568
R6587 VSS.n9982 VSS.n6213 0.0545568
R6588 VSS.n6746 VSS.n6745 0.0545568
R6589 VSS.n6766 VSS.n6692 0.0545568
R6590 VSS.n8099 VSS.n8037 0.0545568
R6591 VSS.n8088 VSS.n8036 0.0545568
R6592 VSS.n8147 VSS.n8146 0.0545568
R6593 VSS.n8073 VSS.n8001 0.0545568
R6594 VSS.n8878 VSS.n8877 0.0545568
R6595 VSS.n8898 VSS.n7948 0.0545568
R6596 VSS.n8811 VSS.n8186 0.0545568
R6597 VSS.n8831 VSS.n8162 0.0545568
R6598 VSS.n9549 VSS.n7567 0.0545568
R6599 VSS.n9595 VSS.n7551 0.0545568
R6600 VSS.n9294 VSS.n9291 0.0545568
R6601 VSS.n9521 VSS.n8994 0.0545568
R6602 VSS.n9509 VSS.n9508 0.0545568
R6603 VSS.n7216 VSS.n7184 0.0545568
R6604 VSS.n9843 VSS.n7158 0.0545568
R6605 VSS.n9831 VSS.n9830 0.0545568
R6606 VSS.n7260 VSS.n7211 0.0545568
R6607 VSS.n7364 VSS.n7262 0.0545568
R6608 VSS.n7312 VSS.n7261 0.0545568
R6609 VSS.n9269 VSS.n9160 0.0545568
R6610 VSS.n9235 VSS.n9187 0.0545568
R6611 VSS.n9260 VSS.n9246 0.0545568
R6612 VSS.n7849 VSS.n7808 0.0545568
R6613 VSS.n8942 VSS.n7850 0.0545568
R6614 VSS.n8954 VSS.n8953 0.0545568
R6615 VSS.n7729 VSS.n7640 0.0545568
R6616 VSS.n8983 VSS.n8982 0.0545568
R6617 VSS.n7804 VSS.n7803 0.0545568
R6618 VSS.n7694 VSS.n7675 0.0545568
R6619 VSS.n7773 VSS.n7772 0.0545568
R6620 VSS.n7725 VSS.n7724 0.0545568
R6621 VSS.n9897 VSS.n7070 0.0545568
R6622 VSS.n7134 VSS.n7089 0.0545568
R6623 VSS.n7112 VSS.n7088 0.0545568
R6624 VSS.n7939 VSS.n7936 0.0545568
R6625 VSS.n8917 VSS.n7940 0.0545568
R6626 VSS.n8937 VSS.n7872 0.0545568
R6627 VSS.n6912 VSS.n6609 0.0545568
R6628 VSS.n6850 VSS.n6628 0.0545568
R6629 VSS.n6903 VSS.n6902 0.0545568
R6630 VSS.n6917 VSS.n6580 0.0545568
R6631 VSS.n6976 VSS.n6975 0.0545568
R6632 VSS.n6538 VSS.n6510 0.0545568
R6633 VSS.n6990 VSS.n6539 0.0545568
R6634 VSS.n7036 VSS.n7035 0.0545568
R6635 VSS.n6481 VSS.n6292 0.0545568
R6636 VSS.n7049 VSS.n6482 0.0545568
R6637 VSS.n7065 VSS.n6271 0.0545568
R6638 VSS.n6459 VSS.n6297 0.0545568
R6639 VSS.n6418 VSS.n6316 0.0545568
R6640 VSS.n6366 VSS.n6315 0.0545568
R6641 VSS.n6835 VSS.n6834 0.0545568
R6642 VSS.n6782 VSS.n6675 0.0545568
R6643 VSS.n6845 VSS.n6657 0.0545568
R6644 VSS.n6386 VSS.n6347 0.0545568
R6645 VSS.n11025 VSS.n11024 0.0545568
R6646 VSS.n10992 VSS.n3853 0.0545568
R6647 VSS.n10952 VSS.n10900 0.0545568
R6648 VSS.n7332 VSS.n7293 0.0545568
R6649 VSS.n10874 VSS.n10873 0.0545568
R6650 VSS.n4444 VSS.n4132 0.0545568
R6651 VSS.n4401 VSS.n4400 0.0545568
R6652 VSS.n4377 VSS.n4376 0.0545568
R6653 VSS.n4266 VSS.n4259 0.0545568
R6654 VSS.n4323 VSS.n4262 0.0545568
R6655 VSS.n4349 VSS.n4230 0.0545568
R6656 VSS.n4208 VSS.n4201 0.0545568
R6657 VSS.n4432 VSS.n4131 0.0545568
R6658 VSS.n10770 VSS.n10769 0.0545568
R6659 VSS.n1400 VSS.n862 0.0545568
R6660 VSS.n14225 VSS.n14224 0.0545568
R6661 VSS.n1136 VSS.n1135 0.0545568
R6662 VSS.n1156 VSS.n910 0.0545568
R6663 VSS.n14197 VSS.n14196 0.0545568
R6664 VSS.n12419 VSS.n2480 0.0545568
R6665 VSS.n13042 VSS.n2482 0.0545568
R6666 VSS.n2531 VSS.n2481 0.0545568
R6667 VSS.n13097 VSS.n2350 0.0545568
R6668 VSS.n2391 VSS.n2390 0.0545568
R6669 VSS.n13091 VSS.n13090 0.0545568
R6670 VSS.n13138 VSS.n1911 0.0545568
R6671 VSS.n2327 VSS.n1930 0.0545568
R6672 VSS.n2296 VSS.n1929 0.0545568
R6673 VSS.n14157 VSS.n14154 0.0545568
R6674 VSS.n2419 VSS.n2403 0.0545568
R6675 VSS.n1161 VSS.n881 0.0545568
R6676 VSS.n1391 VSS.n1390 0.0545568
R6677 VSS.n1672 VSS.n1461 0.0545568
R6678 VSS.n14120 VSS.n628 0.0545568
R6679 VSS.n14108 VSS.n14107 0.0545568
R6680 VSS.n13694 VSS.n13672 0.0545568
R6681 VSS.n14077 VSS.n14076 0.0545568
R6682 VSS.n13702 VSS.n13652 0.0545568
R6683 VSS.n13908 VSS.n13204 0.0545568
R6684 VSS.n13640 VSS.n13223 0.0545568
R6685 VSS.n13530 VSS.n13222 0.0545568
R6686 VSS.n1439 VSS.n813 0.0545568
R6687 VSS.n1405 VSS.n840 0.0545568
R6688 VSS.n1430 VSS.n1416 0.0545568
R6689 VSS.n2206 VSS.n2054 0.0545568
R6690 VSS.n2250 VSS.n1983 0.0545568
R6691 VSS.n2238 VSS.n2237 0.0545568
R6692 VSS.n2122 VSS.n2103 0.0545568
R6693 VSS.n2185 VSS.n2058 0.0545568
R6694 VSS.n2173 VSS.n2172 0.0545568
R6695 VSS.n12645 VSS.n1851 0.0545568
R6696 VSS.n13184 VSS.n1852 0.0545568
R6697 VSS.n13200 VSS.n1831 0.0545568
R6698 VSS.n12692 VSS.n1813 0.0545568
R6699 VSS.n13931 VSS.n1771 0.0545568
R6700 VSS.n1812 VSS.n1811 0.0545568
R6701 VSS.n2033 VSS.n1977 0.0545568
R6702 VSS.n2317 VSS.n2316 0.0545568
R6703 VSS.n2276 VSS.n2275 0.0545568
R6704 VSS.n2722 VSS.n2661 0.0545568
R6705 VSS.n12990 VSS.n2562 0.0545568
R6706 VSS.n12978 VSS.n12977 0.0545568
R6707 VSS.n12947 VSS.n12946 0.0545568
R6708 VSS.n2820 VSS.n2770 0.0545568
R6709 VSS.n12913 VSS.n2743 0.0545568
R6710 VSS.n12901 VSS.n12900 0.0545568
R6711 VSS.n12635 VSS.n3056 0.0545568
R6712 VSS.n12870 VSS.n12869 0.0545568
R6713 VSS.n12643 VSS.n3036 0.0545568
R6714 VSS.n3083 VSS.n3018 0.0545568
R6715 VSS.n12726 VSS.n2949 0.0545568
R6716 VSS.n3017 VSS.n3016 0.0545568
R6717 VSS.n2640 VSS.n2590 0.0545568
R6718 VSS.n13022 VSS.n13021 0.0545568
R6719 VSS.n2631 VSS.n2630 0.0545568
R6720 VSS.n2997 VSS.n2943 0.0545568
R6721 VSS.n12779 VSS.n12778 0.0545568
R6722 VSS.n13988 VSS.n1759 0.0545568
R6723 VSS.n14021 VSS.n1716 0.0545568
R6724 VSS.n13551 VSS.n13510 0.0545568
R6725 VSS.n13608 VSS.n13481 0.0545568
R6726 VSS.n11760 VSS 0.0542143
R6727 VSS.n3 VSS 0.0539905
R6728 VSS.n3340 VSS 0.0539905
R6729 VSS.n11785 VSS 0.0539905
R6730 VSS.n11534 VSS 0.0539905
R6731 VSS.n3418 VSS 0.0537667
R6732 VSS.n11904 VSS 0.0537667
R6733 VSS.n3616 VSS 0.0537667
R6734 VSS.n12351 VSS.n11547 0.0537275
R6735 VSS.n13627 VSS.n13626 0.0530835
R6736 VSS.n13941 VSS.n1708 0.0530835
R6737 VSS.n13992 VSS.n1756 0.0530835
R6738 VSS.n3273 VSS.n2923 0.0530835
R6739 VSS.n13002 VSS.n2550 0.0530835
R6740 VSS.n10843 VSS.n3916 0.0530835
R6741 VSS.n10966 VSS.n10965 0.0530835
R6742 VSS.n10996 VSS.n3850 0.0530835
R6743 VSS.n11125 VSS.n11124 0.0530835
R6744 VSS.n11125 VSS 0.0530835
R6745 VSS.n3850 VSS 0.0530835
R6746 VSS.n10966 VSS 0.0530835
R6747 VSS.n3916 VSS 0.0530835
R6748 VSS VSS.n2550 0.0530835
R6749 VSS.n3273 VSS 0.0530835
R6750 VSS.n1756 VSS 0.0530835
R6751 VSS.n13941 VSS 0.0530835
R6752 VSS.n13627 VSS 0.0530835
R6753 VSS VSS.n8759 0.0530834
R6754 VSS.n9945 VSS 0.0530834
R6755 VSS VSS.n8838 0.0530834
R6756 VSS VSS.n7593 0.0530834
R6757 VSS VSS.n9603 0.0530834
R6758 VSS VSS.n8517 0.0530834
R6759 VSS VSS.n9456 0.0530834
R6760 VSS VSS.n9799 0.0530834
R6761 VSS VSS.n9147 0.0530834
R6762 VSS.n9528 VSS 0.0530834
R6763 VSS VSS.n7152 0.0530834
R6764 VSS VSS.n9855 0.0530834
R6765 VSS.n9538 VSS 0.0530834
R6766 VSS.n9933 VSS 0.0530834
R6767 VSS.n9925 VSS 0.0530834
R6768 VSS.n9917 VSS 0.0530834
R6769 VSS.n9909 VSS 0.0530834
R6770 VSS.n9939 VSS 0.0530834
R6771 VSS.n9998 VSS 0.0530834
R6772 VSS.n10007 VSS 0.0530834
R6773 VSS.n10016 VSS 0.0530834
R6774 VSS.n10025 VSS 0.0530834
R6775 VSS VSS.n10032 0.0530834
R6776 VSS.n9989 VSS 0.0530834
R6777 VSS VSS.n3818 0.0530834
R6778 VSS VSS.n3847 0.0530834
R6779 VSS VSS.n3886 0.0530834
R6780 VSS VSS.n3914 0.0530834
R6781 VSS VSS.n14244 0.0530834
R6782 VSS VSS.n1905 0.0530834
R6783 VSS VSS.n611 0.0530834
R6784 VSS.n14145 VSS 0.0530834
R6785 VSS VSS.n1359 0.0530834
R6786 VSS VSS.n1118 0.0530834
R6787 VSS.n1634 VSS 0.0530834
R6788 VSS VSS.n13867 0.0530834
R6789 VSS VSS.n800 0.0530834
R6790 VSS.n14127 VSS 0.0530834
R6791 VSS VSS.n14051 0.0530834
R6792 VSS.n14042 VSS 0.0530834
R6793 VSS.n14137 VSS 0.0530834
R6794 VSS.n13158 VSS 0.0530834
R6795 VSS.n13167 VSS 0.0530834
R6796 VSS VSS.n13174 0.0530834
R6797 VSS VSS.n12699 0.0530834
R6798 VSS.n13149 VSS 0.0530834
R6799 VSS.n12997 VSS 0.0530834
R6800 VSS VSS.n2734 0.0530834
R6801 VSS.n12920 VSS 0.0530834
R6802 VSS VSS.n2914 0.0530834
R6803 VSS.n12843 VSS 0.0530834
R6804 VSS.n12426 VSS 0.0530834
R6805 VSS.n12838 VSS 0.0530834
R6806 VSS VSS.n1753 0.0530834
R6807 VSS.n14037 VSS 0.0530834
R6808 VSS VSS.n13616 0.0530834
R6809 VSS.n12613 VSS.n12611 0.0530834
R6810 VSS.n12850 VSS.n2905 0.0530834
R6811 VSS.n12918 VSS.n12917 0.0530834
R6812 VSS.n12927 VSS.n2725 0.0530834
R6813 VSS.n12995 VSS.n12994 0.0530834
R6814 VSS.n2588 VSS.n1900 0.0530834
R6815 VSS.n12709 VSS.n12708 0.0530834
R6816 VSS.n13180 VSS.n1882 0.0530834
R6817 VSS.n2822 VSS.n1891 0.0530834
R6818 VSS.n2666 VSS.n1896 0.0530834
R6819 VSS.n2009 VSS.n620 0.0530834
R6820 VSS.n13914 VSS.n13913 0.0530834
R6821 VSS.n14057 VSS.n1698 0.0530834
R6822 VSS.n14125 VSS.n14124 0.0530834
R6823 VSS.n811 VSS.n810 0.0530834
R6824 VSS.n13876 VSS.n13875 0.0530834
R6825 VSS.n1639 VSS.n1638 0.0530834
R6826 VSS.n6048 VSS.n4656 0.0530834
R6827 VSS.n10042 VSS.n10041 0.0530834
R6828 VSS.n5251 VSS.n4639 0.0530834
R6829 VSS.n5431 VSS.n4644 0.0530834
R6830 VSS.n5611 VSS.n4648 0.0530834
R6831 VSS.n5792 VSS.n4652 0.0530834
R6832 VSS.n6813 VSS.n6246 0.0530834
R6833 VSS.n9901 VSS.n7067 0.0530834
R6834 VSS.n7014 VSS.n6263 0.0530834
R6835 VSS.n6928 VSS.n6258 0.0530834
R6836 VSS.n6861 VSS.n6253 0.0530834
R6837 VSS.n7919 VSS.n7597 0.0530834
R6838 VSS.n9865 VSS.n9864 0.0530834
R6839 VSS.n9847 VSS.n7155 0.0530834
R6840 VSS.n9526 VSS.n9525 0.0530834
R6841 VSS.n9158 VSS.n9157 0.0530834
R6842 VSS.n9808 VSS.n9807 0.0530834
R6843 VSS.n9467 VSS.n9466 0.0530834
R6844 VSS.n8526 VSS.n8409 0.0530834
R6845 VSS.n9609 VSS.n9597 0.0530834
R6846 VSS.n8770 VSS.n8769 0.0530834
R6847 VSS.n8770 VSS 0.0530834
R6848 VSS.n8848 VSS.n8847 0.0530834
R6849 VSS.n6738 VSS.n6239 0.0530834
R6850 VSS.n6738 VSS 0.0530834
R6851 VSS.n8848 VSS 0.0530834
R6852 VSS.n9545 VSS.n7590 0.0530834
R6853 VSS VSS.n7590 0.0530834
R6854 VSS VSS.n9597 0.0530834
R6855 VSS VSS.n8409 0.0530834
R6856 VSS.n9467 VSS 0.0530834
R6857 VSS.n9808 VSS 0.0530834
R6858 VSS.n9158 VSS 0.0530834
R6859 VSS VSS.n9526 0.0530834
R6860 VSS.n7155 VSS 0.0530834
R6861 VSS.n9865 VSS 0.0530834
R6862 VSS.n7919 VSS 0.0530834
R6863 VSS.n6861 VSS 0.0530834
R6864 VSS.n6928 VSS 0.0530834
R6865 VSS.n7014 VSS 0.0530834
R6866 VSS.n7067 VSS 0.0530834
R6867 VSS.n6813 VSS 0.0530834
R6868 VSS.n5792 VSS 0.0530834
R6869 VSS.n5611 VSS 0.0530834
R6870 VSS.n5431 VSS 0.0530834
R6871 VSS.n5251 VSS 0.0530834
R6872 VSS.n10042 VSS 0.0530834
R6873 VSS.n6048 VSS 0.0530834
R6874 VSS.n1129 VSS.n1128 0.0530834
R6875 VSS.n1368 VSS.n1367 0.0530834
R6876 VSS.n14250 VSS.n537 0.0530834
R6877 VSS VSS.n537 0.0530834
R6878 VSS.n14152 VSS.n608 0.0530834
R6879 VSS.n13142 VSS.n1908 0.0530834
R6880 VSS.n1908 VSS 0.0530834
R6881 VSS VSS.n608 0.0530834
R6882 VSS.n2325 VSS.n617 0.0530834
R6883 VSS.n2325 VSS 0.0530834
R6884 VSS.n1368 VSS 0.0530834
R6885 VSS.n1129 VSS 0.0530834
R6886 VSS.n1639 VSS 0.0530834
R6887 VSS.n13876 VSS 0.0530834
R6888 VSS.n811 VSS 0.0530834
R6889 VSS VSS.n14125 0.0530834
R6890 VSS VSS.n1698 0.0530834
R6891 VSS.n13914 VSS 0.0530834
R6892 VSS.n2009 VSS 0.0530834
R6893 VSS.n2666 VSS 0.0530834
R6894 VSS.n2822 VSS 0.0530834
R6895 VSS VSS.n1882 0.0530834
R6896 VSS.n12709 VSS 0.0530834
R6897 VSS.n2588 VSS 0.0530834
R6898 VSS VSS.n12995 0.0530834
R6899 VSS VSS.n2725 0.0530834
R6900 VSS VSS.n12918 0.0530834
R6901 VSS VSS.n2905 0.0530834
R6902 VSS.n12611 VSS 0.0530834
R6903 VSS.n1501 VSS 0.0526476
R6904 VSS.n13750 VSS 0.0526476
R6905 VSS.n13419 VSS 0.0526476
R6906 VSS.n13288 VSS 0.0526476
R6907 VSS.n1238 VSS 0.0526476
R6908 VSS.n8762 VSS 0.0525833
R6909 VSS VSS.n6237 0.0525833
R6910 VSS VSS.n8844 0.0525833
R6911 VSS VSS.n9542 0.0525833
R6912 VSS.n9604 VSS 0.0525833
R6913 VSS.n8519 VSS 0.0525833
R6914 VSS.n9459 VSS 0.0525833
R6915 VSS.n9802 VSS 0.0525833
R6916 VSS.n9150 VSS 0.0525833
R6917 VSS VSS.n7600 0.0525833
R6918 VSS.n9850 VSS 0.0525833
R6919 VSS VSS.n9861 0.0525833
R6920 VSS.n9530 VSS 0.0525833
R6921 VSS VSS.n6251 0.0525833
R6922 VSS VSS.n6256 0.0525833
R6923 VSS VSS.n6261 0.0525833
R6924 VSS VSS.n9908 0.0525833
R6925 VSS VSS.n6244 0.0525833
R6926 VSS VSS.n4651 0.0525833
R6927 VSS VSS.n4647 0.0525833
R6928 VSS VSS.n4643 0.0525833
R6929 VSS VSS.n4641 0.0525833
R6930 VSS VSS.n10038 0.0525833
R6931 VSS VSS.n4655 0.0525833
R6932 VSS VSS.n11121 0.0525833
R6933 VSS.n10999 VSS 0.0525833
R6934 VSS VSS.n10962 0.0525833
R6935 VSS.n10846 VSS 0.0525833
R6936 VSS VSS.n14247 0.0525833
R6937 VSS.n13146 VSS 0.0525833
R6938 VSS VSS.n14149 0.0525833
R6939 VSS VSS.n615 0.0525833
R6940 VSS.n1362 VSS 0.0525833
R6941 VSS.n1121 VSS 0.0525833
R6942 VSS VSS.n1631 0.0525833
R6943 VSS.n13870 VSS 0.0525833
R6944 VSS.n803 VSS 0.0525833
R6945 VSS VSS.n623 0.0525833
R6946 VSS.n14052 VSS 0.0525833
R6947 VSS VSS.n14041 0.0525833
R6948 VSS.n14129 VSS 0.0525833
R6949 VSS VSS.n1895 0.0525833
R6950 VSS VSS.n1893 0.0525833
R6951 VSS.n13175 VSS 0.0525833
R6952 VSS VSS.n12705 0.0525833
R6953 VSS VSS.n1899 0.0525833
R6954 VSS VSS.n2557 0.0525833
R6955 VSS VSS.n12924 0.0525833
R6956 VSS VSS.n2738 0.0525833
R6957 VSS VSS.n12847 0.0525833
R6958 VSS VSS.n12842 0.0525833
R6959 VSS VSS.n12425 0.0525833
R6960 VSS.n12831 VSS 0.0525833
R6961 VSS.n13995 VSS 0.0525833
R6962 VSS.n14030 VSS 0.0525833
R6963 VSS.n13619 VSS 0.0525833
R6964 VSS.n2298 VSS.n1900 0.0525626
R6965 VSS.n1402 VSS.n620 0.0525626
R6966 VSS.n810 VSS.n797 0.0525626
R6967 VSS.n6768 VSS.n4656 0.0525626
R6968 VSS.n8900 VSS.n6246 0.0525626
R6969 VSS.n9232 VSS.n7597 0.0525626
R6970 VSS.n9157 VSS.n9144 0.0525626
R6971 VSS.n8527 VSS.n8526 0.0525626
R6972 VSS.n8049 VSS.n6239 0.0525626
R6973 VSS.n8847 VSS.n8008 0.0525626
R6974 VSS.n9546 VSS.n9545 0.0525626
R6975 VSS.n8939 VSS.n6253 0.0525626
R6976 VSS.n6847 VSS.n4652 0.0525626
R6977 VSS.n6914 VSS.n4648 0.0525626
R6978 VSS.n6987 VSS.n4644 0.0525626
R6979 VSS.n7046 VSS.n4639 0.0525626
R6980 VSS.n1128 VSS.n1115 0.0525626
R6981 VSS.n14251 VSS.n14250 0.0525626
R6982 VSS.n13142 VSS.n13141 0.0525626
R6983 VSS.n1158 VSS.n617 0.0525626
R6984 VSS.n2252 VSS.n1896 0.0525626
R6985 VSS.n2187 VSS.n1891 0.0525626
R6986 VSS.n12994 VSS.n12993 0.0525626
R6987 VSS.n12928 VSS.n12927 0.0525626
R6988 VSS.n12917 VSS.n12916 0.0525626
R6989 VSS.n12851 VSS.n12850 0.0525626
R6990 VSS.n12614 VSS.n12613 0.0525626
R6991 VSS.n13626 VSS.n13397 0.0525625
R6992 VSS.n13548 VSS.n1708 0.0525625
R6993 VSS.n13992 VSS.n13991 0.0525625
R6994 VSS.n2974 VSS.n2923 0.0525625
R6995 VSS.n13003 VSS.n13002 0.0525625
R6996 VSS.n12708 VSS.n12695 0.0525625
R6997 VSS.n13181 VSS.n13180 0.0525625
R6998 VSS.n13913 VSS.n13911 0.0525625
R6999 VSS.n14058 VSS.n14057 0.0525625
R7000 VSS.n14124 VSS.n14123 0.0525625
R7001 VSS.n13875 VSS.n13862 0.0525625
R7002 VSS.n1638 VSS.n1637 0.0525625
R7003 VSS.n10843 VSS.n10841 0.0525625
R7004 VSS.n10965 VSS.n3882 0.0525625
R7005 VSS.n10996 VSS.n10995 0.0525625
R7006 VSS.n11124 VSS.n3814 0.0525625
R7007 VSS.n10041 VSS.n4632 0.0525625
R7008 VSS.n9901 VSS.n9900 0.0525625
R7009 VSS.n7754 VSS.n6263 0.0525625
R7010 VSS.n8964 VSS.n6258 0.0525625
R7011 VSS.n9864 VSS.n7146 0.0525625
R7012 VSS.n9847 VSS.n9846 0.0525625
R7013 VSS.n9525 VSS.n9524 0.0525625
R7014 VSS.n9807 VSS.n9794 0.0525625
R7015 VSS.n9466 VSS.n9453 0.0525625
R7016 VSS.n9610 VSS.n9609 0.0525625
R7017 VSS.n8769 VSS.n8756 0.0525625
R7018 VSS.n1367 VSS.n1354 0.0525625
R7019 VSS.n14153 VSS.n14152 0.0525625
R7020 VSS.n14375 VSS 0.0524238
R7021 VSS.n980 VSS 0.0524238
R7022 VSS.n700 VSS 0.0524238
R7023 VSS.n11143 VSS.n3713 0.0520625
R7024 VSS.n13373 VSS.n13371 0.0515417
R7025 VSS.n13838 VSS.n13836 0.0515417
R7026 VSS.n1598 VSS.n1596 0.0515417
R7027 VSS.n12042 VSS.n11781 0.0515417
R7028 VSS.n10639 VSS.n10638 0.0513775
R7029 VSS.n12334 VSS.n11547 0.0513775
R7030 VSS.n14461 VSS.n23 0.05126
R7031 VSS.n3344 VSS.n3343 0.05126
R7032 VSS.n11907 VSS.n11906 0.05126
R7033 VSS.n11763 VSS.n11762 0.05126
R7034 VSS.n3619 VSS.n3618 0.05126
R7035 VSS.n4486 VSS.n4484 0.05126
R7036 VSS.n1054 VSS.n476 0.05126
R7037 VSS.n13816 VSS.n485 0.05126
R7038 VSS.n13353 VSS.n490 0.05126
R7039 VSS.n14381 VSS.n487 0.05126
R7040 VSS.n1576 VSS.n481 0.05126
R7041 VSS.n453 VSS.n449 0.05126
R7042 VSS.n1304 VSS.n446 0.05126
R7043 VSS.n14340 VSS.n494 0.05126
R7044 VSS.n14380 VSS.n14378 0.05126
R7045 VSS.n14381 VSS.n498 0.05126
R7046 VSS.n11538 VSS.n11537 0.05126
R7047 VSS.n11789 VSS.n11788 0.05126
R7048 VSS.n3422 VSS.n3421 0.05126
R7049 VSS.n14511 VSS.n14510 0.051025
R7050 VSS.n12327 VSS.n12326 0.050555
R7051 VSS.n3331 VSS.n3330 0.0505002
R7052 VSS.n9771 VSS.n9770 0.0499792
R7053 VSS.n10786 VSS.n10784 0.0494583
R7054 VSS.n11291 VSS.n11290 0.0489848
R7055 VSS.n11293 VSS.n11292 0.0489848
R7056 VSS.n14362 VSS.n14360 0.0489375
R7057 VSS.n11079 VSS 0.0487365
R7058 VSS.n11566 VSS.n11565 0.047735
R7059 VSS.n3614 VSS 0.0475
R7060 VSS.n292 VSS 0.0475
R7061 VSS.n4531 VSS 0.0475
R7062 VSS.n4505 VSS 0.0475
R7063 VSS.n4458 VSS 0.0475
R7064 VSS.n4491 VSS 0.0475
R7065 VSS.n4469 VSS 0.0475
R7066 VSS.n4482 VSS 0.0475
R7067 VSS.n373 VSS 0.0475
R7068 VSS.n171 VSS 0.0475
R7069 VSS.n28 VSS 0.0475
R7070 VSS.n335 VSS 0.0475
R7071 VSS.n262 VSS 0.0475
R7072 VSS.n150 VSS 0.0475
R7073 VSS.n89 VSS 0.0475
R7074 VSS.n2 VSS 0.0475
R7075 VSS.n11532 VSS.n11525 0.047265
R7076 VSS.n3570 VSS.n3569 0.0469125
R7077 VSS.n14370 VSS.n14368 0.0468542
R7078 VSS.n1314 VSS.n1312 0.046795
R7079 VSS.n11150 VSS.n11149 0.0464425
R7080 VSS.n9426 VSS.n9424 0.0463333
R7081 VSS.n12281 VSS.n12280 0.046325
R7082 VSS.n12038 VSS.n12031 0.046325
R7083 VSS.n1063 VSS.n1062 0.0452675
R7084 VSS.n5788 VSS.n5786 0.0447708
R7085 VSS.n3363 VSS.n3362 0.04468
R7086 VSS.n1312 VSS 0.0445116
R7087 VSS.n1062 VSS 0.0444436
R7088 VSS.n14348 VSS 0.0443757
R7089 VSS.n13824 VSS 0.0443757
R7090 VSS.n13361 VSS 0.0443757
R7091 VSS.n1584 VSS 0.0443757
R7092 VSS.n469 VSS 0.0443757
R7093 VSS.n691 VSS.n690 0.0442502
R7094 VSS.n3342 VSS 0.0439131
R7095 VSS.n3420 VSS 0.0439131
R7096 VSS.n11903 VSS 0.0439131
R7097 VSS.n11787 VSS 0.0439131
R7098 VSS.n11759 VSS 0.0439131
R7099 VSS.n11536 VSS 0.0439131
R7100 VSS.n3615 VSS 0.0439131
R7101 VSS.n480 VSS 0.0439131
R7102 VSS.n291 VSS 0.0439131
R7103 VSS.n493 VSS 0.0439131
R7104 VSS.n4517 VSS 0.0439131
R7105 VSS.n4457 VSS 0.0439131
R7106 VSS.n4468 VSS 0.0439131
R7107 VSS.n4479 VSS 0.0439131
R7108 VSS.n4485 VSS 0.0439131
R7109 VSS.n4489 VSS 0.0439131
R7110 VSS.n4503 VSS 0.0439131
R7111 VSS.n475 VSS 0.0439131
R7112 VSS.n484 VSS 0.0439131
R7113 VSS.n488 VSS 0.0439131
R7114 VSS.n489 VSS 0.0439131
R7115 VSS.n372 VSS 0.0439131
R7116 VSS.n14457 VSS 0.0439131
R7117 VSS.n14454 VSS 0.0439131
R7118 VSS.n448 VSS 0.0439131
R7119 VSS.n445 VSS 0.0439131
R7120 VSS.n499 VSS 0.0439131
R7121 VSS.n14379 VSS 0.0439131
R7122 VSS.n348 VSS 0.0439131
R7123 VSS.n275 VSS 0.0439131
R7124 VSS.n165 VSS 0.0439131
R7125 VSS.n38 VSS 0.0439131
R7126 VSS.n6152 VSS.n6150 0.0437292
R7127 VSS.n5969 VSS.n5967 0.0437292
R7128 VSS.n4526 VSS 0.0437243
R7129 VSS.n1585 VSS.n1584 0.0436225
R7130 VSS.n13825 VSS.n13824 0.0436225
R7131 VSS.n13365 VSS.n13361 0.0436225
R7132 VSS.n469 VSS.n468 0.0436225
R7133 VSS.n10107 VSS.n10106 0.043505
R7134 VSS.n12202 VSS.n12201 0.043505
R7135 VSS.n14354 VSS.n14348 0.043035
R7136 VSS.n5597 VSS.n5595 0.042095
R7137 VSS.n12574 VSS.n12570 0.0415075
R7138 VSS.n12166 VSS.n12165 0.04139
R7139 VSS.n12468 VSS.n12467 0.0405675
R7140 VSS.n13417 VSS.n490 0.0400873
R7141 VSS.n9116 VSS.n9055 0.0400833
R7142 VSS.n5564 VSS.n5563 0.0396275
R7143 VSS.n10100 VSS.n4571 0.0390417
R7144 VSS.n12206 VSS.n11752 0.0390417
R7145 VSS.n4490 VSS.n4488 0.03904
R7146 VSS.n4504 VSS.n4502 0.03904
R7147 VSS.n4518 VSS.n4516 0.03904
R7148 VSS.n3914 VSS.n3913 0.0389306
R7149 VSS.n13616 VSS.n13615 0.0389306
R7150 VSS.n4488 VSS.n4481 0.0383507
R7151 VSS.n13421 VSS.n13420 0.038335
R7152 VSS.n13420 VSS.n13419 0.038221
R7153 VSS.n9946 VSS.n9945 0.0381806
R7154 VSS.n8838 VSS.n8837 0.0381806
R7155 VSS.n8841 VSS.n7593 0.0381806
R7156 VSS.n9603 VSS.n9602 0.0381806
R7157 VSS.n8759 VSS.n8758 0.0381806
R7158 VSS.n8517 VSS.n8516 0.0381806
R7159 VSS.n9799 VSS.n9798 0.0381806
R7160 VSS.n9456 VSS.n9455 0.0381806
R7161 VSS.n9147 VSS.n9146 0.0381806
R7162 VSS.n7603 VSS.n7152 0.0381806
R7163 VSS.n9855 VSS.n9854 0.0381806
R7164 VSS.n9529 VSS.n9528 0.0381806
R7165 VSS.n9539 VSS.n9538 0.0381806
R7166 VSS.n9910 VSS.n9909 0.0381806
R7167 VSS.n9918 VSS.n9917 0.0381806
R7168 VSS.n9926 VSS.n9925 0.0381806
R7169 VSS.n9934 VSS.n9933 0.0381806
R7170 VSS.n9940 VSS.n9939 0.0381806
R7171 VSS.n10032 VSS.n10031 0.0381806
R7172 VSS.n10025 VSS.n10024 0.0381806
R7173 VSS.n10016 VSS.n10015 0.0381806
R7174 VSS.n10007 VSS.n10006 0.0381806
R7175 VSS.n9998 VSS.n9997 0.0381806
R7176 VSS.n9989 VSS.n9988 0.0381806
R7177 VSS.n10035 VSS.n3818 0.0381806
R7178 VSS.n9905 VSS.n3847 0.0381806
R7179 VSS.n9858 VSS.n3886 0.0381806
R7180 VSS.n14244 VSS.n14243 0.0381806
R7181 VSS.n13064 VSS.n1905 0.0381806
R7182 VSS.n2425 VSS.n611 0.0381806
R7183 VSS.n14146 VSS.n14145 0.0381806
R7184 VSS.n1359 VSS.n1358 0.0381806
R7185 VSS.n1118 VSS.n1117 0.0381806
R7186 VSS.n13867 VSS.n13866 0.0381806
R7187 VSS.n1634 VSS.n1633 0.0381806
R7188 VSS.n800 VSS.n799 0.0381806
R7189 VSS.n14051 VSS.n14050 0.0381806
R7190 VSS.n14043 VSS.n14042 0.0381806
R7191 VSS.n14128 VSS.n14127 0.0381806
R7192 VSS.n14138 VSS.n14137 0.0381806
R7193 VSS.n12699 VSS.n1886 0.0381806
R7194 VSS.n13174 VSS.n13173 0.0381806
R7195 VSS.n13167 VSS.n13166 0.0381806
R7196 VSS.n13158 VSS.n13157 0.0381806
R7197 VSS.n13149 VSS.n13148 0.0381806
R7198 VSS.n12844 VSS.n12843 0.0381806
R7199 VSS.n2914 VSS.n2913 0.0381806
R7200 VSS.n12921 VSS.n12920 0.0381806
R7201 VSS.n2734 VSS.n2733 0.0381806
R7202 VSS.n12998 VSS.n12997 0.0381806
R7203 VSS.n12427 VSS.n12426 0.0381806
R7204 VSS.n12839 VSS.n12838 0.0381806
R7205 VSS.n12702 VSS.n1753 0.0381806
R7206 VSS.n14038 VSS.n14037 0.0381806
R7207 VSS.n3440 VSS.n3417 0.0381
R7208 VSS.n5237 VSS.n5235 0.0379825
R7209 VSS.n11999 VSS.n11998 0.037395
R7210 VSS.n5384 VSS.n5383 0.0370425
R7211 VSS.n3308 VSS.n3307 0.0370425
R7212 VSS.n14505 VSS.n14504 0.0370425
R7213 VSS VSS 0.0369583
R7214 VSS.n11925 VSS.n11902 0.03669
R7215 VSS.n5744 VSS.n5743 0.0365725
R7216 VSS.n27 VSS.n25 0.03622
R7217 VSS.n3613 VSS.n47 0.0361104
R7218 VSS.n5417 VSS.n5415 0.0361025
R7219 VSS.n6210 VSS.n4659 0.0356744
R7220 VSS.n9949 VSS.n6234 0.0356744
R7221 VSS.n8159 VSS.n8013 0.0356744
R7222 VSS.n4275 VSS.n4204 0.0356744
R7223 VSS.n4160 VSS.n4158 0.0356744
R7224 VSS.n12430 VSS.n12395 0.0356744
R7225 VSS.n13061 VSS.n2459 0.0356744
R7226 VSS.n2428 VSS.n2395 0.0356744
R7227 VSS.n10152 VSS.n10151 0.0351625
R7228 VSS.n9985 VSS.n4659 0.035093
R7229 VSS.n8123 VSS.n6234 0.035093
R7230 VSS.n8834 VSS.n8013 0.035093
R7231 VSS.n4358 VSS.n4204 0.035093
R7232 VSS.n4435 VSS.n4158 0.035093
R7233 VSS.n12422 VSS.n12395 0.035093
R7234 VSS.n13067 VSS.n2459 0.035093
R7235 VSS.n2422 VSS.n2395 0.035093
R7236 VSS.n11797 VSS.n11796 0.0348752
R7237 VSS.n3646 VSS 0.0343542
R7238 VSS.n11212 VSS 0.0343542
R7239 VSS.n8490 VSS.n8411 0.0341111
R7240 VSS.n4659 VSS.n4658 0.0341111
R7241 VSS.n9947 VSS.n6234 0.0341111
R7242 VSS.n9942 VSS.n9941 0.0341111
R7243 VSS.n8013 VSS.n8012 0.0341111
R7244 VSS.n8842 VSS.n8010 0.0341111
R7245 VSS.n7595 VSS.n7592 0.0341111
R7246 VSS.n9607 VSS.n9606 0.0341111
R7247 VSS.n8767 VSS.n8766 0.0341111
R7248 VSS.n8524 VSS.n8523 0.0341111
R7249 VSS.n9805 VSS.n9804 0.0341111
R7250 VSS.n9464 VSS.n9463 0.0341111
R7251 VSS.n9155 VSS.n9154 0.0341111
R7252 VSS.n9860 VSS.n7149 0.0341111
R7253 VSS.n7151 VSS.n7150 0.0341111
R7254 VSS.n7607 VSS.n7606 0.0341111
R7255 VSS.n9534 VSS.n9533 0.0341111
R7256 VSS.n9907 VSS.n9903 0.0341111
R7257 VSS.n9914 VSS.n9913 0.0341111
R7258 VSS.n9922 VSS.n9921 0.0341111
R7259 VSS.n9930 VSS.n9929 0.0341111
R7260 VSS.n9936 VSS.n9935 0.0341111
R7261 VSS.n10037 VSS.n4635 0.0341111
R7262 VSS.n10029 VSS.n4636 0.0341111
R7263 VSS.n10020 VSS.n4642 0.0341111
R7264 VSS.n10011 VSS.n4646 0.0341111
R7265 VSS.n10002 VSS.n4650 0.0341111
R7266 VSS.n9993 VSS.n4654 0.0341111
R7267 VSS.n3820 VSS.n3817 0.0341111
R7268 VSS.n3846 VSS.n3845 0.0341111
R7269 VSS.n3888 VSS.n3885 0.0341111
R7270 VSS.n3912 VSS.n3911 0.0341111
R7271 VSS.n4205 VSS.n4204 0.0341111
R7272 VSS.n4158 VSS.n4157 0.0341111
R7273 VSS.n14238 VSS.n542 0.0341111
R7274 VSS.n14246 VSS.n541 0.0341111
R7275 VSS.n12428 VSS.n12395 0.0341111
R7276 VSS.n13063 VSS.n2459 0.0341111
R7277 VSS.n1904 VSS.n1902 0.0341111
R7278 VSS.n2426 VSS.n2395 0.0341111
R7279 VSS.n14147 VSS.n610 0.0341111
R7280 VSS.n14142 VSS.n14141 0.0341111
R7281 VSS.n1365 VSS.n1364 0.0341111
R7282 VSS.n1126 VSS.n1125 0.0341111
R7283 VSS.n13873 VSS.n13872 0.0341111
R7284 VSS.n1628 VSS.n1627 0.0341111
R7285 VSS.n808 VSS.n807 0.0341111
R7286 VSS.n14040 VSS.n1706 0.0341111
R7287 VSS.n14055 VSS.n14054 0.0341111
R7288 VSS.n14048 VSS.n14045 0.0341111
R7289 VSS.n14133 VSS.n14132 0.0341111
R7290 VSS.n12704 VSS.n12698 0.0341111
R7291 VSS.n13178 VSS.n13177 0.0341111
R7292 VSS.n13171 VSS.n1888 0.0341111
R7293 VSS.n13162 VSS.n1894 0.0341111
R7294 VSS.n13153 VSS.n1898 0.0341111
R7295 VSS.n12841 VSS.n2921 0.0341111
R7296 VSS.n2916 VSS.n2907 0.0341111
R7297 VSS.n2909 VSS.n2908 0.0341111
R7298 VSS.n2736 VSS.n2727 0.0341111
R7299 VSS.n2729 VSS.n2728 0.0341111
R7300 VSS.n13000 VSS.n12999 0.0341111
R7301 VSS.n12834 VSS.n12833 0.0341111
R7302 VSS.n1752 VSS.n1751 0.0341111
R7303 VSS.n14033 VSS.n14032 0.0341111
R7304 VSS.n13624 VSS.n13623 0.0341111
R7305 VSS.n5204 VSS.n5203 0.034105
R7306 VSS.n8515 VSS.n8411 0.0335556
R7307 VSS.n9987 VSS.n4659 0.0335556
R7308 VSS.n6235 VSS.n6234 0.0335556
R7309 VSS.n9942 VSS.n6240 0.0335556
R7310 VSS.n8836 VSS.n8013 0.0335556
R7311 VSS.n8839 VSS.n8010 0.0335556
R7312 VSS.n9541 VSS.n7592 0.0335556
R7313 VSS.n9607 VSS.n9601 0.0335556
R7314 VSS.n8767 VSS.n8764 0.0335556
R7315 VSS.n8524 VSS.n8521 0.0335556
R7316 VSS.n9805 VSS.n9797 0.0335556
R7317 VSS.n9464 VSS.n9461 0.0335556
R7318 VSS.n9155 VSS.n9152 0.0335556
R7319 VSS.n9857 VSS.n7149 0.0335556
R7320 VSS.n9853 VSS.n7151 0.0335556
R7321 VSS.n7607 VSS.n7602 0.0335556
R7322 VSS.n9534 VSS.n7598 0.0335556
R7323 VSS.n9904 VSS.n9903 0.0335556
R7324 VSS.n9914 VSS.n6264 0.0335556
R7325 VSS.n9922 VSS.n6259 0.0335556
R7326 VSS.n9930 VSS.n6254 0.0335556
R7327 VSS.n9936 VSS.n6247 0.0335556
R7328 VSS.n10034 VSS.n4635 0.0335556
R7329 VSS.n10030 VSS.n10029 0.0335556
R7330 VSS.n10023 VSS.n10020 0.0335556
R7331 VSS.n10014 VSS.n10011 0.0335556
R7332 VSS.n10005 VSS.n10002 0.0335556
R7333 VSS.n9996 VSS.n9993 0.0335556
R7334 VSS.n11120 VSS.n3817 0.0335556
R7335 VSS.n11002 VSS.n3846 0.0335556
R7336 VSS.n10961 VSS.n3885 0.0335556
R7337 VSS.n10848 VSS.n3912 0.0335556
R7338 VSS.n4356 VSS.n4204 0.0335556
R7339 VSS.n4437 VSS.n4158 0.0335556
R7340 VSS.n14242 VSS.n542 0.0335556
R7341 VSS.n541 VSS.n540 0.0335556
R7342 VSS.n12424 VSS.n12395 0.0335556
R7343 VSS.n13065 VSS.n2459 0.0335556
R7344 VSS.n13147 VSS.n1904 0.0335556
R7345 VSS.n2424 VSS.n2395 0.0335556
R7346 VSS.n612 VSS.n610 0.0335556
R7347 VSS.n14142 VSS.n618 0.0335556
R7348 VSS.n1365 VSS.n1357 0.0335556
R7349 VSS.n1126 VSS.n1123 0.0335556
R7350 VSS.n13873 VSS.n13865 0.0335556
R7351 VSS.n1630 VSS.n1628 0.0335556
R7352 VSS.n808 VSS.n805 0.0335556
R7353 VSS.n1707 VSS.n1706 0.0335556
R7354 VSS.n14055 VSS.n1701 0.0335556
R7355 VSS.n14049 VSS.n14048 0.0335556
R7356 VSS.n14133 VSS.n621 0.0335556
R7357 VSS.n12701 VSS.n12698 0.0335556
R7358 VSS.n13178 VSS.n1885 0.0335556
R7359 VSS.n13172 VSS.n13171 0.0335556
R7360 VSS.n13165 VSS.n13162 0.0335556
R7361 VSS.n13156 VSS.n13153 0.0335556
R7362 VSS.n2922 VSS.n2921 0.0335556
R7363 VSS.n12846 VSS.n2907 0.0335556
R7364 VSS.n2912 VSS.n2909 0.0335556
R7365 VSS.n12923 VSS.n2727 0.0335556
R7366 VSS.n2732 VSS.n2729 0.0335556
R7367 VSS.n13000 VSS.n2553 0.0335556
R7368 VSS.n12834 VSS.n2925 0.0335556
R7369 VSS.n13998 VSS.n1752 0.0335556
R7370 VSS.n14033 VSS.n1710 0.0335556
R7371 VSS.n13624 VSS.n13621 0.0335556
R7372 VSS.n11354 VSS 0.0330521
R7373 VSS.n11344 VSS 0.0330521
R7374 VSS VSS.n11487 0.0330521
R7375 VSS VSS.n11276 0.0330521
R7376 VSS.n5605 VSS.n4691 0.0327917
R7377 VSS.n6142 VSS.n6138 0.032695
R7378 VSS.n5959 VSS.n5956 0.032695
R7379 VSS.n5778 VSS.n5775 0.03246
R7380 VSS.n5187 VSS.n5186 0.0322708
R7381 VSS.n11525 VSS.n11524 0.031755
R7382 VSS.n8763 VSS 0.03175
R7383 VSS VSS.n8760 0.03175
R7384 VSS VSS.n8761 0.03175
R7385 VSS.n8761 VSS 0.03175
R7386 VSS.n6241 VSS 0.03175
R7387 VSS VSS.n6238 0.03175
R7388 VSS VSS.n9944 0.03175
R7389 VSS.n9944 VSS 0.03175
R7390 VSS.n8840 VSS 0.03175
R7391 VSS VSS.n8011 0.03175
R7392 VSS.n8845 VSS 0.03175
R7393 VSS.n8845 VSS 0.03175
R7394 VSS.n9540 VSS 0.03175
R7395 VSS VSS.n7589 0.03175
R7396 VSS.n9543 VSS 0.03175
R7397 VSS.n9543 VSS 0.03175
R7398 VSS VSS.n7548 0.03175
R7399 VSS VSS.n9599 0.03175
R7400 VSS.n9599 VSS 0.03175
R7401 VSS.n9605 VSS 0.03175
R7402 VSS.n8520 VSS 0.03175
R7403 VSS VSS.n8364 0.03175
R7404 VSS VSS.n8518 0.03175
R7405 VSS.n8518 VSS 0.03175
R7406 VSS.n9460 VSS 0.03175
R7407 VSS VSS.n9457 0.03175
R7408 VSS VSS.n9458 0.03175
R7409 VSS.n9458 VSS 0.03175
R7410 VSS VSS.n9800 0.03175
R7411 VSS VSS.n9801 0.03175
R7412 VSS.n9801 VSS 0.03175
R7413 VSS.n9803 VSS 0.03175
R7414 VSS.n9151 VSS 0.03175
R7415 VSS VSS.n9148 0.03175
R7416 VSS VSS.n9149 0.03175
R7417 VSS.n9149 VSS 0.03175
R7418 VSS.n7605 VSS 0.03175
R7419 VSS VSS.n7601 0.03175
R7420 VSS VSS.n9527 0.03175
R7421 VSS.n9527 VSS 0.03175
R7422 VSS.n9852 VSS 0.03175
R7423 VSS VSS.n7153 0.03175
R7424 VSS VSS.n9849 0.03175
R7425 VSS.n9849 VSS 0.03175
R7426 VSS.n9862 VSS 0.03175
R7427 VSS VSS.n7148 0.03175
R7428 VSS.n7148 VSS 0.03175
R7429 VSS.n9859 VSS 0.03175
R7430 VSS.n9531 VSS 0.03175
R7431 VSS.n7596 VSS 0.03175
R7432 VSS.n9536 VSS 0.03175
R7433 VSS.n9536 VSS 0.03175
R7434 VSS.n9928 VSS 0.03175
R7435 VSS VSS.n6252 0.03175
R7436 VSS VSS.n9932 0.03175
R7437 VSS.n9932 VSS 0.03175
R7438 VSS.n9919 VSS 0.03175
R7439 VSS VSS.n6257 0.03175
R7440 VSS VSS.n9924 0.03175
R7441 VSS.n9924 VSS 0.03175
R7442 VSS.n9911 VSS 0.03175
R7443 VSS VSS.n6262 0.03175
R7444 VSS VSS.n9916 0.03175
R7445 VSS.n9916 VSS 0.03175
R7446 VSS VSS.n6266 0.03175
R7447 VSS VSS.n6267 0.03175
R7448 VSS VSS.n6267 0.03175
R7449 VSS.n9906 VSS 0.03175
R7450 VSS.n6248 VSS 0.03175
R7451 VSS VSS.n6245 0.03175
R7452 VSS VSS.n9938 0.03175
R7453 VSS.n9938 VSS 0.03175
R7454 VSS.n10004 VSS 0.03175
R7455 VSS VSS.n4653 0.03175
R7456 VSS.n10000 VSS 0.03175
R7457 VSS.n10000 VSS 0.03175
R7458 VSS.n10013 VSS 0.03175
R7459 VSS VSS.n4649 0.03175
R7460 VSS.n10009 VSS 0.03175
R7461 VSS.n10009 VSS 0.03175
R7462 VSS.n10022 VSS 0.03175
R7463 VSS VSS.n4645 0.03175
R7464 VSS.n10018 VSS 0.03175
R7465 VSS.n10018 VSS 0.03175
R7466 VSS.n4637 VSS 0.03175
R7467 VSS VSS.n4640 0.03175
R7468 VSS.n10027 VSS 0.03175
R7469 VSS.n10027 VSS 0.03175
R7470 VSS.n10039 VSS 0.03175
R7471 VSS VSS.n4634 0.03175
R7472 VSS.n4634 VSS 0.03175
R7473 VSS.n10036 VSS 0.03175
R7474 VSS.n9995 VSS 0.03175
R7475 VSS VSS.n4657 0.03175
R7476 VSS.n9991 VSS 0.03175
R7477 VSS.n9991 VSS 0.03175
R7478 VSS.n11119 VSS 0.03175
R7479 VSS.n11122 VSS 0.03175
R7480 VSS VSS.n3816 0.03175
R7481 VSS.n3816 VSS 0.03175
R7482 VSS.n11001 VSS 0.03175
R7483 VSS VSS.n3848 0.03175
R7484 VSS VSS.n10998 0.03175
R7485 VSS.n10998 VSS 0.03175
R7486 VSS.n10960 VSS 0.03175
R7487 VSS.n10963 VSS 0.03175
R7488 VSS VSS.n3884 0.03175
R7489 VSS.n3884 VSS 0.03175
R7490 VSS.n10847 VSS 0.03175
R7491 VSS VSS.n3915 0.03175
R7492 VSS VSS.n10845 0.03175
R7493 VSS.n10845 VSS 0.03175
R7494 VSS.n14245 VSS 0.03175
R7495 VSS VSS.n536 0.03175
R7496 VSS.n14248 VSS 0.03175
R7497 VSS.n14248 VSS 0.03175
R7498 VSS.n1903 VSS 0.03175
R7499 VSS VSS.n1906 0.03175
R7500 VSS VSS.n13144 0.03175
R7501 VSS.n13144 VSS 0.03175
R7502 VSS.n613 VSS 0.03175
R7503 VSS VSS.n607 0.03175
R7504 VSS.n14150 VSS 0.03175
R7505 VSS.n14150 VSS 0.03175
R7506 VSS.n14140 VSS 0.03175
R7507 VSS VSS.n616 0.03175
R7508 VSS VSS.n14144 0.03175
R7509 VSS.n14144 VSS 0.03175
R7510 VSS VSS.n1360 0.03175
R7511 VSS VSS.n1361 0.03175
R7512 VSS.n1361 VSS 0.03175
R7513 VSS.n1363 VSS 0.03175
R7514 VSS.n1122 VSS 0.03175
R7515 VSS VSS.n1119 0.03175
R7516 VSS VSS.n1120 0.03175
R7517 VSS.n1120 VSS 0.03175
R7518 VSS.n1629 VSS 0.03175
R7519 VSS.n1636 VSS 0.03175
R7520 VSS VSS.n1632 0.03175
R7521 VSS.n1632 VSS 0.03175
R7522 VSS VSS.n13868 0.03175
R7523 VSS VSS.n13869 0.03175
R7524 VSS.n13869 VSS 0.03175
R7525 VSS.n13871 VSS 0.03175
R7526 VSS.n804 VSS 0.03175
R7527 VSS VSS.n801 0.03175
R7528 VSS VSS.n802 0.03175
R7529 VSS.n802 VSS 0.03175
R7530 VSS.n14046 VSS 0.03175
R7531 VSS VSS.n624 0.03175
R7532 VSS VSS.n14126 0.03175
R7533 VSS.n14126 VSS 0.03175
R7534 VSS.n14044 VSS 0.03175
R7535 VSS VSS.n1697 0.03175
R7536 VSS VSS.n1700 0.03175
R7537 VSS.n1700 VSS 0.03175
R7538 VSS VSS.n1703 0.03175
R7539 VSS VSS.n1704 0.03175
R7540 VSS VSS.n1704 0.03175
R7541 VSS.n14039 VSS 0.03175
R7542 VSS.n14130 VSS 0.03175
R7543 VSS.n619 VSS 0.03175
R7544 VSS.n14135 VSS 0.03175
R7545 VSS.n14135 VSS 0.03175
R7546 VSS.n13164 VSS 0.03175
R7547 VSS VSS.n1897 0.03175
R7548 VSS.n13160 VSS 0.03175
R7549 VSS.n13160 VSS 0.03175
R7550 VSS.n1889 VSS 0.03175
R7551 VSS VSS.n1892 0.03175
R7552 VSS.n13169 VSS 0.03175
R7553 VSS.n13169 VSS 0.03175
R7554 VSS.n1887 VSS 0.03175
R7555 VSS VSS.n1881 0.03175
R7556 VSS VSS.n1884 0.03175
R7557 VSS.n1884 VSS 0.03175
R7558 VSS.n12706 VSS 0.03175
R7559 VSS VSS.n12697 0.03175
R7560 VSS.n12697 VSS 0.03175
R7561 VSS.n12703 VSS 0.03175
R7562 VSS.n13155 VSS 0.03175
R7563 VSS VSS.n1901 0.03175
R7564 VSS.n13151 VSS 0.03175
R7565 VSS.n13151 VSS 0.03175
R7566 VSS.n2731 VSS 0.03175
R7567 VSS VSS.n2558 0.03175
R7568 VSS VSS.n12996 0.03175
R7569 VSS.n12996 VSS 0.03175
R7570 VSS.n12922 VSS 0.03175
R7571 VSS VSS.n2724 0.03175
R7572 VSS.n12925 VSS 0.03175
R7573 VSS.n12925 VSS 0.03175
R7574 VSS.n2911 VSS 0.03175
R7575 VSS VSS.n2739 0.03175
R7576 VSS VSS.n12919 0.03175
R7577 VSS.n12919 VSS 0.03175
R7578 VSS.n12845 VSS 0.03175
R7579 VSS VSS.n2904 0.03175
R7580 VSS.n12848 VSS 0.03175
R7581 VSS.n12848 VSS 0.03175
R7582 VSS VSS.n2918 0.03175
R7583 VSS VSS.n2919 0.03175
R7584 VSS VSS.n2919 0.03175
R7585 VSS.n12840 VSS 0.03175
R7586 VSS.n2554 VSS 0.03175
R7587 VSS VSS.n2549 0.03175
R7588 VSS VSS.n2552 0.03175
R7589 VSS.n2552 VSS 0.03175
R7590 VSS.n12830 VSS 0.03175
R7591 VSS.n2924 VSS 0.03175
R7592 VSS.n12836 VSS 0.03175
R7593 VSS.n12836 VSS 0.03175
R7594 VSS.n13997 VSS 0.03175
R7595 VSS VSS.n1754 0.03175
R7596 VSS VSS.n13994 0.03175
R7597 VSS.n13994 VSS 0.03175
R7598 VSS.n14029 VSS 0.03175
R7599 VSS.n1709 VSS 0.03175
R7600 VSS.n14035 VSS 0.03175
R7601 VSS.n14035 VSS 0.03175
R7602 VSS.n13620 VSS 0.03175
R7603 VSS VSS.n13617 0.03175
R7604 VSS VSS.n13618 0.03175
R7605 VSS.n13618 VSS 0.03175
R7606 VSS.n6239 VSS.n6236 0.0316203
R7607 VSS.n9943 VSS.n6239 0.0316203
R7608 VSS.n8847 VSS.n8009 0.0316203
R7609 VSS.n8847 VSS.n8846 0.0316203
R7610 VSS.n9545 VSS.n7591 0.0316203
R7611 VSS.n9545 VSS.n9544 0.0316203
R7612 VSS.n9609 VSS.n9598 0.0316203
R7613 VSS.n9609 VSS.n9608 0.0316203
R7614 VSS.n8769 VSS.n8757 0.0316203
R7615 VSS.n8769 VSS.n8768 0.0316203
R7616 VSS.n8526 VSS.n8410 0.0316203
R7617 VSS.n8526 VSS.n8525 0.0316203
R7618 VSS.n9807 VSS.n9795 0.0316203
R7619 VSS.n9807 VSS.n9806 0.0316203
R7620 VSS.n9466 VSS.n9454 0.0316203
R7621 VSS.n9466 VSS.n9465 0.0316203
R7622 VSS.n9157 VSS.n9145 0.0316203
R7623 VSS.n9157 VSS.n9156 0.0316203
R7624 VSS.n9864 VSS.n7147 0.0316203
R7625 VSS.n9864 VSS.n9863 0.0316203
R7626 VSS.n9847 VSS.n7154 0.0316203
R7627 VSS.n9848 VSS.n9847 0.0316203
R7628 VSS.n9525 VSS.n7599 0.0316203
R7629 VSS.n9525 VSS.n7608 0.0316203
R7630 VSS.n9537 VSS.n7597 0.0316203
R7631 VSS.n9535 VSS.n7597 0.0316203
R7632 VSS.n9901 VSS.n6265 0.0316203
R7633 VSS.n9902 VSS.n9901 0.0316203
R7634 VSS.n6263 VSS.n6260 0.0316203
R7635 VSS.n9915 VSS.n6263 0.0316203
R7636 VSS.n6258 VSS.n6255 0.0316203
R7637 VSS.n9923 VSS.n6258 0.0316203
R7638 VSS.n6253 VSS.n6250 0.0316203
R7639 VSS.n9931 VSS.n6253 0.0316203
R7640 VSS.n6246 VSS.n6243 0.0316203
R7641 VSS.n9937 VSS.n6246 0.0316203
R7642 VSS.n10041 VSS.n4633 0.0316203
R7643 VSS.n10041 VSS.n10040 0.0316203
R7644 VSS.n10026 VSS.n4639 0.0316203
R7645 VSS.n10028 VSS.n4639 0.0316203
R7646 VSS.n10017 VSS.n4644 0.0316203
R7647 VSS.n10019 VSS.n4644 0.0316203
R7648 VSS.n10008 VSS.n4648 0.0316203
R7649 VSS.n10010 VSS.n4648 0.0316203
R7650 VSS.n9999 VSS.n4652 0.0316203
R7651 VSS.n10001 VSS.n4652 0.0316203
R7652 VSS.n9990 VSS.n4656 0.0316203
R7653 VSS.n9992 VSS.n4656 0.0316203
R7654 VSS.n11124 VSS.n3815 0.0316203
R7655 VSS.n11124 VSS.n11123 0.0316203
R7656 VSS.n10996 VSS.n3849 0.0316203
R7657 VSS.n10997 VSS.n10996 0.0316203
R7658 VSS.n10965 VSS.n3883 0.0316203
R7659 VSS.n10965 VSS.n10964 0.0316203
R7660 VSS.n10844 VSS.n10843 0.0316203
R7661 VSS.n10843 VSS.n10842 0.0316203
R7662 VSS.n14250 VSS.n538 0.0316203
R7663 VSS.n14250 VSS.n14249 0.0316203
R7664 VSS.n13142 VSS.n1907 0.0316203
R7665 VSS.n13143 VSS.n13142 0.0316203
R7666 VSS.n14152 VSS.n609 0.0316203
R7667 VSS.n14152 VSS.n14151 0.0316203
R7668 VSS.n617 VSS.n614 0.0316203
R7669 VSS.n14143 VSS.n617 0.0316203
R7670 VSS.n1367 VSS.n1355 0.0316203
R7671 VSS.n1367 VSS.n1366 0.0316203
R7672 VSS.n1128 VSS.n1116 0.0316203
R7673 VSS.n1128 VSS.n1127 0.0316203
R7674 VSS.n13875 VSS.n13863 0.0316203
R7675 VSS.n13875 VSS.n13874 0.0316203
R7676 VSS.n810 VSS.n798 0.0316203
R7677 VSS.n810 VSS.n809 0.0316203
R7678 VSS.n13913 VSS.n1702 0.0316203
R7679 VSS.n13913 VSS.n13912 0.0316203
R7680 VSS.n14057 VSS.n1699 0.0316203
R7681 VSS.n14057 VSS.n14056 0.0316203
R7682 VSS.n14124 VSS.n622 0.0316203
R7683 VSS.n14124 VSS.n625 0.0316203
R7684 VSS.n14136 VSS.n620 0.0316203
R7685 VSS.n14134 VSS.n620 0.0316203
R7686 VSS.n12708 VSS.n12696 0.0316203
R7687 VSS.n12708 VSS.n12707 0.0316203
R7688 VSS.n13180 VSS.n1883 0.0316203
R7689 VSS.n13180 VSS.n13179 0.0316203
R7690 VSS.n13168 VSS.n1891 0.0316203
R7691 VSS.n13170 VSS.n1891 0.0316203
R7692 VSS.n13159 VSS.n1896 0.0316203
R7693 VSS.n13161 VSS.n1896 0.0316203
R7694 VSS.n13150 VSS.n1900 0.0316203
R7695 VSS.n13152 VSS.n1900 0.0316203
R7696 VSS.n12613 VSS.n2917 0.0316203
R7697 VSS.n12613 VSS.n12612 0.0316203
R7698 VSS.n12850 VSS.n2906 0.0316203
R7699 VSS.n12850 VSS.n12849 0.0316203
R7700 VSS.n12917 VSS.n2737 0.0316203
R7701 VSS.n12917 VSS.n2740 0.0316203
R7702 VSS.n12927 VSS.n2726 0.0316203
R7703 VSS.n12927 VSS.n12926 0.0316203
R7704 VSS.n12994 VSS.n2556 0.0316203
R7705 VSS.n12994 VSS.n2559 0.0316203
R7706 VSS.n13002 VSS.n2551 0.0316203
R7707 VSS.n13002 VSS.n13001 0.0316203
R7708 VSS.n12837 VSS.n2923 0.0316203
R7709 VSS.n12835 VSS.n2923 0.0316203
R7710 VSS.n13992 VSS.n1755 0.0316203
R7711 VSS.n13993 VSS.n13992 0.0316203
R7712 VSS.n14036 VSS.n1708 0.0316203
R7713 VSS.n14034 VSS.n1708 0.0316203
R7714 VSS.n13626 VSS.n13398 0.0316203
R7715 VSS.n13626 VSS.n13625 0.0316203
R7716 VSS.n702 VSS.n700 0.0314025
R7717 VSS.n4028 VSS.n3969 0.0307083
R7718 VSS.n12579 VSS.n3173 0.0307083
R7719 VSS.n3212 VSS.n3191 0.0307083
R7720 VSS.n3343 VSS.n3341 0.0303642
R7721 VSS.n3421 VSS.n3419 0.0303642
R7722 VSS.n11788 VSS.n11786 0.0303642
R7723 VSS.n11537 VSS.n11535 0.0303642
R7724 VSS.n979 VSS.n494 0.0303642
R7725 VSS.n13749 VSS.n481 0.0303642
R7726 VSS.n13287 VSS.n485 0.0303642
R7727 VSS.n1500 VSS.n449 0.0303642
R7728 VSS.n699 VSS.n446 0.0303642
R7729 VSS.n1237 VSS.n476 0.0303642
R7730 VSS.n14380 VSS.n14376 0.0303642
R7731 VSS.n3618 VSS.n3617 0.0303642
R7732 VSS.n11762 VSS.n11761 0.0303642
R7733 VSS.n11906 VSS.n11905 0.0303642
R7734 VSS.n14460 VSS.n14459 0.0303642
R7735 VSS.n3957 VSS.n3956 0.0286252
R7736 VSS.n5427 VSS.n5425 0.028625
R7737 VSS.n6107 VSS.n6106 0.0283475
R7738 VSS.n5925 VSS.n5924 0.0283475
R7739 VSS.n11396 VSS 0.0278438
R7740 VSS.n11378 VSS 0.0278438
R7741 VSS.n11360 VSS 0.0278438
R7742 VSS.n11118 VSS.n3821 0.0278438
R7743 VSS.n11003 VSS.n3843 0.0278438
R7744 VSS.n10959 VSS.n3889 0.0278438
R7745 VSS.n10850 VSS.n10849 0.0278438
R7746 VSS.n4355 VSS.n4206 0.0278438
R7747 VSS.n4438 VSS.n4156 0.0278438
R7748 VSS.n12829 VSS.n2926 0.0278438
R7749 VSS.n13999 VSS.n1749 0.0278438
R7750 VSS.n14028 VSS.n1711 0.0278438
R7751 VSS.n13614 VSS.n13613 0.0278438
R7752 VSS.n10135 VSS.n10134 0.0275833
R7753 VSS.n5557 VSS.n5556 0.0270627
R7754 VSS.n12463 VSS.n12364 0.0265417
R7755 VSS.n10715 VSS.n10652 0.0265417
R7756 VSS.n11931 VSS.n11929 0.0260208
R7757 VSS.n317 VSS.n277 0.02588
R7758 VSS.n14444 VSS.n261 0.02588
R7759 VSS.n14396 VSS.n306 0.02588
R7760 VSS.n14444 VSS.n279 0.02588
R7761 VSS.n14394 VSS.n334 0.02588
R7762 VSS.n14394 VSS.n352 0.02588
R7763 VSS.n14381 VSS.n444 0.02588
R7764 VSS.n14381 VSS.n491 0.02588
R7765 VSS.n14381 VSS.n483 0.02588
R7766 VSS.n14393 VSS.n14391 0.02588
R7767 VSS.n14394 VSS.n368 0.02588
R7768 VSS.n14455 VSS.n149 0.02588
R7769 VSS.n232 VSS.n188 0.02588
R7770 VSS.n14455 VSS.n167 0.02588
R7771 VSS.n125 VSS.n123 0.02588
R7772 VSS.n14455 VSS.n14453 0.02588
R7773 VSS.n198 VSS.n182 0.02588
R7774 VSS.n328 VSS.n303 0.02588
R7775 VSS.n14444 VSS.n304 0.02588
R7776 VSS.n14444 VSS.n308 0.02588
R7777 VSS.n14455 VSS.n196 0.02588
R7778 VSS.n203 VSS.n184 0.02588
R7779 VSS.n214 VSS.n192 0.02588
R7780 VSS.n14443 VSS.n14441 0.02588
R7781 VSS.n387 VSS.n370 0.02588
R7782 VSS.n14394 VSS.n364 0.02588
R7783 VSS.n396 VSS.n366 0.02588
R7784 VSS.n14381 VSS.n479 0.02588
R7785 VSS.n14381 VSS.n477 0.02588
R7786 VSS.n14381 VSS.n473 0.02588
R7787 VSS.n436 VSS.n357 0.02588
R7788 VSS.n427 VSS.n354 0.02588
R7789 VSS.n14394 VSS.n362 0.02588
R7790 VSS.n14394 VSS.n358 0.02588
R7791 VSS.n14425 VSS.n284 0.02588
R7792 VSS.n14406 VSS.n281 0.02588
R7793 VSS.n14444 VSS.n289 0.02588
R7794 VSS.n14444 VSS.n285 0.02588
R7795 VSS.n223 VSS.n195 0.02588
R7796 VSS.n14455 VSS.n186 0.02588
R7797 VSS.n14455 VSS.n190 0.02588
R7798 VSS.n79 VSS.n77 0.02588
R7799 VSS.n64 VSS.n62 0.02588
R7800 VSS.n253 VSS.n169 0.02588
R7801 VSS.n242 VSS.n163 0.02588
R7802 VSS.n14418 VSS.n288 0.02588
R7803 VSS.n408 VSS.n361 0.02588
R7804 VSS.n417 VSS.n350 0.02588
R7805 VSS.n14381 VSS.n500 0.02588
R7806 VSS.n14394 VSS.n347 0.02588
R7807 VSS.n14444 VSS.n274 0.02588
R7808 VSS.n14455 VSS.n164 0.02588
R7809 VSS.n67 VSS.n51 0.02588
R7810 VSS.n112 VSS.n110 0.02588
R7811 VSS.n138 VSS.n136 0.02588
R7812 VSS.n14461 VSS.n49 0.02588
R7813 VSS.n984 VSS.n980 0.0252925
R7814 VSS.n13751 VSS.n13750 0.0245875
R7815 VSS.n13289 VSS.n13288 0.0245875
R7816 VSS.n1505 VSS.n1501 0.0245875
R7817 VSS.n24 VSS 0.024
R7818 VSS VSS 0.024
R7819 VSS.n4522 VSS 0.024
R7820 VSS.n4531 VSS 0.024
R7821 VSS.n4482 VSS 0.024
R7822 VSS.n4480 VSS 0.024
R7823 VSS VSS 0.024
R7824 VSS VSS 0.024
R7825 VSS VSS 0.024
R7826 VSS VSS.n496 0.024
R7827 VSS.n11355 VSS 0.0239375
R7828 VSS.n3665 VSS 0.0239375
R7829 VSS.n3657 VSS 0.0239375
R7830 VSS VSS.n11243 0.0239375
R7831 VSS.n11251 VSS 0.0239375
R7832 VSS.n11495 VSS.n11494 0.0233646
R7833 VSS.n1239 VSS.n1238 0.023295
R7834 VSS.n8430 VSS.n8429 0.0228958
R7835 VSS.n8627 VSS.n8625 0.0228958
R7836 VSS.n8711 VSS.n8710 0.0228958
R7837 VSS.n9702 VSS.n9700 0.0228958
R7838 VSS.n11351 VSS 0.0226354
R7839 VSS.n3670 VSS 0.0226354
R7840 VSS.n11236 VSS 0.0226354
R7841 VSS.n276 VSS 0.0224565
R7842 VSS.n273 VSS 0.0224565
R7843 VSS.n287 VSS 0.0224565
R7844 VSS.n278 VSS 0.0224565
R7845 VSS.n305 VSS 0.0224565
R7846 VSS.n290 VSS 0.0224565
R7847 VSS.n302 VSS 0.0224565
R7848 VSS.n309 VSS 0.0224565
R7849 VSS.n360 VSS 0.0224565
R7850 VSS.n351 VSS 0.0224565
R7851 VSS.n369 VSS 0.0224565
R7852 VSS.n367 VSS 0.0224565
R7853 VSS.n501 VSS 0.0224565
R7854 VSS.n492 VSS 0.0224565
R7855 VSS.n482 VSS 0.0224565
R7856 VSS.n486 VSS 0.0224565
R7857 VSS.n14392 VSS 0.0224565
R7858 VSS.n371 VSS 0.0224565
R7859 VSS.n168 VSS 0.0224565
R7860 VSS.n166 VSS 0.0224565
R7861 VSS.n187 VSS 0.0224565
R7862 VSS.n170 VSS 0.0224565
R7863 VSS.n124 VSS 0.0224565
R7864 VSS.n42 VSS 0.0224565
R7865 VSS.n137 VSS 0.0224565
R7866 VSS.n41 VSS 0.0224565
R7867 VSS.n48 VSS 0.0224565
R7868 VSS.n46 VSS 0.0224565
R7869 VSS.n181 VSS 0.0224565
R7870 VSS.n197 VSS 0.0224565
R7871 VSS.n14442 VSS 0.0224565
R7872 VSS.n307 VSS 0.0224565
R7873 VSS.n183 VSS 0.0224565
R7874 VSS.n185 VSS 0.0224565
R7875 VSS.n191 VSS 0.0224565
R7876 VSS.n193 VSS 0.0224565
R7877 VSS.n365 VSS 0.0224565
R7878 VSS.n363 VSS 0.0224565
R7879 VSS.n478 VSS 0.0224565
R7880 VSS.n447 VSS 0.0224565
R7881 VSS.n474 VSS 0.0224565
R7882 VSS.n356 VSS 0.0224565
R7883 VSS.n355 VSS 0.0224565
R7884 VSS.n353 VSS 0.0224565
R7885 VSS.n359 VSS 0.0224565
R7886 VSS.n283 VSS 0.0224565
R7887 VSS.n282 VSS 0.0224565
R7888 VSS.n280 VSS 0.0224565
R7889 VSS.n286 VSS 0.0224565
R7890 VSS.n194 VSS 0.0224565
R7891 VSS.n189 VSS 0.0224565
R7892 VSS.n66 VSS 0.0224565
R7893 VSS.n44 VSS 0.0224565
R7894 VSS.n111 VSS 0.0224565
R7895 VSS.n40 VSS 0.0224565
R7896 VSS.n63 VSS 0.0224565
R7897 VSS.n39 VSS 0.0224565
R7898 VSS.n50 VSS 0.0224565
R7899 VSS.n43 VSS 0.0224565
R7900 VSS.n162 VSS 0.0224565
R7901 VSS.n161 VSS 0.0224565
R7902 VSS.n349 VSS 0.0224565
R7903 VSS.n346 VSS 0.0224565
R7904 VSS.n4487 VSS.n4482 0.0220983
R7905 VSS.n13419 VSS 0.0216803
R7906 VSS.n8340 VSS.n8339 0.0213335
R7907 VSS.n8322 VSS.n8321 0.0213335
R7908 VSS.n7517 VSS.n7516 0.0213335
R7909 VSS.n9726 VSS.n9725 0.0213335
R7910 VSS VSS.n13240 0.0213333
R7911 VSS.n13942 VSS 0.0213333
R7912 VSS.n12750 VSS 0.0213333
R7913 VSS.n3274 VSS 0.0213333
R7914 VSS.n12586 VSS.n12585 0.0213333
R7915 VSS.n3561 VSS.n3560 0.0213333
R7916 VSS.n11989 VSS.n11988 0.0213333
R7917 VSS.n12157 VSS.n12156 0.0213333
R7918 VSS.n12852 VSS.n2903 0.0213333
R7919 VSS.n12915 VSS.n2741 0.0213333
R7920 VSS.n768 VSS.n767 0.0213333
R7921 VSS.n11357 VSS 0.0213333
R7922 VSS VSS.n7351 0.0213333
R7923 VSS.n10967 VSS 0.0213333
R7924 VSS VSS.n6405 0.0213333
R7925 VSS.n11126 VSS 0.0213333
R7926 VSS.n10097 VSS.n10095 0.0213333
R7927 VSS.n5363 VSS.n5361 0.0213333
R7928 VSS.n5543 VSS.n5541 0.0213333
R7929 VSS.n5723 VSS.n5721 0.0213333
R7930 VSS.n6988 VSS.n6986 0.0213333
R7931 VSS.n9115 VSS.n9114 0.0213333
R7932 VSS.n9703 VSS.n9695 0.0213333
R7933 VSS.n9121 VSS.n9120 0.0213333
R7934 VSS.n9143 VSS.n9142 0.0213333
R7935 VSS.n9233 VSS.n7565 0.0213333
R7936 VSS VSS.n7999 0.0213333
R7937 VSS.n8563 VSS.n8562 0.0213333
R7938 VSS VSS.n8509 0.0213333
R7939 VSS VSS.n8389 0.0213333
R7940 VSS VSS.n8408 0.0213333
R7941 VSS.n8708 VSS.n8707 0.0213333
R7942 VSS.n9640 VSS.n9639 0.0213333
R7943 VSS.n9612 VSS.n9611 0.0213333
R7944 VSS.n8628 VSS.n8620 0.0213333
R7945 VSS.n8734 VSS.n8733 0.0213333
R7946 VSS.n8755 VSS.n8754 0.0213333
R7947 VSS VSS.n8285 0.0213333
R7948 VSS.n8771 VSS 0.0213333
R7949 VSS.n9547 VSS.n7588 0.0213333
R7950 VSS.n8795 VSS.n8794 0.0213333
R7951 VSS VSS.n6737 0.0213333
R7952 VSS VSS.n6208 0.0213333
R7953 VSS.n6739 VSS 0.0213333
R7954 VSS.n6769 VSS.n6767 0.0213333
R7955 VSS.n9951 VSS 0.0213333
R7956 VSS VSS.n8157 0.0213333
R7957 VSS.n8087 VSS.n8075 0.0213333
R7958 VSS.n8075 VSS.n8074 0.0213333
R7959 VSS.n8000 VSS 0.0213333
R7960 VSS.n8901 VSS.n8899 0.0213333
R7961 VSS.n8849 VSS 0.0213333
R7962 VSS VSS.n8007 0.0213333
R7963 VSS.n8810 VSS.n8795 0.0213333
R7964 VSS.n9548 VSS.n9547 0.0213333
R7965 VSS VSS.n7549 0.0213333
R7966 VSS VSS.n9596 0.0213333
R7967 VSS.n8529 VSS.n8528 0.0213333
R7968 VSS.n8434 VSS 0.0213333
R7969 VSS.n9793 VSS.n9792 0.0213333
R7970 VSS.n9427 VSS.n9420 0.0213333
R7971 VSS.n9776 VSS.n9775 0.0213333
R7972 VSS.n10840 VSS.n10839 0.0213333
R7973 VSS.n7478 VSS.n7477 0.0213333
R7974 VSS.n10823 VSS.n10822 0.0213333
R7975 VSS.n4025 VSS.n4024 0.0213333
R7976 VSS.n9431 VSS.n9430 0.0213333
R7977 VSS.n9452 VSS.n9451 0.0213333
R7978 VSS.n9845 VSS.n7156 0.0213333
R7979 VSS.n9271 VSS 0.0213333
R7980 VSS.n9487 VSS 0.0213333
R7981 VSS VSS.n9486 0.0213333
R7982 VSS.n7241 VSS.n7240 0.0213333
R7983 VSS.n9845 VSS.n9844 0.0213333
R7984 VSS.n7242 VSS.n7241 0.0213333
R7985 VSS.n7363 VSS 0.0213333
R7986 VSS.n7330 VSS.n7329 0.0213333
R7987 VSS VSS.n7380 0.0213333
R7988 VSS.n9809 VSS 0.0213333
R7989 VSS VSS.n9270 0.0213333
R7990 VSS.n9234 VSS.n9233 0.0213333
R7991 VSS.n9523 VSS.n8992 0.0213333
R7992 VSS.n9523 VSS.n9522 0.0213333
R7993 VSS VSS.n7918 0.0213333
R7994 VSS.n8965 VSS.n8963 0.0213333
R7995 VSS VSS.n7609 0.0213333
R7996 VSS VSS.n8991 0.0213333
R7997 VSS.n7755 VSS.n7753 0.0213333
R7998 VSS.n8966 VSS.n8965 0.0213333
R7999 VSS.n7782 VSS 0.0213333
R8000 VSS VSS.n7781 0.0213333
R8001 VSS.n9899 VSS.n7068 0.0213333
R8002 VSS.n7756 VSS.n7755 0.0213333
R8003 VSS.n9899 VSS.n9898 0.0213333
R8004 VSS VSS.n3881 0.0213333
R8005 VSS.n10994 VSS.n3851 0.0213333
R8006 VSS.n9866 VSS 0.0213333
R8007 VSS VSS.n7145 0.0213333
R8008 VSS.n7920 VSS 0.0213333
R8009 VSS.n8916 VSS.n8901 0.0213333
R8010 VSS.n8940 VSS.n8938 0.0213333
R8011 VSS.n8941 VSS.n8940 0.0213333
R8012 VSS.n6915 VSS.n6913 0.0213333
R8013 VSS VSS.n6812 0.0213333
R8014 VSS.n6881 VSS 0.0213333
R8015 VSS VSS.n6880 0.0213333
R8016 VSS.n6916 VSS.n6915 0.0213333
R8017 VSS.n6954 VSS 0.0213333
R8018 VSS VSS.n6953 0.0213333
R8019 VSS.n7047 VSS.n7045 0.0213333
R8020 VSS.n6989 VSS.n6988 0.0213333
R8021 VSS.n7034 VSS 0.0213333
R8022 VSS VSS.n7033 0.0213333
R8023 VSS.n6462 VSS.n6461 0.0213333
R8024 VSS.n7048 VSS.n7047 0.0213333
R8025 VSS.n6461 VSS.n6460 0.0213333
R8026 VSS.n6417 VSS 0.0213333
R8027 VSS.n6384 VSS.n6383 0.0213333
R8028 VSS VSS.n6269 0.0213333
R8029 VSS VSS.n7066 0.0213333
R8030 VSS.n6814 VSS 0.0213333
R8031 VSS.n6781 VSS.n6769 0.0213333
R8032 VSS.n6848 VSS.n6846 0.0213333
R8033 VSS.n6849 VSS.n6848 0.0213333
R8034 VSS.n5904 VSS.n5902 0.0213333
R8035 VSS VSS.n6047 0.0213333
R8036 VSS.n6033 VSS.n5970 0.0213333
R8037 VSS.n5850 VSS 0.0213333
R8038 VSS VSS.n5849 0.0213333
R8039 VSS.n5835 VSS.n5789 0.0213333
R8040 VSS.n5669 VSS 0.0213333
R8041 VSS VSS.n5668 0.0213333
R8042 VSS.n5654 VSS.n5608 0.0213333
R8043 VSS.n5489 VSS 0.0213333
R8044 VSS VSS.n5488 0.0213333
R8045 VSS.n5474 VSS.n5428 0.0213333
R8046 VSS.n5309 VSS 0.0213333
R8047 VSS VSS.n5308 0.0213333
R8048 VSS.n5294 VSS.n5248 0.0213333
R8049 VSS.n10099 VSS.n4573 0.0213333
R8050 VSS VSS.n3813 0.0213333
R8051 VSS.n3784 VSS.n3783 0.0213333
R8052 VSS VSS.n4631 0.0213333
R8053 VSS.n10043 VSS 0.0213333
R8054 VSS.n6049 VSS 0.0213333
R8055 VSS.n6086 VSS.n6084 0.0213333
R8056 VSS.n5727 VSS.n5726 0.0213333
R8057 VSS.n11142 VSS.n11141 0.0213333
R8058 VSS VSS.n11112 0.0213333
R8059 VSS.n6385 VSS.n6384 0.0213333
R8060 VSS.n11008 VSS 0.0213333
R8061 VSS.n10994 VSS.n10993 0.0213333
R8062 VSS VSS.n10953 0.0213333
R8063 VSS.n7331 VSS.n7330 0.0213333
R8064 VSS.n10857 VSS 0.0213333
R8065 VSS VSS.n4088 0.0213333
R8066 VSS VSS.n10782 0.0213333
R8067 VSS.n4384 VSS 0.0213333
R8068 VSS.n4277 VSS 0.0213333
R8069 VSS VSS.n4350 0.0213333
R8070 VSS VSS.n4411 0.0213333
R8071 VSS.n10748 VSS 0.0213333
R8072 VSS.n1327 VSS.n1301 0.0213333
R8073 VSS.n774 VSS.n773 0.0213333
R8074 VSS.n796 VSS.n795 0.0213333
R8075 VSS.n1077 VSS.n1052 0.0213333
R8076 VSS.n1332 VSS.n1331 0.0213333
R8077 VSS.n1353 VSS.n1352 0.0213333
R8078 VSS.n1403 VSS.n1401 0.0213333
R8079 VSS VSS.n955 0.0213333
R8080 VSS VSS.n2324 0.0213333
R8081 VSS.n1082 VSS.n1081 0.0213333
R8082 VSS.n14208 VSS 0.0213333
R8083 VSS VSS.n14235 0.0213333
R8084 VSS VSS.n10709 0.0213333
R8085 VSS.n14367 VSS.n14280 0.0213333
R8086 VSS.n14253 VSS.n14252 0.0213333
R8087 VSS VSS.n14207 0.0213333
R8088 VSS.n1130 VSS 0.0213333
R8089 VSS.n1159 VSS.n1157 0.0213333
R8090 VSS.n14175 VSS.n14174 0.0213333
R8091 VSS VSS.n13029 0.0213333
R8092 VSS.n12432 VSS 0.0213333
R8093 VSS.n13041 VSS 0.0213333
R8094 VSS.n13004 VSS.n2548 0.0213333
R8095 VSS VSS.n13059 0.0213333
R8096 VSS.n2446 VSS 0.0213333
R8097 VSS.n13140 VSS.n1909 0.0213333
R8098 VSS.n13140 VSS.n13139 0.0213333
R8099 VSS.n2326 VSS 0.0213333
R8100 VSS.n2299 VSS.n2297 0.0213333
R8101 VSS.n13107 VSS 0.0213333
R8102 VSS VSS.n13106 0.0213333
R8103 VSS.n14174 VSS.n14173 0.0213333
R8104 VSS.n1160 VSS.n1159 0.0213333
R8105 VSS VSS.n1196 0.0213333
R8106 VSS.n1369 VSS 0.0213333
R8107 VSS.n1114 VSS.n1113 0.0213333
R8108 VSS.n14363 VSS.n14337 0.0213333
R8109 VSS.n13861 VSS.n13860 0.0213333
R8110 VSS.n1599 VSS.n1574 0.0213333
R8111 VSS.n13844 VSS.n13843 0.0213333
R8112 VSS.n13396 VSS.n13395 0.0213333
R8113 VSS.n13839 VSS.n13814 0.0213333
R8114 VSS.n13379 VSS.n13378 0.0213333
R8115 VSS.n13374 VSS.n13349 0.0213333
R8116 VSS.n1603 VSS.n1602 0.0213333
R8117 VSS.n1624 VSS.n1623 0.0213333
R8118 VSS.n14059 VSS.n1696 0.0213333
R8119 VSS.n1441 VSS 0.0213333
R8120 VSS.n14086 VSS 0.0213333
R8121 VSS VSS.n14085 0.0213333
R8122 VSS.n13910 VSS.n13202 0.0213333
R8123 VSS.n14060 VSS.n14059 0.0213333
R8124 VSS.n13910 VSS.n13909 0.0213333
R8125 VSS.n13639 VSS 0.0213333
R8126 VSS.n13549 VSS.n13547 0.0213333
R8127 VSS.n13877 VSS 0.0213333
R8128 VSS VSS.n13703 0.0213333
R8129 VSS VSS.n1440 0.0213333
R8130 VSS.n1404 VSS.n1403 0.0213333
R8131 VSS.n14122 VSS.n626 0.0213333
R8132 VSS.n14122 VSS.n14121 0.0213333
R8133 VSS.n2035 VSS 0.0213333
R8134 VSS.n2205 VSS.n2188 0.0213333
R8135 VSS.n2216 VSS 0.0213333
R8136 VSS.n2084 VSS 0.0213333
R8137 VSS.n13182 VSS.n1880 0.0213333
R8138 VSS.n2188 VSS.n2186 0.0213333
R8139 VSS.n2151 VSS 0.0213333
R8140 VSS VSS.n2150 0.0213333
R8141 VSS.n12694 VSS.n12668 0.0213333
R8142 VSS.n13183 VSS.n13182 0.0213333
R8143 VSS.n12694 VSS.n12693 0.0213333
R8144 VSS VSS.n13940 0.0213333
R8145 VSS.n13990 VSS.n1757 0.0213333
R8146 VSS.n13915 VSS 0.0213333
R8147 VSS VSS.n13201 0.0213333
R8148 VSS VSS.n2034 0.0213333
R8149 VSS.n2300 VSS.n2299 0.0213333
R8150 VSS.n2254 VSS.n2253 0.0213333
R8151 VSS.n2253 VSS.n2251 0.0213333
R8152 VSS.n12929 VSS.n2723 0.0213333
R8153 VSS.n2642 VSS 0.0213333
R8154 VSS.n12956 VSS 0.0213333
R8155 VSS VSS.n12955 0.0213333
R8156 VSS.n12930 VSS.n12929 0.0213333
R8157 VSS VSS.n2821 0.0213333
R8158 VSS.n2823 VSS 0.0213333
R8159 VSS.n12915 VSS.n12914 0.0213333
R8160 VSS.n12879 VSS 0.0213333
R8161 VSS VSS.n12878 0.0213333
R8162 VSS.n12616 VSS.n12615 0.0213333
R8163 VSS.n12853 VSS.n12852 0.0213333
R8164 VSS.n12615 VSS.n3084 0.0213333
R8165 VSS VSS.n12735 0.0213333
R8166 VSS.n3000 VSS.n2999 0.0213333
R8167 VSS.n12710 VSS 0.0213333
R8168 VSS VSS.n12644 0.0213333
R8169 VSS VSS.n2641 0.0213333
R8170 VSS.n13005 VSS.n13004 0.0213333
R8171 VSS.n12992 VSS.n2560 0.0213333
R8172 VSS.n12992 VSS.n12991 0.0213333
R8173 VSS.n12264 VSS.n12263 0.0213333
R8174 VSS.n11637 VSS 0.0213333
R8175 VSS.n12341 VSS.n11681 0.0213333
R8176 VSS.n12211 VSS 0.0213333
R8177 VSS.n11706 VSS 0.0213333
R8178 VSS.n12208 VSS.n11750 0.0213333
R8179 VSS.n12104 VSS 0.0213333
R8180 VSS VSS.n12103 0.0213333
R8181 VSS.n12089 VSS.n12044 0.0213333
R8182 VSS.n11936 VSS 0.0213333
R8183 VSS.n11838 VSS 0.0213333
R8184 VSS.n11933 VSS.n11882 0.0213333
R8185 VSS.n3508 VSS 0.0213333
R8186 VSS VSS.n3507 0.0213333
R8187 VSS.n3493 VSS.n3448 0.0213333
R8188 VSS.n12583 VSS.n3171 0.0213333
R8189 VSS VSS.n3272 0.0213333
R8190 VSS.n3244 VSS.n3188 0.0213333
R8191 VSS VSS.n3085 0.0213333
R8192 VSS VSS.n12610 0.0213333
R8193 VSS VSS.n11636 0.0213333
R8194 VSS.n12343 VSS.n11568 0.0213333
R8195 VSS.n3288 VSS.n3287 0.0213333
R8196 VSS VSS.n12823 0.0213333
R8197 VSS.n2999 VSS.n2998 0.0213333
R8198 VSS.n12762 VSS 0.0213333
R8199 VSS.n13990 VSS.n13989 0.0213333
R8200 VSS VSS.n14022 0.0213333
R8201 VSS.n13550 VSS.n13549 0.0213333
R8202 VSS VSS.n13609 0.0213333
R8203 VSS.n13430 VSS 0.0213333
R8204 VSS.n3 VSS.n2 0.0211485
R8205 VSS VSS.n3 0.0211485
R8206 VSS.n11080 VSS.n11079 0.0208125
R8207 VSS.n14375 VSS.n14374 0.0205925
R8208 VSS.n5247 VSS.n5245 0.0202917
R8209 VSS.n3203 VSS.n3201 0.02024
R8210 VSS.n3204 VSS.n3203 0.02024
R8211 VSS.n3350 VSS.n3348 0.02024
R8212 VSS.n3351 VSS.n3350 0.02024
R8213 VSS.n11913 VSS.n11911 0.02024
R8214 VSS.n11914 VSS.n11913 0.02024
R8215 VSS.n11769 VSS.n11767 0.02024
R8216 VSS.n11770 VSS.n11769 0.02024
R8217 VSS.n1059 VSS.n1058 0.02024
R8218 VSS.n1060 VSS.n1059 0.02024
R8219 VSS.n13821 VSS.n13820 0.02024
R8220 VSS.n13822 VSS.n13821 0.02024
R8221 VSS.n13358 VSS.n13357 0.02024
R8222 VSS.n13359 VSS.n13358 0.02024
R8223 VSS.n1581 VSS.n1580 0.02024
R8224 VSS.n1582 VSS.n1581 0.02024
R8225 VSS.n451 VSS.n450 0.02024
R8226 VSS.n470 VSS.n450 0.02024
R8227 VSS.n1309 VSS.n1308 0.02024
R8228 VSS.n1310 VSS.n1309 0.02024
R8229 VSS.n14345 VSS.n14344 0.02024
R8230 VSS.n14346 VSS.n14345 0.02024
R8231 VSS.n11544 VSS.n11542 0.02024
R8232 VSS.n11545 VSS.n11544 0.02024
R8233 VSS.n11793 VSS.n11792 0.02024
R8234 VSS.n11794 VSS.n11793 0.02024
R8235 VSS.n3428 VSS.n3426 0.02024
R8236 VSS.n3429 VSS.n3428 0.02024
R8237 VSS.n4534 VSS 0.0198529
R8238 VSS.n4525 VSS 0.0198529
R8239 VSS.n295 VSS 0.0195238
R8240 VSS.n4524 VSS.n4522 0.0195238
R8241 VSS.n4519 VSS 0.0195238
R8242 VSS VSS.n4530 0.0195238
R8243 VSS.n4533 VSS.n4531 0.0195238
R8244 VSS.n4462 VSS 0.0195238
R8245 VSS.n4473 VSS 0.0195238
R8246 VSS VSS.n4497 0.0195238
R8247 VSS VSS.n4511 0.0195238
R8248 VSS VSS.n13418 0.0195238
R8249 VSS.n377 VSS 0.0195238
R8250 VSS.n31 VSS 0.0195238
R8251 VSS.n174 VSS 0.0195238
R8252 VSS.n497 VSS 0.0195238
R8253 VSS VSS.n342 0.0195238
R8254 VSS VSS.n269 0.0195238
R8255 VSS VSS.n157 0.0195238
R8256 VSS VSS.n96 0.0195238
R8257 VSS.n3446 VSS.n3444 0.01925
R8258 VSS.n3292 VSS.n3291 0.0187292
R8259 VSS.n12811 VSS.n12810 0.0187292
R8260 VSS.n5367 VSS.n5366 0.0182083
R8261 VSS.n13574 VSS.n13240 0.0178611
R8262 VSS.n13962 VSS.n13942 0.0178611
R8263 VSS.n12751 VSS.n12750 0.0178611
R8264 VSS.n3275 VSS.n3274 0.0178611
R8265 VSS.n767 VSS.n766 0.0178611
R8266 VSS.n7351 VSS.n7279 0.0178611
R8267 VSS.n10983 VSS.n10967 0.0178611
R8268 VSS.n6405 VSS.n6333 0.0178611
R8269 VSS.n11127 VSS.n11126 0.0178611
R8270 VSS.n9114 VSS.n9113 0.0178611
R8271 VSS.n9695 VSS.n9694 0.0178611
R8272 VSS.n7999 VSS.n7998 0.0178611
R8273 VSS.n8509 VSS.n8508 0.0178611
R8274 VSS.n8408 VSS.n8407 0.0178611
R8275 VSS.n8707 VSS.n8706 0.0178611
R8276 VSS.n8620 VSS.n8619 0.0178611
R8277 VSS.n8285 VSS.n8284 0.0178611
R8278 VSS.n6737 VSS.n6736 0.0178611
R8279 VSS.n6208 VSS.n6207 0.0178611
R8280 VSS.n9971 VSS.n9951 0.0178611
R8281 VSS.n8157 VSS.n8156 0.0178611
R8282 VSS.n8849 VSS.n8004 0.0178611
R8283 VSS.n9207 VSS.n7549 0.0178611
R8284 VSS.n8435 VSS.n8434 0.0178611
R8285 VSS.n9420 VSS.n9419 0.0178611
R8286 VSS.n7477 VSS.n7476 0.0178611
R8287 VSS.n4024 VSS.n4023 0.0178611
R8288 VSS.n9288 VSS.n9271 0.0178611
R8289 VSS.n9486 VSS.n9468 0.0178611
R8290 VSS.n7380 VSS.n7379 0.0178611
R8291 VSS.n7918 VSS.n7894 0.0178611
R8292 VSS.n8991 VSS.n7610 0.0178611
R8293 VSS.n7781 VSS.n7645 0.0178611
R8294 VSS.n9886 VSS.n9866 0.0178611
R8295 VSS.n6812 VSS.n6794 0.0178611
R8296 VSS.n6880 VSS.n6862 0.0178611
R8297 VSS.n6953 VSS.n6929 0.0178611
R8298 VSS.n7033 VSS.n7015 0.0178611
R8299 VSS.n6448 VSS.n6269 0.0178611
R8300 VSS.n6047 VSS.n6046 0.0178611
R8301 VSS.n5849 VSS.n5848 0.0178611
R8302 VSS.n5668 VSS.n5667 0.0178611
R8303 VSS.n5488 VSS.n5487 0.0178611
R8304 VSS.n5308 VSS.n5307 0.0178611
R8305 VSS.n4631 VSS.n4630 0.0178611
R8306 VSS.n10782 VSS.n4107 0.0178611
R8307 VSS.n4297 VSS.n4277 0.0178611
R8308 VSS.n4411 VSS.n4410 0.0178611
R8309 VSS.n1301 VSS.n1300 0.0178611
R8310 VSS.n1052 VSS.n1051 0.0178611
R8311 VSS.n955 VSS.n954 0.0178611
R8312 VSS.n2324 VSS.n2323 0.0178611
R8313 VSS.n14235 VSS.n14234 0.0178611
R8314 VSS.n10709 VSS.n10708 0.0178611
R8315 VSS.n14207 VSS.n14206 0.0178611
R8316 VSS.n13029 VSS.n13028 0.0178611
R8317 VSS.n12433 VSS.n12432 0.0178611
R8318 VSS.n13059 VSS.n13058 0.0178611
R8319 VSS.n2447 VSS.n2446 0.0178611
R8320 VSS.n13127 VSS.n13107 0.0178611
R8321 VSS.n1196 VSS.n1195 0.0178611
R8322 VSS.n14337 VSS.n14336 0.0178611
R8323 VSS.n1574 VSS.n1573 0.0178611
R8324 VSS.n13814 VSS.n13813 0.0178611
R8325 VSS.n13349 VSS.n13348 0.0178611
R8326 VSS.n1458 VSS.n1441 0.0178611
R8327 VSS.n14085 VSS.n1640 0.0178611
R8328 VSS.n13897 VSS.n13877 0.0178611
R8329 VSS.n2052 VSS.n2035 0.0178611
R8330 VSS.n2101 VSS.n2084 0.0178611
R8331 VSS.n2150 VSS.n2132 0.0178611
R8332 VSS.n13915 VSS.n1816 0.0178611
R8333 VSS.n2659 VSS.n2642 0.0178611
R8334 VSS.n12955 VSS.n2667 0.0178611
R8335 VSS.n2840 VSS.n2823 0.0178611
R8336 VSS.n12878 VSS.n2847 0.0178611
R8337 VSS.n12710 VSS.n3021 0.0178611
R8338 VSS.n11638 VSS.n11637 0.0178611
R8339 VSS.n11707 VSS.n11706 0.0178611
R8340 VSS.n12103 VSS.n12102 0.0178611
R8341 VSS.n11839 VSS.n11838 0.0178611
R8342 VSS.n3507 VSS.n3506 0.0178611
R8343 VSS.n3158 VSS.n3085 0.0178611
R8344 VSS.n11814 VSS.n11813 0.0176877
R8345 VSS.n8514 VSS.n8489 0.0175455
R8346 VSS.n8514 VSS 0.0175455
R8347 VSS VSS.n8512 0.0175455
R8348 VSS.n8512 VSS 0.0175455
R8349 VSS.n9986 VSS.n4660 0.0175455
R8350 VSS.n9986 VSS 0.0175455
R8351 VSS VSS.n6211 0.0175455
R8352 VSS.n6211 VSS 0.0175455
R8353 VSS.n8122 VSS.n8121 0.0175455
R8354 VSS.n8122 VSS 0.0175455
R8355 VSS.n9948 VSS 0.0175455
R8356 VSS.n9948 VSS 0.0175455
R8357 VSS.n8835 VSS.n8014 0.0175455
R8358 VSS.n8835 VSS 0.0175455
R8359 VSS VSS.n8160 0.0175455
R8360 VSS.n8160 VSS 0.0175455
R8361 VSS VSS.n8563 0.0175455
R8362 VSS.n8629 VSS 0.0175455
R8363 VSS.n8733 VSS 0.0175455
R8364 VSS.n8320 VSS 0.0175455
R8365 VSS VSS.n9640 0.0175455
R8366 VSS.n9704 VSS 0.0175455
R8367 VSS.n9120 VSS 0.0175455
R8368 VSS.n9053 VSS 0.0175455
R8369 VSS.n10822 VSS 0.0175455
R8370 VSS.n3955 VSS 0.0175455
R8371 VSS.n9775 VSS.n7419 0.0175455
R8372 VSS.n9775 VSS 0.0175455
R8373 VSS.n7420 VSS 0.0175455
R8374 VSS.n9430 VSS 0.0175455
R8375 VSS.n9428 VSS 0.0175455
R8376 VSS.n6086 VSS 0.0175455
R8377 VSS VSS.n5970 0.0175455
R8378 VSS.n5970 VSS 0.0175455
R8379 VSS.n5904 VSS 0.0175455
R8380 VSS VSS.n5789 0.0175455
R8381 VSS.n5789 VSS 0.0175455
R8382 VSS.n5723 VSS 0.0175455
R8383 VSS VSS.n5608 0.0175455
R8384 VSS.n5608 VSS 0.0175455
R8385 VSS.n5543 VSS 0.0175455
R8386 VSS VSS.n5428 0.0175455
R8387 VSS.n5428 VSS 0.0175455
R8388 VSS.n5363 VSS 0.0175455
R8389 VSS VSS.n5248 0.0175455
R8390 VSS.n5248 VSS 0.0175455
R8391 VSS.n10097 VSS 0.0175455
R8392 VSS.n10099 VSS 0.0175455
R8393 VSS VSS.n10099 0.0175455
R8394 VSS.n3783 VSS 0.0175455
R8395 VSS.n11142 VSS 0.0175455
R8396 VSS VSS.n11142 0.0175455
R8397 VSS.n11116 VSS.n3823 0.0175455
R8398 VSS.n11116 VSS 0.0175455
R8399 VSS.n11113 VSS 0.0175455
R8400 VSS VSS.n11113 0.0175455
R8401 VSS.n11005 VSS.n3842 0.0175455
R8402 VSS.n11005 VSS 0.0175455
R8403 VSS VSS.n3844 0.0175455
R8404 VSS.n3844 VSS 0.0175455
R8405 VSS.n10957 VSS.n3891 0.0175455
R8406 VSS.n10957 VSS 0.0175455
R8407 VSS.n10954 VSS 0.0175455
R8408 VSS VSS.n10954 0.0175455
R8409 VSS.n10854 VSS.n3909 0.0175455
R8410 VSS.n10854 VSS 0.0175455
R8411 VSS VSS.n10852 0.0175455
R8412 VSS.n10852 VSS 0.0175455
R8413 VSS.n4090 VSS 0.0175455
R8414 VSS.n4155 VSS.n4152 0.0175455
R8415 VSS.n4155 VSS 0.0175455
R8416 VSS.n4440 VSS 0.0175455
R8417 VSS.n4440 VSS 0.0175455
R8418 VSS.n4357 VSS.n4203 0.0175455
R8419 VSS.n4357 VSS 0.0175455
R8420 VSS.n4274 VSS 0.0175455
R8421 VSS.n4274 VSS 0.0175455
R8422 VSS.n4227 VSS.n4226 0.0175455
R8423 VSS.n4226 VSS 0.0175455
R8424 VSS.n4353 VSS 0.0175455
R8425 VSS.n4353 VSS 0.0175455
R8426 VSS.n4436 VSS.n4159 0.0175455
R8427 VSS.n4436 VSS 0.0175455
R8428 VSS VSS.n4413 0.0175455
R8429 VSS.n4413 VSS 0.0175455
R8430 VSS.n14241 VSS.n543 0.0175455
R8431 VSS.n14241 VSS 0.0175455
R8432 VSS VSS.n14239 0.0175455
R8433 VSS.n14239 VSS 0.0175455
R8434 VSS.n12423 VSS.n12396 0.0175455
R8435 VSS.n12423 VSS 0.0175455
R8436 VSS.n12429 VSS 0.0175455
R8437 VSS.n12429 VSS 0.0175455
R8438 VSS.n13066 VSS.n2458 0.0175455
R8439 VSS.n13066 VSS 0.0175455
R8440 VSS.n13062 VSS 0.0175455
R8441 VSS.n13062 VSS 0.0175455
R8442 VSS.n2423 VSS.n2396 0.0175455
R8443 VSS.n2423 VSS 0.0175455
R8444 VSS.n2427 VSS 0.0175455
R8445 VSS.n2427 VSS 0.0175455
R8446 VSS.n14368 VSS.n14367 0.0175455
R8447 VSS.n14367 VSS 0.0175455
R8448 VSS.n14364 VSS 0.0175455
R8449 VSS.n1081 VSS.n995 0.0175455
R8450 VSS.n1081 VSS 0.0175455
R8451 VSS.n1078 VSS 0.0175455
R8452 VSS.n1331 VSS.n1246 0.0175455
R8453 VSS.n1331 VSS 0.0175455
R8454 VSS.n1328 VSS 0.0175455
R8455 VSS.n773 VSS 0.0175455
R8456 VSS.n687 VSS 0.0175455
R8457 VSS.n13378 VSS.n13294 0.0175455
R8458 VSS.n13378 VSS 0.0175455
R8459 VSS.n13375 VSS 0.0175455
R8460 VSS.n13843 VSS.n13757 0.0175455
R8461 VSS.n13843 VSS 0.0175455
R8462 VSS.n13840 VSS 0.0175455
R8463 VSS.n1602 VSS.n1516 0.0175455
R8464 VSS.n1602 VSS 0.0175455
R8465 VSS.n1600 VSS 0.0175455
R8466 VSS.n12344 VSS.n12343 0.0175455
R8467 VSS.n12343 VSS 0.0175455
R8468 VSS.n12341 VSS 0.0175455
R8469 VSS.n12341 VSS 0.0175455
R8470 VSS.n12264 VSS 0.0175455
R8471 VSS VSS.n12208 0.0175455
R8472 VSS.n12208 VSS 0.0175455
R8473 VSS.n12157 VSS 0.0175455
R8474 VSS VSS.n12044 0.0175455
R8475 VSS.n12044 VSS 0.0175455
R8476 VSS.n11989 VSS 0.0175455
R8477 VSS VSS.n11933 0.0175455
R8478 VSS.n11933 VSS 0.0175455
R8479 VSS.n3561 VSS 0.0175455
R8480 VSS VSS.n3448 0.0175455
R8481 VSS.n3448 VSS 0.0175455
R8482 VSS.n12585 VSS 0.0175455
R8483 VSS.n12583 VSS 0.0175455
R8484 VSS.n12583 VSS 0.0175455
R8485 VSS VSS.n3188 0.0175455
R8486 VSS.n3288 VSS 0.0175455
R8487 VSS.n3288 VSS 0.0175455
R8488 VSS.n12827 VSS.n2928 0.0175455
R8489 VSS.n12827 VSS 0.0175455
R8490 VSS.n12824 VSS 0.0175455
R8491 VSS VSS.n12824 0.0175455
R8492 VSS.n14001 VSS.n1746 0.0175455
R8493 VSS.n14001 VSS 0.0175455
R8494 VSS VSS.n1750 0.0175455
R8495 VSS.n1750 VSS 0.0175455
R8496 VSS.n14026 VSS.n1713 0.0175455
R8497 VSS.n14026 VSS 0.0175455
R8498 VSS.n14023 VSS 0.0175455
R8499 VSS VSS.n14023 0.0175455
R8500 VSS.n13612 VSS.n13401 0.0175455
R8501 VSS.n13612 VSS 0.0175455
R8502 VSS VSS.n13400 0.0175455
R8503 VSS VSS.n13400 0.0175455
R8504 VSS.n13478 VSS.n13477 0.0173919
R8505 VSS.n13591 VSS.n13590 0.0173919
R8506 VSS.n14004 VSS.n1745 0.0173919
R8507 VSS.n12802 VSS.n12801 0.0173919
R8508 VSS.n12587 VSS.n12586 0.0173919
R8509 VSS.n3560 VSS.n3559 0.0173919
R8510 VSS.n11988 VSS.n11987 0.0173919
R8511 VSS.n12156 VSS.n12155 0.0173919
R8512 VSS.n2903 VSS.n2902 0.0173919
R8513 VSS.n2789 VSS.n2741 0.0173919
R8514 VSS.n4059 VSS.n4058 0.0173919
R8515 VSS.n10897 VSS.n10896 0.0173919
R8516 VSS.n10941 VSS.n10921 0.0173919
R8517 VSS.n11048 VSS.n11047 0.0173919
R8518 VSS.n10095 VSS.n10094 0.0173919
R8519 VSS.n5361 VSS.n5360 0.0173919
R8520 VSS.n5541 VSS.n5540 0.0173919
R8521 VSS.n5721 VSS.n5720 0.0173919
R8522 VSS.n6986 VSS.n6985 0.0173919
R8523 VSS.n9122 VSS.n9121 0.0173919
R8524 VSS.n9142 VSS.n9141 0.0173919
R8525 VSS.n9684 VSS.n9683 0.0173919
R8526 VSS.n9563 VSS.n7565 0.0173919
R8527 VSS.n8562 VSS.n8561 0.0173919
R8528 VSS.n8487 VSS.n8486 0.0173919
R8529 VSS.n8389 VSS.n8388 0.0173919
R8530 VSS.n9639 VSS.n9638 0.0173919
R8531 VSS.n9613 VSS.n9612 0.0173919
R8532 VSS.n8696 VSS.n8695 0.0173919
R8533 VSS.n8735 VSS.n8734 0.0173919
R8534 VSS.n8607 VSS.n8606 0.0173919
R8535 VSS.n8754 VSS.n8753 0.0173919
R8536 VSS.n8772 VSS.n8771 0.0173919
R8537 VSS.n8237 VSS.n7588 0.0173919
R8538 VSS.n8794 VSS.n8793 0.0173919
R8539 VSS.n9983 VSS.n9982 0.0173919
R8540 VSS.n6746 VSS.n6739 0.0173919
R8541 VSS.n6767 VSS.n6766 0.0173919
R8542 VSS.n8099 VSS.n8007 0.0173919
R8543 VSS.n8088 VSS.n8087 0.0173919
R8544 VSS.n8146 VSS.n8125 0.0173919
R8545 VSS.n8074 VSS.n8073 0.0173919
R8546 VSS.n8878 VSS.n8000 0.0173919
R8547 VSS.n8899 VSS.n8898 0.0173919
R8548 VSS.n8811 VSS.n8810 0.0173919
R8549 VSS.n8832 VSS.n8831 0.0173919
R8550 VSS.n9549 VSS.n9548 0.0173919
R8551 VSS.n9596 VSS.n9595 0.0173919
R8552 VSS.n8530 VSS.n8529 0.0173919
R8553 VSS.n9792 VSS.n9791 0.0173919
R8554 VSS.n9407 VSS.n9406 0.0173919
R8555 VSS.n9777 VSS.n9776 0.0173919
R8556 VSS.n10839 VSS.n10838 0.0173919
R8557 VSS.n7464 VSS.n7463 0.0173919
R8558 VSS.n10824 VSS.n10823 0.0173919
R8559 VSS.n9432 VSS.n9431 0.0173919
R8560 VSS.n9101 VSS.n9100 0.0173919
R8561 VSS.n9451 VSS.n9450 0.0173919
R8562 VSS.n9294 VSS.n7156 0.0173919
R8563 VSS.n9522 VSS.n9521 0.0173919
R8564 VSS.n9508 VSS.n9487 0.0173919
R8565 VSS.n7240 VSS.n7216 0.0173919
R8566 VSS.n9844 VSS.n9843 0.0173919
R8567 VSS.n9830 VSS.n9809 0.0173919
R8568 VSS.n7242 VSS.n7211 0.0173919
R8569 VSS.n7364 VSS.n7363 0.0173919
R8570 VSS.n7329 VSS.n7312 0.0173919
R8571 VSS.n9270 VSS.n9269 0.0173919
R8572 VSS.n9235 VSS.n9234 0.0173919
R8573 VSS.n9260 VSS.n8992 0.0173919
R8574 VSS.n8963 VSS.n7808 0.0173919
R8575 VSS.n8942 VSS.n8941 0.0173919
R8576 VSS.n8953 VSS.n7609 0.0173919
R8577 VSS.n7753 VSS.n7729 0.0173919
R8578 VSS.n8982 VSS.n8966 0.0173919
R8579 VSS.n7803 VSS.n7782 0.0173919
R8580 VSS.n7694 VSS.n7068 0.0173919
R8581 VSS.n7772 VSS.n7756 0.0173919
R8582 VSS.n7724 VSS.n7145 0.0173919
R8583 VSS.n9898 VSS.n9897 0.0173919
R8584 VSS.n7134 VSS.n3881 0.0173919
R8585 VSS.n7112 VSS.n3851 0.0173919
R8586 VSS.n7936 VSS.n7920 0.0173919
R8587 VSS.n8917 VSS.n8916 0.0173919
R8588 VSS.n8938 VSS.n8937 0.0173919
R8589 VSS.n6913 VSS.n6912 0.0173919
R8590 VSS.n6850 VSS.n6849 0.0173919
R8591 VSS.n6902 VSS.n6881 0.0173919
R8592 VSS.n6917 VSS.n6916 0.0173919
R8593 VSS.n6975 VSS.n6954 0.0173919
R8594 VSS.n7045 VSS.n6510 0.0173919
R8595 VSS.n6990 VSS.n6989 0.0173919
R8596 VSS.n7035 VSS.n7034 0.0173919
R8597 VSS.n6462 VSS.n6292 0.0173919
R8598 VSS.n7049 VSS.n7048 0.0173919
R8599 VSS.n7066 VSS.n7065 0.0173919
R8600 VSS.n6460 VSS.n6459 0.0173919
R8601 VSS.n6418 VSS.n6417 0.0173919
R8602 VSS.n6383 VSS.n6366 0.0173919
R8603 VSS.n6834 VSS.n6814 0.0173919
R8604 VSS.n6782 VSS.n6781 0.0173919
R8605 VSS.n6846 VSS.n6845 0.0173919
R8606 VSS.n5902 VSS.n5901 0.0173919
R8607 VSS.n6034 VSS.n6033 0.0173919
R8608 VSS.n5851 VSS.n5850 0.0173919
R8609 VSS.n5836 VSS.n5835 0.0173919
R8610 VSS.n5670 VSS.n5669 0.0173919
R8611 VSS.n5655 VSS.n5654 0.0173919
R8612 VSS.n5490 VSS.n5489 0.0173919
R8613 VSS.n5475 VSS.n5474 0.0173919
R8614 VSS.n5310 VSS.n5309 0.0173919
R8615 VSS.n5295 VSS.n5294 0.0173919
R8616 VSS.n10044 VSS.n10043 0.0173919
R8617 VSS.n4581 VSS.n4573 0.0173919
R8618 VSS.n3813 VSS.n3812 0.0173919
R8619 VSS.n3785 VSS.n3784 0.0173919
R8620 VSS.n6050 VSS.n6049 0.0173919
R8621 VSS.n6084 VSS.n6083 0.0173919
R8622 VSS.n6156 VSS.n6155 0.0173919
R8623 VSS.n11083 VSS.n11082 0.0173919
R8624 VSS.n11141 VSS.n11140 0.0173919
R8625 VSS.n11112 VSS.n11111 0.0173919
R8626 VSS.n6386 VSS.n6385 0.0173919
R8627 VSS.n11024 VSS.n11008 0.0173919
R8628 VSS.n10993 VSS.n10992 0.0173919
R8629 VSS.n10953 VSS.n10952 0.0173919
R8630 VSS.n7332 VSS.n7331 0.0173919
R8631 VSS.n10873 VSS.n10857 0.0173919
R8632 VSS.n3976 VSS.n3975 0.0173919
R8633 VSS.n4088 VSS.n4087 0.0173919
R8634 VSS.n4444 VSS.n4443 0.0173919
R8635 VSS.n4400 VSS.n4384 0.0173919
R8636 VSS.n4376 VSS.n4360 0.0173919
R8637 VSS.n4332 VSS.n4259 0.0173919
R8638 VSS.n4324 VSS.n4323 0.0173919
R8639 VSS.n4350 VSS.n4349 0.0173919
R8640 VSS.n4225 VSS.n4208 0.0173919
R8641 VSS.n4433 VSS.n4432 0.0173919
R8642 VSS.n10769 VSS.n10748 0.0173919
R8643 VSS.n775 VSS.n774 0.0173919
R8644 VSS.n795 VSS.n794 0.0173919
R8645 VSS.n1290 VSS.n1289 0.0173919
R8646 VSS.n1333 VSS.n1332 0.0173919
R8647 VSS.n1039 VSS.n1038 0.0173919
R8648 VSS.n1352 VSS.n1351 0.0173919
R8649 VSS.n1401 VSS.n1400 0.0173919
R8650 VSS.n1083 VSS.n1082 0.0173919
R8651 VSS.n14308 VSS.n14307 0.0173919
R8652 VSS.n14224 VSS.n14208 0.0173919
R8653 VSS.n14280 VSS.n14279 0.0173919
R8654 VSS.n14254 VSS.n14253 0.0173919
R8655 VSS.n10698 VSS.n10697 0.0173919
R8656 VSS.n1136 VSS.n1130 0.0173919
R8657 VSS.n1157 VSS.n1156 0.0173919
R8658 VSS.n14196 VSS.n14175 0.0173919
R8659 VSS.n12420 VSS.n12419 0.0173919
R8660 VSS.n13042 VSS.n13041 0.0173919
R8661 VSS.n2548 VSS.n2531 0.0173919
R8662 VSS.n13106 VSS.n2350 0.0173919
R8663 VSS.n2390 VSS.n1909 0.0173919
R8664 VSS.n13090 VSS.n13069 0.0173919
R8665 VSS.n13139 VSS.n13138 0.0173919
R8666 VSS.n2327 VSS.n2326 0.0173919
R8667 VSS.n2297 VSS.n2296 0.0173919
R8668 VSS.n14173 VSS.n14154 0.0173919
R8669 VSS.n2420 VSS.n2419 0.0173919
R8670 VSS.n1161 VSS.n1160 0.0173919
R8671 VSS.n1390 VSS.n1369 0.0173919
R8672 VSS.n1113 VSS.n1112 0.0173919
R8673 VSS.n13860 VSS.n13859 0.0173919
R8674 VSS.n1561 VSS.n1560 0.0173919
R8675 VSS.n13845 VSS.n13844 0.0173919
R8676 VSS.n13395 VSS.n13394 0.0173919
R8677 VSS.n13801 VSS.n13800 0.0173919
R8678 VSS.n13380 VSS.n13379 0.0173919
R8679 VSS.n1604 VSS.n1603 0.0173919
R8680 VSS.n754 VSS.n753 0.0173919
R8681 VSS.n1623 VSS.n1622 0.0173919
R8682 VSS.n1696 VSS.n1672 0.0173919
R8683 VSS.n14121 VSS.n14120 0.0173919
R8684 VSS.n14107 VSS.n14086 0.0173919
R8685 VSS.n13672 VSS.n13202 0.0173919
R8686 VSS.n14076 VSS.n14060 0.0173919
R8687 VSS.n13703 VSS.n13702 0.0173919
R8688 VSS.n13909 VSS.n13908 0.0173919
R8689 VSS.n13640 VSS.n13639 0.0173919
R8690 VSS.n13547 VSS.n13530 0.0173919
R8691 VSS.n1440 VSS.n1439 0.0173919
R8692 VSS.n1405 VSS.n1404 0.0173919
R8693 VSS.n1430 VSS.n626 0.0173919
R8694 VSS.n2206 VSS.n2205 0.0173919
R8695 VSS.n2251 VSS.n2250 0.0173919
R8696 VSS.n2237 VSS.n2216 0.0173919
R8697 VSS.n2122 VSS.n1880 0.0173919
R8698 VSS.n2186 VSS.n2185 0.0173919
R8699 VSS.n2172 VSS.n2151 0.0173919
R8700 VSS.n12668 VSS.n12645 0.0173919
R8701 VSS.n13184 VSS.n13183 0.0173919
R8702 VSS.n13201 VSS.n13200 0.0173919
R8703 VSS.n12693 VSS.n12692 0.0173919
R8704 VSS.n13940 VSS.n1771 0.0173919
R8705 VSS.n1811 VSS.n1757 0.0173919
R8706 VSS.n2034 VSS.n2033 0.0173919
R8707 VSS.n2316 VSS.n2300 0.0173919
R8708 VSS.n2275 VSS.n2254 0.0173919
R8709 VSS.n2723 VSS.n2722 0.0173919
R8710 VSS.n12991 VSS.n12990 0.0173919
R8711 VSS.n12977 VSS.n12956 0.0173919
R8712 VSS.n12946 VSS.n12930 0.0173919
R8713 VSS.n2821 VSS.n2820 0.0173919
R8714 VSS.n12914 VSS.n12913 0.0173919
R8715 VSS.n12900 VSS.n12879 0.0173919
R8716 VSS.n12616 VSS.n3056 0.0173919
R8717 VSS.n12869 VSS.n12853 0.0173919
R8718 VSS.n12644 VSS.n12643 0.0173919
R8719 VSS.n3084 VSS.n3083 0.0173919
R8720 VSS.n12735 VSS.n2949 0.0173919
R8721 VSS.n3016 VSS.n3000 0.0173919
R8722 VSS.n2641 VSS.n2640 0.0173919
R8723 VSS.n13021 VSS.n13005 0.0173919
R8724 VSS.n2630 VSS.n2560 0.0173919
R8725 VSS.n12263 VSS.n12262 0.0173919
R8726 VSS.n11681 VSS.n11680 0.0173919
R8727 VSS.n12212 VSS.n12211 0.0173919
R8728 VSS.n11750 VSS.n11749 0.0173919
R8729 VSS.n12105 VSS.n12104 0.0173919
R8730 VSS.n12090 VSS.n12089 0.0173919
R8731 VSS.n11937 VSS.n11936 0.0173919
R8732 VSS.n11882 VSS.n11881 0.0173919
R8733 VSS.n3509 VSS.n3508 0.0173919
R8734 VSS.n3494 VSS.n3493 0.0173919
R8735 VSS.n12610 VSS.n12609 0.0173919
R8736 VSS.n3171 VSS.n3170 0.0173919
R8737 VSS.n3272 VSS.n3271 0.0173919
R8738 VSS.n3245 VSS.n3244 0.0173919
R8739 VSS.n11636 VSS.n11635 0.0173919
R8740 VSS.n11598 VSS.n11568 0.0173919
R8741 VSS.n12458 VSS.n12457 0.0173919
R8742 VSS.n12816 VSS.n12815 0.0173919
R8743 VSS.n3287 VSS.n3286 0.0173919
R8744 VSS.n12823 VSS.n12822 0.0173919
R8745 VSS.n2998 VSS.n2997 0.0173919
R8746 VSS.n12778 VSS.n12762 0.0173919
R8747 VSS.n13989 VSS.n13988 0.0173919
R8748 VSS.n14022 VSS.n14021 0.0173919
R8749 VSS.n13551 VSS.n13550 0.0173919
R8750 VSS.n13609 VSS.n13608 0.0173919
R8751 VSS.n13303 VSS.n13302 0.0173919
R8752 VSS.n13431 VSS.n13430 0.0173919
R8753 VSS.n3200 VSS 0.017343
R8754 VSS.n3205 VSS 0.017343
R8755 VSS.n3347 VSS 0.017343
R8756 VSS.n3352 VSS 0.017343
R8757 VSS.n3425 VSS 0.017343
R8758 VSS.n3430 VSS 0.017343
R8759 VSS.n11910 VSS 0.017343
R8760 VSS.n11915 VSS 0.017343
R8761 VSS VSS.n11784 0.017343
R8762 VSS VSS.n11795 0.017343
R8763 VSS.n11795 VSS 0.017343
R8764 VSS.n11766 VSS 0.017343
R8765 VSS.n11771 VSS 0.017343
R8766 VSS.n11541 VSS 0.017343
R8767 VSS.n11546 VSS 0.017343
R8768 VSS.n3206 VSS.n3205 0.0171826
R8769 VSS.n3353 VSS.n3352 0.0171826
R8770 VSS.n11916 VSS.n11915 0.0171826
R8771 VSS.n11772 VSS.n11771 0.0171826
R8772 VSS.n11547 VSS.n11546 0.0171826
R8773 VSS.n11993 VSS.n11992 0.0171667
R8774 VSS.n3431 VSS.n3430 0.0170222
R8775 VSS VSS.n14511 0.0168222
R8776 VSS.n5377 VSS.n5376 0.016646
R8777 VSS.n14445 VSS.n240 0.0163425
R8778 VSS.n14382 VSS.n393 0.0163425
R8779 VSS.n14382 VSS.n443 0.0163425
R8780 VSS.n14435 VSS.n14434 0.0163425
R8781 VSS.n14445 VSS.n230 0.0163425
R8782 VSS.n14445 VSS.n260 0.0163425
R8783 VSS.n14435 VSS.n14424 0.0163425
R8784 VSS.n14435 VSS.n14414 0.0163425
R8785 VSS.n14382 VSS.n413 0.0163425
R8786 VSS.n11783 VSS.n47 0.0163425
R8787 VSS.n11912 VSS.n47 0.0163425
R8788 VSS.n3427 VSS.n47 0.0163425
R8789 VSS.n3349 VSS.n47 0.0163425
R8790 VSS.n3202 VSS.n47 0.0163425
R8791 VSS.n3299 VSS.n3298 0.0161252
R8792 VSS.n5 VSS.n4 0.0161252
R8793 VSS.n8628 VSS 0.016125
R8794 VSS VSS.n8708 0.016125
R8795 VSS.n9703 VSS 0.016125
R8796 VSS VSS.n9115 0.016125
R8797 VSS VSS.n4025 0.016125
R8798 VSS VSS.n7478 0.016125
R8799 VSS.n9427 VSS 0.016125
R8800 VSS.n14363 VSS 0.016125
R8801 VSS.n1077 VSS 0.016125
R8802 VSS.n1327 VSS 0.016125
R8803 VSS VSS.n768 0.016125
R8804 VSS.n13374 VSS 0.016125
R8805 VSS.n13839 VSS 0.016125
R8806 VSS.n1599 VSS 0.016125
R8807 VSS.n319 VSS.n272 0.0157702
R8808 VSS.n14399 VSS.n284 0.0157702
R8809 VSS.n14389 VSS.n370 0.0157702
R8810 VSS.n236 VSS.n169 0.0157702
R8811 VSS.n121 VSS.n112 0.0157702
R8812 VSS.n200 VSS.n184 0.0157702
R8813 VSS.n14443 VSS.n310 0.0157702
R8814 VSS.n205 VSS.n192 0.0157702
R8815 VSS.n216 VSS.n195 0.0157702
R8816 VSS.n311 VSS.n306 0.0157702
R8817 VSS.n386 VSS.n366 0.0157702
R8818 VSS.n398 VSS.n357 0.0157702
R8819 VSS.n438 VSS.n354 0.0157702
R8820 VSS.n429 VSS.n361 0.0157702
R8821 VSS.n14427 VSS.n281 0.0157702
R8822 VSS.n14408 VSS.n288 0.0157702
R8823 VSS.n225 VSS.n188 0.0157702
R8824 VSS.n99 VSS.n88 0.0157702
R8825 VSS.n60 VSS.n51 0.0157702
R8826 VSS.n252 VSS.n163 0.0157702
R8827 VSS.n244 VSS.n160 0.0157702
R8828 VSS.n14417 VSS.n277 0.0157702
R8829 VSS.n407 VSS.n350 0.0157702
R8830 VSS.n419 VSS.n345 0.0157702
R8831 VSS.n77 VSS.n76 0.0157702
R8832 VSS.n101 VSS.n64 0.0157702
R8833 VSS.n127 VSS.n125 0.0157702
R8834 VSS.n140 VSS.n138 0.0157702
R8835 VSS.n3444 VSS.n3399 0.0156042
R8836 VSS.n14435 VSS.n324 0.0155925
R8837 VSS.n14435 VSS.n14404 0.0155925
R8838 VSS.n14383 VSS.n14382 0.0155925
R8839 VSS.n14456 VSS.n113 0.0155925
R8840 VSS.n14456 VSS.n126 0.0155925
R8841 VSS.n14456 VSS.n148 0.0155925
R8842 VSS.n14446 VSS.n14445 0.0155925
R8843 VSS.n14445 VSS.n220 0.0155925
R8844 VSS.n14445 VSS.n210 0.0155925
R8845 VSS.n14436 VSS.n14435 0.0155925
R8846 VSS.n14435 VSS.n333 0.0155925
R8847 VSS.n14382 VSS.n403 0.0155925
R8848 VSS.n14382 VSS.n433 0.0155925
R8849 VSS.n14456 VSS.n100 0.0155925
R8850 VSS.n14456 VSS.n78 0.0155925
R8851 VSS.n14456 VSS.n65 0.0155925
R8852 VSS.n14456 VSS.n52 0.0155925
R8853 VSS.n14445 VSS.n250 0.0155925
R8854 VSS.n14382 VSS.n423 0.0155925
R8855 VSS.n11543 VSS.n47 0.0155925
R8856 VSS.n11768 VSS.n47 0.0155925
R8857 VSS.n14376 VSS.n14375 0.0151004
R8858 VSS.n980 VSS.n979 0.0151004
R8859 VSS.n700 VSS.n699 0.0151004
R8860 VSS.n11502 VSS.n11501 0.0150187
R8861 VSS.n11525 VSS 0.0149369
R8862 VSS.n1501 VSS.n1500 0.0148765
R8863 VSS.n13750 VSS.n13749 0.0148765
R8864 VSS.n13288 VSS.n13287 0.0148765
R8865 VSS.n1238 VSS.n1237 0.0148765
R8866 VSS.n1312 VSS.n1305 0.0146
R8867 VSS.n5245 VSS.n4714 0.0145625
R8868 VSS.n14511 VSS 0.0144825
R8869 VSS.n1062 VSS.n1055 0.0143762
R8870 VSS.n1584 VSS.n1577 0.0141524
R8871 VSS.n14348 VSS.n14341 0.0141524
R8872 VSS.n4534 VSS.n4533 0.0141524
R8873 VSS.n13824 VSS.n13817 0.0141524
R8874 VSS.n13361 VSS.n13354 0.0141524
R8875 VSS.n469 VSS.n454 0.0141524
R8876 VSS.n13420 VSS 0.01413
R8877 VSS.n3419 VSS.n3418 0.0137575
R8878 VSS.n11905 VSS.n11904 0.0137575
R8879 VSS.n3617 VSS.n3616 0.0137575
R8880 VSS.n11489 VSS.n11488 0.0136341
R8881 VSS.n3341 VSS.n3340 0.0135337
R8882 VSS.n11786 VSS.n11785 0.0135337
R8883 VSS.n11535 VSS.n11534 0.0135337
R8884 VSS.n5737 VSS.n5736 0.013521
R8885 VSS.n8634 VSS.n8633 0.0135208
R8886 VSS.n8729 VSS.n8727 0.0135208
R8887 VSS.n9709 VSS.n9708 0.0135208
R8888 VSS.n7500 VSS.n7499 0.0135208
R8889 VSS.n8635 VSS.n8634 0.0133116
R8890 VSS.n8727 VSS.n8726 0.0133116
R8891 VSS.n9710 VSS.n9709 0.0133116
R8892 VSS.n7501 VSS.n7500 0.0133116
R8893 VSS.n10816 VSS.n10815 0.0133116
R8894 VSS.n11761 VSS.n11760 0.0133099
R8895 VSS.n6091 VSS.n6090 0.0132939
R8896 VSS.n5909 VSS.n5908 0.0132939
R8897 VSS.n5728 VSS.n5727 0.0132939
R8898 VSS.n5548 VSS.n5547 0.0132939
R8899 VSS.n5368 VSS.n5367 0.0132939
R8900 VSS.n5188 VSS.n5187 0.0132939
R8901 VSS.n10136 VSS.n10135 0.0132939
R8902 VSS.n11079 VSS.n11078 0.0132939
R8903 VSS.n11994 VSS.n11993 0.0132939
R8904 VSS.n3293 VSS.n3292 0.0132939
R8905 VSS.n12810 VSS.n10 0.0132939
R8906 VSS.n12161 VSS.n12160 0.013121
R8907 VSS.n3 VSS.n1 0.0130333
R8908 VSS.n3199 VSS.n3198 0.0128095
R8909 VSS.n3346 VSS.n3345 0.0128095
R8910 VSS.n11791 VSS.n11790 0.0128095
R8911 VSS.n11540 VSS.n11539 0.0128095
R8912 VSS.n3621 VSS.n3620 0.0128095
R8913 VSS.n11909 VSS.n11908 0.0125857
R8914 VSS.n11765 VSS.n11764 0.0125857
R8915 VSS.n3424 VSS.n3423 0.0123619
R8916 VSS.n3281 VSS.t1 0.0122949
R8917 VSS VSS.n316 0.01225
R8918 VSS.n321 VSS 0.01225
R8919 VSS.n321 VSS 0.01225
R8920 VSS.n14421 VSS 0.01225
R8921 VSS VSS.n14416 0.01225
R8922 VSS.n14416 VSS 0.01225
R8923 VSS VSS.n14398 0.01225
R8924 VSS.n14401 VSS 0.01225
R8925 VSS.n14401 VSS 0.01225
R8926 VSS.n330 VSS 0.01225
R8927 VSS VSS.n327 0.01225
R8928 VSS.n327 VSS 0.01225
R8929 VSS.n410 VSS 0.01225
R8930 VSS VSS.n406 0.01225
R8931 VSS.n406 VSS 0.01225
R8932 VSS VSS.n385 0.01225
R8933 VSS.n390 VSS 0.01225
R8934 VSS.n390 VSS 0.01225
R8935 VSS VSS.n383 0.01225
R8936 VSS VSS.n14388 0.01225
R8937 VSS.n14388 VSS 0.01225
R8938 VSS VSS.n251 0.01225
R8939 VSS.n256 VSS 0.01225
R8940 VSS.n256 VSS 0.01225
R8941 VSS.n237 VSS 0.01225
R8942 VSS VSS.n235 0.01225
R8943 VSS.n235 VSS 0.01225
R8944 VSS VSS.n114 0.01225
R8945 VSS VSS.n120 0.01225
R8946 VSS.n120 VSS 0.01225
R8947 VSS VSS.n128 0.01225
R8948 VSS VSS.n134 0.01225
R8949 VSS.n134 VSS 0.01225
R8950 VSS.n142 VSS 0.01225
R8951 VSS.n144 VSS 0.01225
R8952 VSS VSS.n144 0.01225
R8953 VSS.n14448 VSS 0.01225
R8954 VSS.n14451 VSS 0.01225
R8955 VSS VSS.n14451 0.01225
R8956 VSS VSS.n313 0.01225
R8957 VSS VSS.n14439 0.01225
R8958 VSS.n14439 VSS 0.01225
R8959 VSS VSS.n202 0.01225
R8960 VSS.n207 VSS 0.01225
R8961 VSS.n207 VSS 0.01225
R8962 VSS.n217 VSS 0.01225
R8963 VSS VSS.n213 0.01225
R8964 VSS.n213 VSS 0.01225
R8965 VSS VSS.n395 0.01225
R8966 VSS.n400 VSS 0.01225
R8967 VSS.n400 VSS 0.01225
R8968 VSS VSS.n435 0.01225
R8969 VSS.n440 VSS 0.01225
R8970 VSS.n440 VSS 0.01225
R8971 VSS.n430 VSS 0.01225
R8972 VSS VSS.n426 0.01225
R8973 VSS.n426 VSS 0.01225
R8974 VSS.n14428 VSS 0.01225
R8975 VSS.n14431 VSS 0.01225
R8976 VSS.n14431 VSS 0.01225
R8977 VSS VSS.n14405 0.01225
R8978 VSS.n14411 VSS 0.01225
R8979 VSS.n14411 VSS 0.01225
R8980 VSS VSS.n222 0.01225
R8981 VSS.n227 VSS 0.01225
R8982 VSS.n227 VSS 0.01225
R8983 VSS VSS.n81 0.01225
R8984 VSS VSS.n87 0.01225
R8985 VSS.n87 VSS 0.01225
R8986 VSS VSS.n102 0.01225
R8987 VSS VSS.n108 0.01225
R8988 VSS.n108 VSS 0.01225
R8989 VSS VSS.n53 0.01225
R8990 VSS VSS.n59 0.01225
R8991 VSS.n59 VSS 0.01225
R8992 VSS VSS.n69 0.01225
R8993 VSS VSS.n75 0.01225
R8994 VSS.n75 VSS 0.01225
R8995 VSS VSS.n241 0.01225
R8996 VSS.n246 VSS 0.01225
R8997 VSS.n246 VSS 0.01225
R8998 VSS.n420 VSS 0.01225
R8999 VSS VSS.n416 0.01225
R9000 VSS.n416 VSS 0.01225
R9001 VSS.n8429 VSS.n8416 0.0119583
R9002 VSS.n8625 VSS.n8622 0.0119583
R9003 VSS.n8711 VSS.n8652 0.0119583
R9004 VSS.n9700 VSS.n9697 0.0119583
R9005 VSS.n692 VSS.n691 0.0114223
R9006 VSS.n9356 VSS.n9355 0.0114072
R9007 VSS.n8341 VSS.n8340 0.0114072
R9008 VSS.n8323 VSS.n8322 0.0114072
R9009 VSS.n7518 VSS.n7517 0.0114072
R9010 VSS.n9727 VSS.n9726 0.0114072
R9011 VSS.n3958 VSS.n3957 0.0114072
R9012 VSS.n5738 VSS.n5737 0.0113921
R9013 VSS.n5558 VSS.n5557 0.0113921
R9014 VSS.n5378 VSS.n5377 0.0113921
R9015 VSS.n5198 VSS.n5197 0.0113921
R9016 VSS.n10146 VSS.n10145 0.0113921
R9017 VSS.n11189 VSS.n11186 0.0113921
R9018 VSS.n12361 VSS.n12360 0.0113921
R9019 VSS.n12275 VSS.n12274 0.0113921
R9020 VSS.n11798 VSS.n11797 0.0113921
R9021 VSS.n11815 VSS.n11814 0.0113921
R9022 VSS.n3386 VSS.n3385 0.0113921
R9023 VSS.n3332 VSS.n3331 0.0113921
R9024 VSS.n3300 VSS.n3299 0.0113921
R9025 VSS.n6 VSS.n5 0.0113921
R9026 VSS.n12347 VSS.n12345 0.0112192
R9027 VSS.n11289 VSS.n11277 0.011
R9028 VSS VSS.n11783 0.0105121
R9029 VSS.n11912 VSS 0.0105121
R9030 VSS.n3427 VSS 0.0105121
R9031 VSS.n3349 VSS 0.0105121
R9032 VSS.n3202 VSS 0.0105121
R9033 VSS VSS.n319 0.0105121
R9034 VSS VSS.n14417 0.0105121
R9035 VSS VSS.n14399 0.0105121
R9036 VSS VSS.n310 0.0105121
R9037 VSS VSS.n407 0.0105121
R9038 VSS VSS.n386 0.0105121
R9039 VSS VSS.n14389 0.0105121
R9040 VSS VSS.n252 0.0105121
R9041 VSS VSS.n236 0.0105121
R9042 VSS VSS.n121 0.0105121
R9043 VSS VSS.n127 0.0105121
R9044 VSS VSS.n140 0.0105121
R9045 VSS VSS.n200 0.0105121
R9046 VSS VSS.n311 0.0105121
R9047 VSS VSS.n205 0.0105121
R9048 VSS VSS.n216 0.0105121
R9049 VSS VSS.n398 0.0105121
R9050 VSS VSS.n438 0.0105121
R9051 VSS VSS.n429 0.0105121
R9052 VSS VSS.n14427 0.0105121
R9053 VSS VSS.n14408 0.0105121
R9054 VSS VSS.n225 0.0105121
R9055 VSS.n88 VSS 0.0105121
R9056 VSS VSS.n101 0.0105121
R9057 VSS VSS.n60 0.0105121
R9058 VSS.n76 VSS 0.0105121
R9059 VSS VSS.n244 0.0105121
R9060 VSS VSS.n419 0.0105121
R9061 VSS.n11543 VSS 0.0105121
R9062 VSS.n11768 VSS 0.0105121
R9063 VSS.n323 VSS.n322 0.01037
R9064 VSS.n14403 VSS.n14395 0.01037
R9065 VSS.n14403 VSS.n14402 0.01037
R9066 VSS.n14385 VSS.n14384 0.01037
R9067 VSS.n239 VSS.n231 0.01037
R9068 VSS.n239 VSS.n238 0.01037
R9069 VSS.n119 VSS.n118 0.01037
R9070 VSS.n14449 VSS.n14447 0.01037
R9071 VSS.n332 VSS.n331 0.01037
R9072 VSS.n209 VSS.n208 0.01037
R9073 VSS.n219 VSS.n218 0.01037
R9074 VSS.n14438 VSS.n14437 0.01037
R9075 VSS.n392 VSS.n391 0.01037
R9076 VSS.n402 VSS.n401 0.01037
R9077 VSS.n442 VSS.n441 0.01037
R9078 VSS.n432 VSS.n431 0.01037
R9079 VSS.n14433 VSS.n14432 0.01037
R9080 VSS.n14413 VSS.n14412 0.01037
R9081 VSS.n229 VSS.n228 0.01037
R9082 VSS.n86 VSS.n85 0.01037
R9083 VSS.n85 VSS.n84 0.01037
R9084 VSS.n58 VSS.n57 0.01037
R9085 VSS.n57 VSS.n56 0.01037
R9086 VSS.n259 VSS.n257 0.01037
R9087 VSS.n259 VSS.n258 0.01037
R9088 VSS.n249 VSS.n247 0.01037
R9089 VSS.n249 VSS.n248 0.01037
R9090 VSS.n14423 VSS.n14422 0.01037
R9091 VSS.n412 VSS.n411 0.01037
R9092 VSS.n422 VSS.n421 0.01037
R9093 VSS.n72 VSS.n71 0.01037
R9094 VSS.n72 VSS.n70 0.01037
R9095 VSS.n107 VSS.n106 0.01037
R9096 VSS.n106 VSS.n103 0.01037
R9097 VSS.n133 VSS.n132 0.01037
R9098 VSS.n132 VSS.n129 0.01037
R9099 VSS.n147 VSS.n139 0.01037
R9100 VSS.t0 VSS.n14462 0.0101281
R9101 VSS.n709 VSS.n706 0.0100354
R9102 VSS VSS.n318 0.0100119
R9103 VSS VSS.n320 0.0100119
R9104 VSS VSS.n14419 0.0100119
R9105 VSS VSS.n14415 0.0100119
R9106 VSS VSS.n14397 0.0100119
R9107 VSS VSS.n14400 0.0100119
R9108 VSS VSS.n329 0.0100119
R9109 VSS VSS.n325 0.0100119
R9110 VSS VSS.n409 0.0100119
R9111 VSS VSS.n404 0.0100119
R9112 VSS VSS.n388 0.0100119
R9113 VSS VSS.n389 0.0100119
R9114 VSS VSS.n14342 0.0100119
R9115 VSS VSS.n1056 0.0100119
R9116 VSS VSS.n13818 0.0100119
R9117 VSS VSS.n13355 0.0100119
R9118 VSS.n14390 VSS 0.0100119
R9119 VSS VSS.n14386 0.0100119
R9120 VSS VSS.n254 0.0100119
R9121 VSS VSS.n255 0.0100119
R9122 VSS VSS.n233 0.0100119
R9123 VSS VSS.n234 0.0100119
R9124 VSS.n122 VSS 0.0100119
R9125 VSS.n116 VSS 0.0100119
R9126 VSS.n135 VSS 0.0100119
R9127 VSS.n130 VSS 0.0100119
R9128 VSS VSS.n141 0.0100119
R9129 VSS.n145 VSS 0.0100119
R9130 VSS VSS.n199 0.0100119
R9131 VSS.n14452 VSS 0.0100119
R9132 VSS.n14440 VSS 0.0100119
R9133 VSS VSS.n314 0.0100119
R9134 VSS VSS.n204 0.0100119
R9135 VSS VSS.n206 0.0100119
R9136 VSS VSS.n215 0.0100119
R9137 VSS VSS.n211 0.0100119
R9138 VSS VSS.n397 0.0100119
R9139 VSS VSS.n399 0.0100119
R9140 VSS VSS.n1578 0.0100119
R9141 VSS.n472 VSS 0.0100119
R9142 VSS VSS.n1306 0.0100119
R9143 VSS VSS.n437 0.0100119
R9144 VSS VSS.n439 0.0100119
R9145 VSS VSS.n428 0.0100119
R9146 VSS VSS.n424 0.0100119
R9147 VSS VSS.n14426 0.0100119
R9148 VSS VSS.n14430 0.0100119
R9149 VSS VSS.n14407 0.0100119
R9150 VSS VSS.n14410 0.0100119
R9151 VSS VSS.n224 0.0100119
R9152 VSS VSS.n226 0.0100119
R9153 VSS VSS.n80 0.0100119
R9154 VSS.n82 VSS 0.0100119
R9155 VSS.n109 VSS 0.0100119
R9156 VSS.n104 VSS 0.0100119
R9157 VSS.n61 VSS 0.0100119
R9158 VSS.n54 VSS 0.0100119
R9159 VSS VSS.n68 0.0100119
R9160 VSS VSS.n74 0.0100119
R9161 VSS VSS.n243 0.0100119
R9162 VSS VSS.n245 0.0100119
R9163 VSS VSS.n418 0.0100119
R9164 VSS VSS.n414 0.0100119
R9165 VSS.n4495 VSS.n4494 0.00946062
R9166 VSS.n4509 VSS.n4508 0.00946062
R9167 VSS.n340 VSS.n339 0.00946062
R9168 VSS.n267 VSS.n266 0.00946062
R9169 VSS.n155 VSS.n154 0.00946062
R9170 VSS.n94 VSS.n93 0.00946062
R9171 VSS.n298 VSS.n297 0.00946026
R9172 VSS.n4475 VSS.n4471 0.00946026
R9173 VSS.n4464 VSS.n4461 0.00946026
R9174 VSS.n379 VSS.n375 0.00946026
R9175 VSS.n34 VSS.n33 0.00946026
R9176 VSS.n177 VSS.n176 0.00946026
R9177 VSS.n14459 VSS.n14458 0.00946026
R9178 VSS.n4525 VSS.n4524 0.00922857
R9179 VSS.n3564 VSS.n3396 0.00897165
R9180 VSS.n298 VSS.n296 0.00896
R9181 VSS.n4529 VSS.n4528 0.00896
R9182 VSS.n4464 VSS.n4463 0.00896
R9183 VSS.n4475 VSS.n4474 0.00896
R9184 VSS.n4496 VSS.n4495 0.00896
R9185 VSS.n4510 VSS.n4509 0.00896
R9186 VSS.n4521 VSS.n4520 0.00896
R9187 VSS.n379 VSS.n378 0.00896
R9188 VSS.n34 VSS.n32 0.00896
R9189 VSS.n177 VSS.n175 0.00896
R9190 VSS.n498 VSS.n495 0.00896
R9191 VSS.n341 VSS.n340 0.00896
R9192 VSS.n268 VSS.n267 0.00896
R9193 VSS.n156 VSS.n155 0.00896
R9194 VSS.n95 VSS.n94 0.00896
R9195 VSS.n11929 VSS.n11884 0.00883333
R9196 VSS.n12463 VSS.n12462 0.0083125
R9197 VSS.n10715 VSS.n10714 0.0083125
R9198 VSS.n12267 VSS.n11692 0.00810719
R9199 VSS.n3358 VSS.n3357 0.0079343
R9200 VSS.n5547 VSS.n5546 0.00779167
R9201 VSS.n14343 VSS 0.0076315
R9202 VSS.n14347 VSS 0.0076315
R9203 VSS VSS.n14347 0.0076315
R9204 VSS.n1057 VSS 0.0076315
R9205 VSS.n1061 VSS 0.0076315
R9206 VSS VSS.n1061 0.0076315
R9207 VSS.n13819 VSS 0.0076315
R9208 VSS.n13823 VSS 0.0076315
R9209 VSS VSS.n13823 0.0076315
R9210 VSS.n13356 VSS 0.0076315
R9211 VSS.n13360 VSS 0.0076315
R9212 VSS VSS.n13360 0.0076315
R9213 VSS.n1579 VSS 0.0076315
R9214 VSS.n1583 VSS 0.0076315
R9215 VSS VSS.n1583 0.0076315
R9216 VSS VSS.n452 0.0076315
R9217 VSS VSS.n471 0.0076315
R9218 VSS.n471 VSS 0.0076315
R9219 VSS.n1307 VSS 0.0076315
R9220 VSS.n1311 VSS 0.0076315
R9221 VSS VSS.n1311 0.0076315
R9222 VSS.n9361 VSS.n9360 0.00742521
R9223 VSS.n10794 VSS.n4100 0.007315
R9224 VSS.n10739 VSS.n4535 0.007315
R9225 VSS.n10145 VSS.n10144 0.00727101
R9226 VSS.n9361 VSS.n9358 0.00638643
R9227 VSS.n10818 VSS.n10816 0.00622917
R9228 VSS.n5425 VSS.n4702 0.00622917
R9229 VSS.n293 VSS.n292 0.00610795
R9230 VSS.n293 VSS 0.00610795
R9231 VSS.n300 VSS 0.00610795
R9232 VSS.n300 VSS 0.00610795
R9233 VSS.n4459 VSS.n4458 0.00610795
R9234 VSS.n4459 VSS 0.00610795
R9235 VSS.n4466 VSS 0.00610795
R9236 VSS.n4466 VSS 0.00610795
R9237 VSS.n4477 VSS.n4469 0.00610795
R9238 VSS.n4477 VSS 0.00610795
R9239 VSS.n4472 VSS 0.00610795
R9240 VSS VSS.n4472 0.00610795
R9241 VSS.n4492 VSS.n4491 0.00610795
R9242 VSS.n4492 VSS 0.00610795
R9243 VSS.n4499 VSS 0.00610795
R9244 VSS.n4499 VSS 0.00610795
R9245 VSS.n4506 VSS.n4505 0.00610795
R9246 VSS.n4506 VSS 0.00610795
R9247 VSS.n4513 VSS 0.00610795
R9248 VSS.n4513 VSS 0.00610795
R9249 VSS.n381 VSS.n373 0.00610795
R9250 VSS.n381 VSS 0.00610795
R9251 VSS.n376 VSS 0.00610795
R9252 VSS VSS.n376 0.00610795
R9253 VSS.n36 VSS.n28 0.00610795
R9254 VSS.n36 VSS 0.00610795
R9255 VSS.n30 VSS 0.00610795
R9256 VSS VSS.n30 0.00610795
R9257 VSS.n179 VSS.n171 0.00610795
R9258 VSS.n179 VSS 0.00610795
R9259 VSS.n173 VSS 0.00610795
R9260 VSS VSS.n173 0.00610795
R9261 VSS.n336 VSS.n335 0.00610795
R9262 VSS.n336 VSS 0.00610795
R9263 VSS.n343 VSS 0.00610795
R9264 VSS.n343 VSS 0.00610795
R9265 VSS.n263 VSS.n262 0.00610795
R9266 VSS.n263 VSS 0.00610795
R9267 VSS.n270 VSS 0.00610795
R9268 VSS.n270 VSS 0.00610795
R9269 VSS.n151 VSS.n150 0.00610795
R9270 VSS.n151 VSS 0.00610795
R9271 VSS.n158 VSS 0.00610795
R9272 VSS.n158 VSS 0.00610795
R9273 VSS.n90 VSS.n89 0.00610795
R9274 VSS.n90 VSS 0.00610795
R9275 VSS.n97 VSS 0.00610795
R9276 VSS.n97 VSS 0.00610795
R9277 VSS.n47 VSS.n45 0.00600571
R9278 VSS.n11189 VSS.n11188 0.00585961
R9279 VSS.n3357 VSS.n3356 0.00585961
R9280 VSS.n12268 VSS.n12267 0.00568672
R9281 VSS VSS.n3424 0.00563311
R9282 VSS.n11194 VSS.n11193 0.00557629
R9283 VSS.n11333 VSS.n11332 0.00557629
R9284 VSS VSS.n11909 0.0054727
R9285 VSS VSS.n11765 0.0054727
R9286 VSS.n14435 VSS.n14394 0.0053175
R9287 VSS.n14456 VSS.n14455 0.0053175
R9288 VSS.n14445 VSS.n14444 0.0053175
R9289 VSS.n14382 VSS.n14381 0.0053175
R9290 VSS VSS.n3199 0.00531229
R9291 VSS VSS.n3346 0.00531229
R9292 VSS VSS.n11791 0.00531229
R9293 VSS VSS.n11540 0.00531229
R9294 VSS VSS.n3621 0.00531229
R9295 VSS.n4534 VSS.n4527 0.00526062
R9296 VSS.n240 VSS.n239 0.00523021
R9297 VSS.n393 VSS.n392 0.00523021
R9298 VSS.n443 VSS.n442 0.00523021
R9299 VSS.n14434 VSS.n14433 0.00523021
R9300 VSS.n230 VSS.n229 0.00523021
R9301 VSS.n260 VSS.n259 0.00523021
R9302 VSS.n14424 VSS.n14423 0.00523021
R9303 VSS.n14414 VSS.n14413 0.00523021
R9304 VSS.n413 VSS.n412 0.00523021
R9305 VSS.n11793 VSS.n11783 0.00523021
R9306 VSS.n11913 VSS.n11912 0.00523021
R9307 VSS.n3428 VSS.n3427 0.00523021
R9308 VSS.n3350 VSS.n3349 0.00523021
R9309 VSS.n3203 VSS.n3202 0.00523021
R9310 VSS.n324 VSS.n323 0.00523013
R9311 VSS.n14404 VSS.n14403 0.00523013
R9312 VSS.n14384 VSS.n14383 0.00523013
R9313 VSS.n118 VSS.n113 0.00523013
R9314 VSS.n132 VSS.n126 0.00523013
R9315 VSS.n148 VSS.n147 0.00523013
R9316 VSS.n14447 VSS.n14446 0.00523013
R9317 VSS.n220 VSS.n219 0.00523013
R9318 VSS.n210 VSS.n209 0.00523013
R9319 VSS.n14437 VSS.n14436 0.00523013
R9320 VSS.n333 VSS.n332 0.00523013
R9321 VSS.n403 VSS.n402 0.00523013
R9322 VSS.n433 VSS.n432 0.00523013
R9323 VSS.n106 VSS.n100 0.00523013
R9324 VSS.n85 VSS.n78 0.00523013
R9325 VSS.n72 VSS.n65 0.00523013
R9326 VSS.n57 VSS.n52 0.00523013
R9327 VSS.n250 VSS.n249 0.00523013
R9328 VSS.n423 VSS.n422 0.00523013
R9329 VSS.n11544 VSS.n11543 0.00523013
R9330 VSS.n11769 VSS.n11768 0.00523013
R9331 VSS.n11513 VSS.n11512 0.0052
R9332 VSS.n11512 VSS.n3622 0.0050825
R9333 VSS.n3565 VSS.n3564 0.00482227
R9334 VSS.n4527 VSS.n4526 0.00476029
R9335 VSS.n3343 VSS.n3342 0.00476028
R9336 VSS.n11906 VSS.n11903 0.00476028
R9337 VSS.n11762 VSS.n11759 0.00476028
R9338 VSS.n3618 VSS.n3615 0.00476028
R9339 VSS.n14444 VSS.n291 0.00476028
R9340 VSS.n4518 VSS.n4457 0.00476028
R9341 VSS.n4504 VSS.n4468 0.00476028
R9342 VSS.n4490 VSS.n4479 0.00476028
R9343 VSS.n4486 VSS.n4485 0.00476028
R9344 VSS.n4490 VSS.n4489 0.00476028
R9345 VSS.n4504 VSS.n4503 0.00476028
R9346 VSS.n4518 VSS.n4517 0.00476028
R9347 VSS.n476 VSS.n475 0.00476028
R9348 VSS.n485 VSS.n484 0.00476028
R9349 VSS.n490 VSS.n489 0.00476028
R9350 VSS.n14381 VSS.n488 0.00476028
R9351 VSS.n14394 VSS.n372 0.00476028
R9352 VSS.n14460 VSS.n14457 0.00476028
R9353 VSS.n14455 VSS.n14454 0.00476028
R9354 VSS.n481 VSS.n480 0.00476028
R9355 VSS.n449 VSS.n448 0.00476028
R9356 VSS.n446 VSS.n445 0.00476028
R9357 VSS.n494 VSS.n493 0.00476028
R9358 VSS.n14380 VSS.n14379 0.00476028
R9359 VSS.n14381 VSS.n499 0.00476028
R9360 VSS.n14394 VSS.n348 0.00476028
R9361 VSS.n14444 VSS.n275 0.00476028
R9362 VSS.n14455 VSS.n165 0.00476028
R9363 VSS.n45 VSS.n38 0.00476028
R9364 VSS.n11537 VSS.n11536 0.00476028
R9365 VSS.n11788 VSS.n11787 0.00476028
R9366 VSS.n3421 VSS.n3420 0.00476028
R9367 VSS.n4501 VSS.n4490 0.00473
R9368 VSS.n4515 VSS.n4504 0.00473
R9369 VSS.n4502 VSS.n4501 0.00473
R9370 VSS.n4527 VSS.n4518 0.00473
R9371 VSS.n4516 VSS.n4515 0.00473
R9372 VSS.n1059 VSS.n444 0.00473
R9373 VSS.n13821 VSS.n491 0.00473
R9374 VSS.n13358 VSS.n483 0.00473
R9375 VSS.n14381 VSS.n490 0.00473
R9376 VSS.n14455 VSS.n182 0.00473
R9377 VSS.n14461 VSS.n14456 0.00473
R9378 VSS.n14444 VSS.n303 0.00473
R9379 VSS.n14394 VSS.n14393 0.00473
R9380 VSS.n14444 VSS.n14443 0.00473
R9381 VSS.n14444 VSS.n306 0.00473
R9382 VSS.n14394 VSS.n366 0.00473
R9383 VSS.n14435 VSS.n306 0.00473
R9384 VSS.n14394 VSS.n370 0.00473
R9385 VSS.n14381 VSS.n485 0.00473
R9386 VSS.n14381 VSS.n481 0.00473
R9387 VSS.n14382 VSS.n366 0.00473
R9388 VSS.n1581 VSS.n479 0.00473
R9389 VSS.n1309 VSS.n477 0.00473
R9390 VSS.n473 VSS.n450 0.00473
R9391 VSS.n14381 VSS.n446 0.00473
R9392 VSS.n14381 VSS.n449 0.00473
R9393 VSS.n14394 VSS.n354 0.00473
R9394 VSS.n14394 VSS.n357 0.00473
R9395 VSS.n14444 VSS.n281 0.00473
R9396 VSS.n14444 VSS.n284 0.00473
R9397 VSS.n14455 VSS.n195 0.00473
R9398 VSS.n14456 VSS.n112 0.00473
R9399 VSS.n14455 VSS.n169 0.00473
R9400 VSS.n14456 VSS.n51 0.00473
R9401 VSS.n14444 VSS.n288 0.00473
R9402 VSS.n14444 VSS.n277 0.00473
R9403 VSS.n14445 VSS.n163 0.00473
R9404 VSS.n14394 VSS.n350 0.00473
R9405 VSS.n14394 VSS.n361 0.00473
R9406 VSS.n14381 VSS.n476 0.00473
R9407 VSS.n14381 VSS.n494 0.00473
R9408 VSS.n14345 VSS.n500 0.00473
R9409 VSS.n14381 VSS.n14380 0.00473
R9410 VSS.n14394 VSS.n345 0.00473
R9411 VSS.n14444 VSS.n272 0.00473
R9412 VSS.n14455 VSS.n160 0.00473
R9413 VSS.n14456 VSS.n99 0.00473
R9414 VSS.n85 VSS.n83 0.00473
R9415 VSS.n3618 VSS.n47 0.00473
R9416 VSS.n11537 VSS.n47 0.00473
R9417 VSS.n14455 VSS.n163 0.00473
R9418 VSS.n14456 VSS.n77 0.00473
R9419 VSS.n73 VSS.n72 0.00473
R9420 VSS.n57 VSS.n55 0.00473
R9421 VSS.n11762 VSS.n47 0.00473
R9422 VSS.n11788 VSS.n47 0.00473
R9423 VSS.n14455 VSS.n188 0.00473
R9424 VSS.n14456 VSS.n64 0.00473
R9425 VSS.n106 VSS.n105 0.00473
R9426 VSS.n118 VSS.n117 0.00473
R9427 VSS.n11906 VSS.n47 0.00473
R9428 VSS.n3421 VSS.n47 0.00473
R9429 VSS.n14455 VSS.n192 0.00473
R9430 VSS.n14456 VSS.n125 0.00473
R9431 VSS.n132 VSS.n131 0.00473
R9432 VSS.n3343 VSS.n47 0.00473
R9433 VSS.n14455 VSS.n184 0.00473
R9434 VSS.n14456 VSS.n138 0.00473
R9435 VSS.n147 VSS.n146 0.00473
R9436 VSS.n14461 VSS.n47 0.00473
R9437 VSS.n14461 VSS.n14460 0.00473
R9438 VSS.n14458 VSS.n3 0.00426062
R9439 VSS.n4531 VSS.n4528 0.00426062
R9440 VSS.n4522 VSS.n4521 0.00426062
R9441 VSS.n496 VSS.n495 0.00426062
R9442 VSS.n14461 VSS.n27 0.00426
R9443 VSS.n4028 VSS.n4027 0.00414583
R9444 VSS.n12581 VSS.n12579 0.00414583
R9445 VSS.n3214 VSS.n3212 0.00414583
R9446 VSS.n4481 VSS.n4480 0.00390244
R9447 VSS.n709 VSS.n708 0.00379404
R9448 VSS.n6101 VSS.n6100 0.00378492
R9449 VSS.n5919 VSS.n5918 0.00378492
R9450 VSS.n11336 VSS.n11335 0.00335545
R9451 VSS.n11330 VSS.n11329 0.00335545
R9452 VSS.n11331 VSS.n11330 0.00334133
R9453 VSS.n11335 VSS.n11334 0.00334133
R9454 VSS.n3614 VSS.n3613 0.00327703
R9455 VSS.n4487 VSS.n4486 0.00306417
R9456 VSS.n13308 VSS.n13307 0.00299305
R9457 VSS.n13314 VSS.n13313 0.00299305
R9458 VSS.n13320 VSS.n13319 0.00299305
R9459 VSS.n13324 VSS.n13323 0.00299305
R9460 VSS.n13460 VSS.n13459 0.00299305
R9461 VSS.n13472 VSS.n13471 0.00299305
R9462 VSS.n13474 VSS.n13404 0.00299305
R9463 VSS.n13466 VSS.n13465 0.00299305
R9464 VSS.n13554 VSS.n13512 0.00299305
R9465 VSS.n13517 VSS.n13516 0.00299305
R9466 VSS.n13526 VSS.n13525 0.00299305
R9467 VSS.n13523 VSS.n13520 0.00299305
R9468 VSS.n13594 VSS.n13503 0.00299305
R9469 VSS.n13602 VSS.n13601 0.00299305
R9470 VSS.n13587 VSS.n13501 0.00299305
R9471 VSS.n13508 VSS.n13504 0.00299305
R9472 VSS.n13970 VSS.n13969 0.00299305
R9473 VSS.n13985 VSS.n13984 0.00299305
R9474 VSS.n13982 VSS.n13973 0.00299305
R9475 VSS.n13977 VSS.n13976 0.00299305
R9476 VSS.n14007 VSS.n1738 0.00299305
R9477 VSS.n14015 VSS.n14014 0.00299305
R9478 VSS.n1761 VSS.n1736 0.00299305
R9479 VSS.n1743 VSS.n1739 0.00299305
R9480 VSS.n2979 VSS.n2978 0.00299305
R9481 VSS.n2994 VSS.n2993 0.00299305
R9482 VSS.n2991 VSS.n2982 0.00299305
R9483 VSS.n2986 VSS.n2985 0.00299305
R9484 VSS.n12788 VSS.n12786 0.00299305
R9485 VSS.n12798 VSS.n12797 0.00299305
R9486 VSS.n12784 VSS.n2942 0.00299305
R9487 VSS.n12795 VSS.n12794 0.00299305
R9488 VSS.n2599 VSS.n2593 0.00299305
R9489 VSS.n2637 VSS.n2636 0.00299305
R9490 VSS.n2627 VSS.n2626 0.00299305
R9491 VSS.n2625 VSS.n2624 0.00299305
R9492 VSS.n2617 VSS.n2611 0.00299305
R9493 VSS.n2616 VSS.n2615 0.00299305
R9494 VSS.n2019 VSS.n2013 0.00299305
R9495 VSS.n2030 VSS.n2029 0.00299305
R9496 VSS.n2272 VSS.n2271 0.00299305
R9497 VSS.n2270 VSS.n2269 0.00299305
R9498 VSS.n2262 VSS.n2256 0.00299305
R9499 VSS.n2261 VSS.n2260 0.00299305
R9500 VSS.n1434 VSS.n1433 0.00299305
R9501 VSS.n1428 VSS.n821 0.00299305
R9502 VSS.n1425 VSS.n820 0.00299305
R9503 VSS.n1420 VSS.n819 0.00299305
R9504 VSS.n1619 VSS.n1618 0.00299305
R9505 VSS.n1481 VSS.n1480 0.00299305
R9506 VSS.n1475 VSS.n1474 0.00299305
R9507 VSS.n1469 VSS.n1468 0.00299305
R9508 VSS.n3981 VSS.n3980 0.00299305
R9509 VSS.n3987 VSS.n3986 0.00299305
R9510 VSS.n3993 VSS.n3992 0.00299305
R9511 VSS.n3997 VSS.n3996 0.00299305
R9512 VSS.n4070 VSS.n4069 0.00299305
R9513 VSS.n4082 VSS.n4081 0.00299305
R9514 VSS.n4064 VSS.n4063 0.00299305
R9515 VSS.n4076 VSS.n4075 0.00299305
R9516 VSS.n7335 VSS.n7294 0.00299305
R9517 VSS.n7299 VSS.n7298 0.00299305
R9518 VSS.n7308 VSS.n7307 0.00299305
R9519 VSS.n7305 VSS.n7302 0.00299305
R9520 VSS.n10883 VSS.n10881 0.00299305
R9521 VSS.n10893 VSS.n10892 0.00299305
R9522 VSS.n10879 VSS.n3905 0.00299305
R9523 VSS.n10890 VSS.n10889 0.00299305
R9524 VSS.n3862 VSS.n3861 0.00299305
R9525 VSS.n10989 VSS.n10988 0.00299305
R9526 VSS.n3866 VSS.n3863 0.00299305
R9527 VSS.n3872 VSS.n3871 0.00299305
R9528 VSS.n10929 VSS.n10926 0.00299305
R9529 VSS.n10938 VSS.n10937 0.00299305
R9530 VSS.n10922 VSS.n10918 0.00299305
R9531 VSS.n10935 VSS.n10934 0.00299305
R9532 VSS.n6389 VSS.n6348 0.00299305
R9533 VSS.n6353 VSS.n6352 0.00299305
R9534 VSS.n6362 VSS.n6361 0.00299305
R9535 VSS.n6359 VSS.n6356 0.00299305
R9536 VSS.n11034 VSS.n11032 0.00299305
R9537 VSS.n11044 VSS.n11043 0.00299305
R9538 VSS.n11030 VSS.n3837 0.00299305
R9539 VSS.n11041 VSS.n11040 0.00299305
R9540 VSS.n11137 VSS.n11136 0.00299305
R9541 VSS.n3727 VSS.n3726 0.00299305
R9542 VSS.n3733 VSS.n3732 0.00299305
R9543 VSS.n3737 VSS.n3736 0.00299305
R9544 VSS.n6822 VSS.n6816 0.00299305
R9545 VSS.n6831 VSS.n6792 0.00299305
R9546 VSS.n6842 VSS.n6841 0.00299305
R9547 VSS.n6673 VSS.n6660 0.00299305
R9548 VSS.n6663 VSS.n6662 0.00299305
R9549 VSS.n6667 VSS.n6661 0.00299305
R9550 VSS.n8931 VSS.n8930 0.00299305
R9551 VSS.n8934 VSS.n8933 0.00299305
R9552 VSS.n7887 VSS.n7886 0.00299305
R9553 VSS.n7880 VSS.n7878 0.00299305
R9554 VSS.n9264 VSS.n9263 0.00299305
R9555 VSS.n9258 VSS.n9168 0.00299305
R9556 VSS.n9255 VSS.n9167 0.00299305
R9557 VSS.n9250 VSS.n9166 0.00299305
R9558 VSS.n9447 VSS.n9446 0.00299305
R9559 VSS.n9335 VSS.n9334 0.00299305
R9560 VSS.n9329 VSS.n9328 0.00299305
R9561 VSS.n9323 VSS.n9322 0.00299305
R9562 VSS.n9689 VSS.n9688 0.00299305
R9563 VSS.n9658 VSS.n9657 0.00299305
R9564 VSS.n9652 VSS.n9651 0.00299305
R9565 VSS.n9646 VSS.n9645 0.00299305
R9566 VSS.n9678 VSS.n9674 0.00299305
R9567 VSS.n9672 VSS.n9668 0.00299305
R9568 VSS.n9691 VSS.n9642 0.00299305
R9569 VSS.n9133 VSS.n9132 0.00299305
R9570 VSS.n9127 VSS.n9126 0.00299305
R9571 VSS.n9030 VSS.n9029 0.00299305
R9572 VSS.n9138 VSS.n9020 0.00299305
R9573 VSS.n9046 VSS.n9045 0.00299305
R9574 VSS.n9040 VSS.n9039 0.00299305
R9575 VSS.n9034 VSS.n9033 0.00299305
R9576 VSS.n8825 VSS.n8824 0.00299305
R9577 VSS.n8828 VSS.n8827 0.00299305
R9578 VSS.n8176 VSS.n8175 0.00299305
R9579 VSS.n8169 VSS.n8167 0.00299305
R9580 VSS.n8535 VSS.n8534 0.00299305
R9581 VSS.n8541 VSS.n8540 0.00299305
R9582 VSS.n8547 VSS.n8546 0.00299305
R9583 VSS.n8551 VSS.n8550 0.00299305
R9584 VSS.n8357 VSS.n8353 0.00299305
R9585 VSS.n8363 VSS.n8359 0.00299305
R9586 VSS.n8558 VSS.n8344 0.00299305
R9587 VSS.n8468 VSS.n8467 0.00299305
R9588 VSS.n8483 VSS.n8413 0.00299305
R9589 VSS.n8478 VSS.n8477 0.00299305
R9590 VSS.n8472 VSS.n8471 0.00299305
R9591 VSS.n8505 VSS.n8182 0.00299305
R9592 VSS.n8502 VSS.n8181 0.00299305
R9593 VSS.n8498 VSS.n8180 0.00299305
R9594 VSS.n8492 VSS.n8179 0.00299305
R9595 VSS.n8385 VSS.n8384 0.00299305
R9596 VSS.n8377 VSS.n8368 0.00299305
R9597 VSS.n8375 VSS.n8374 0.00299305
R9598 VSS.n8382 VSS.n8381 0.00299305
R9599 VSS.n8787 VSS.n8786 0.00299305
R9600 VSS.n8790 VSS.n8789 0.00299305
R9601 VSS.n8208 VSS.n8207 0.00299305
R9602 VSS.n8201 VSS.n8199 0.00299305
R9603 VSS.n8404 VSS.n8214 0.00299305
R9604 VSS.n8401 VSS.n8213 0.00299305
R9605 VSS.n8397 VSS.n8212 0.00299305
R9606 VSS.n8391 VSS.n8211 0.00299305
R9607 VSS.n8701 VSS.n8700 0.00299305
R9608 VSS.n8670 VSS.n8669 0.00299305
R9609 VSS.n8664 VSS.n8663 0.00299305
R9610 VSS.n8658 VSS.n8657 0.00299305
R9611 VSS.n8690 VSS.n8686 0.00299305
R9612 VSS.n8684 VSS.n8680 0.00299305
R9613 VSS.n8703 VSS.n8654 0.00299305
R9614 VSS.n9630 VSS.n9629 0.00299305
R9615 VSS.n9635 VSS.n7521 0.00299305
R9616 VSS.n7531 VSS.n7530 0.00299305
R9617 VSS.n9618 VSS.n9617 0.00299305
R9618 VSS.n7547 VSS.n7546 0.00299305
R9619 VSS.n7541 VSS.n7540 0.00299305
R9620 VSS.n7535 VSS.n7534 0.00299305
R9621 VSS.n8750 VSS.n8749 0.00299305
R9622 VSS.n8301 VSS.n8300 0.00299305
R9623 VSS.n8295 VSS.n8294 0.00299305
R9624 VSS.n8289 VSS.n8288 0.00299305
R9625 VSS.n8311 VSS.n8307 0.00299305
R9626 VSS.n8317 VSS.n8313 0.00299305
R9627 VSS.n8738 VSS.n8319 0.00299305
R9628 VSS.n8612 VSS.n8611 0.00299305
R9629 VSS.n8605 VSS.n8604 0.00299305
R9630 VSS.n8599 VSS.n8598 0.00299305
R9631 VSS.n8593 VSS.n8592 0.00299305
R9632 VSS.n8587 VSS.n8586 0.00299305
R9633 VSS.n8581 VSS.n8580 0.00299305
R9634 VSS.n8616 VSS.n8565 0.00299305
R9635 VSS.n8575 VSS.n8574 0.00299305
R9636 VSS.n8255 VSS.n8254 0.00299305
R9637 VSS.n8257 VSS.n8256 0.00299305
R9638 VSS.n8776 VSS.n8775 0.00299305
R9639 VSS.n8241 VSS.n8240 0.00299305
R9640 VSS.n8224 VSS.n8221 0.00299305
R9641 VSS.n8233 VSS.n8232 0.00299305
R9642 VSS.n8227 VSS.n8225 0.00299305
R9643 VSS.n8859 VSS.n8858 0.00299305
R9644 VSS.n8860 VSS.n8005 0.00299305
R9645 VSS.n8867 VSS.n8866 0.00299305
R9646 VSS.n8070 VSS.n8069 0.00299305
R9647 VSS.n8066 VSS.n8065 0.00299305
R9648 VSS.n8059 VSS.n8053 0.00299305
R9649 VSS.n8058 VSS.n8057 0.00299305
R9650 VSS.n9959 VSS.n9953 0.00299305
R9651 VSS.n9967 VSS.n9966 0.00299305
R9652 VSS.n9968 VSS.n6232 0.00299305
R9653 VSS.n9979 VSS.n9978 0.00299305
R9654 VSS.n6217 VSS.n6216 0.00299305
R9655 VSS.n6223 VSS.n6218 0.00299305
R9656 VSS.n6229 VSS.n6228 0.00299305
R9657 VSS.n6189 VSS.n6188 0.00299305
R9658 VSS.n6204 VSS.n4662 0.00299305
R9659 VSS.n6199 VSS.n6198 0.00299305
R9660 VSS.n6747 VSS.n6698 0.00299305
R9661 VSS.n6755 VSS.n6713 0.00299305
R9662 VSS.n6715 VSS.n6714 0.00299305
R9663 VSS.n6751 VSS.n6712 0.00299305
R9664 VSS.n6710 VSS.n6695 0.00299305
R9665 VSS.n6763 VSS.n6762 0.00299305
R9666 VSS.n6709 VSS.n6708 0.00299305
R9667 VSS.n6702 VSS.n6699 0.00299305
R9668 VSS.n8127 VSS.n8126 0.00299305
R9669 VSS.n8143 VSS.n8142 0.00299305
R9670 VSS.n8140 VSS.n8130 0.00299305
R9671 VSS.n8136 VSS.n8135 0.00299305
R9672 VSS.n8153 VSS.n8152 0.00299305
R9673 VSS.n8023 VSS.n8019 0.00299305
R9674 VSS.n8033 VSS.n8022 0.00299305
R9675 VSS.n8024 VSS.n8021 0.00299305
R9676 VSS.n8100 VSS.n8042 0.00299305
R9677 VSS.n8108 VSS.n8093 0.00299305
R9678 VSS.n8095 VSS.n8094 0.00299305
R9679 VSS.n8104 VSS.n8092 0.00299305
R9680 VSS.n8091 VSS.n8040 0.00299305
R9681 VSS.n8046 VSS.n8045 0.00299305
R9682 VSS.n8083 VSS.n8044 0.00299305
R9683 VSS.n8079 VSS.n8043 0.00299305
R9684 VSS.n8879 VSS.n7955 0.00299305
R9685 VSS.n8887 VSS.n7970 0.00299305
R9686 VSS.n7972 VSS.n7971 0.00299305
R9687 VSS.n8883 VSS.n7969 0.00299305
R9688 VSS.n7967 VSS.n7951 0.00299305
R9689 VSS.n8895 VSS.n8894 0.00299305
R9690 VSS.n7966 VSS.n7965 0.00299305
R9691 VSS.n7959 VSS.n7956 0.00299305
R9692 VSS.n8815 VSS.n8814 0.00299305
R9693 VSS.n8798 VSS.n8191 0.00299305
R9694 VSS.n8806 VSS.n8805 0.00299305
R9695 VSS.n8800 VSS.n8799 0.00299305
R9696 VSS.n9553 VSS.n9552 0.00299305
R9697 VSS.n7575 VSS.n7572 0.00299305
R9698 VSS.n7584 VSS.n7583 0.00299305
R9699 VSS.n7581 VSS.n7580 0.00299305
R9700 VSS.n8271 VSS.n8270 0.00299305
R9701 VSS.n8273 VSS.n8264 0.00299305
R9702 VSS.n8278 VSS.n8277 0.00299305
R9703 VSS.n8281 VSS.n8280 0.00299305
R9704 VSS.n9589 VSS.n9588 0.00299305
R9705 VSS.n9592 VSS.n9591 0.00299305
R9706 VSS.n9560 VSS.n7559 0.00299305
R9707 VSS.n9566 VSS.n7560 0.00299305
R9708 VSS.n9568 VSS.n7561 0.00299305
R9709 VSS.n9576 VSS.n9575 0.00299305
R9710 VSS.n9582 VSS.n9581 0.00299305
R9711 VSS.n8445 VSS.n8444 0.00299305
R9712 VSS.n8440 VSS.n8439 0.00299305
R9713 VSS.n8455 VSS.n8454 0.00299305
R9714 VSS.n9412 VSS.n9411 0.00299305
R9715 VSS.n9405 VSS.n9404 0.00299305
R9716 VSS.n9399 VSS.n9398 0.00299305
R9717 VSS.n9393 VSS.n9392 0.00299305
R9718 VSS.n9387 VSS.n9386 0.00299305
R9719 VSS.n9381 VSS.n9380 0.00299305
R9720 VSS.n9416 VSS.n9365 0.00299305
R9721 VSS.n9375 VSS.n9374 0.00299305
R9722 VSS.n7418 VSS.n7417 0.00299305
R9723 VSS.n9782 VSS.n9781 0.00299305
R9724 VSS.n9788 VSS.n9787 0.00299305
R9725 VSS.n7402 VSS.n7401 0.00299305
R9726 VSS.n7408 VSS.n7407 0.00299305
R9727 VSS.n7412 VSS.n7411 0.00299305
R9728 VSS.n7388 VSS.n7384 0.00299305
R9729 VSS.n7469 VSS.n7468 0.00299305
R9730 VSS.n7462 VSS.n7461 0.00299305
R9731 VSS.n7456 VSS.n7455 0.00299305
R9732 VSS.n7450 VSS.n7449 0.00299305
R9733 VSS.n7444 VSS.n7443 0.00299305
R9734 VSS.n7438 VSS.n7437 0.00299305
R9735 VSS.n7473 VSS.n7422 0.00299305
R9736 VSS.n7432 VSS.n7431 0.00299305
R9737 VSS.n3954 VSS.n3953 0.00299305
R9738 VSS.n10829 VSS.n10828 0.00299305
R9739 VSS.n10835 VSS.n10834 0.00299305
R9740 VSS.n3938 VSS.n3937 0.00299305
R9741 VSS.n3944 VSS.n3943 0.00299305
R9742 VSS.n3948 VSS.n3947 0.00299305
R9743 VSS.n3924 VSS.n3920 0.00299305
R9744 VSS.n9345 VSS.n9341 0.00299305
R9745 VSS.n9351 VSS.n9347 0.00299305
R9746 VSS.n9435 VSS.n9353 0.00299305
R9747 VSS.n9106 VSS.n9105 0.00299305
R9748 VSS.n9099 VSS.n9098 0.00299305
R9749 VSS.n9093 VSS.n9092 0.00299305
R9750 VSS.n9087 VSS.n9086 0.00299305
R9751 VSS.n9081 VSS.n9080 0.00299305
R9752 VSS.n9075 VSS.n9074 0.00299305
R9753 VSS.n9110 VSS.n9059 0.00299305
R9754 VSS.n9069 VSS.n9068 0.00299305
R9755 VSS.n9514 VSS.n9015 0.00299305
R9756 VSS.n9518 VSS.n9517 0.00299305
R9757 VSS.n9014 VSS.n9013 0.00299305
R9758 VSS.n9007 VSS.n9005 0.00299305
R9759 VSS.n9274 VSS.n9003 0.00299305
R9760 VSS.n9276 VSS.n9002 0.00299305
R9761 VSS.n9283 VSS.n9001 0.00299305
R9762 VSS.n9285 VSS.n9000 0.00299305
R9763 VSS.n9502 VSS.n9501 0.00299305
R9764 VSS.n9505 VSS.n9504 0.00299305
R9765 VSS.n9313 VSS.n9292 0.00299305
R9766 VSS.n9309 VSS.n9308 0.00299305
R9767 VSS.n9301 VSS.n9295 0.00299305
R9768 VSS.n9300 VSS.n9299 0.00299305
R9769 VSS.n9494 VSS.n9493 0.00299305
R9770 VSS.n9817 VSS.n9811 0.00299305
R9771 VSS.n9825 VSS.n9824 0.00299305
R9772 VSS.n9827 VSS.n9826 0.00299305
R9773 VSS.n7227 VSS.n7226 0.00299305
R9774 VSS.n7233 VSS.n7232 0.00299305
R9775 VSS.n7236 VSS.n7235 0.00299305
R9776 VSS.n9836 VSS.n7179 0.00299305
R9777 VSS.n9840 VSS.n9839 0.00299305
R9778 VSS.n7178 VSS.n7177 0.00299305
R9779 VSS.n7171 VSS.n7169 0.00299305
R9780 VSS.n9471 VSS.n7167 0.00299305
R9781 VSS.n9475 VSS.n7166 0.00299305
R9782 VSS.n9482 VSS.n7165 0.00299305
R9783 VSS.n9479 VSS.n7164 0.00299305
R9784 VSS.n7376 VSS.n7193 0.00299305
R9785 VSS.n7258 VSS.n7257 0.00299305
R9786 VSS.n7213 VSS.n7212 0.00299305
R9787 VSS.n7248 VSS.n7247 0.00299305
R9788 VSS.n7246 VSS.n7245 0.00299305
R9789 VSS.n7276 VSS.n7267 0.00299305
R9790 VSS.n7275 VSS.n7274 0.00299305
R9791 VSS.n7359 VSS.n7273 0.00299305
R9792 VSS.n7321 VSS.n7268 0.00299305
R9793 VSS.n7317 VSS.n7270 0.00299305
R9794 VSS.n7271 VSS.n7265 0.00299305
R9795 VSS.n7325 VSS.n7269 0.00299305
R9796 VSS.n7197 VSS.n7195 0.00299305
R9797 VSS.n7207 VSS.n7196 0.00299305
R9798 VSS.n9171 VSS.n9170 0.00299305
R9799 VSS.n9181 VSS.n9163 0.00299305
R9800 VSS.n9266 VSS.n9164 0.00299305
R9801 VSS.n9239 VSS.n9238 0.00299305
R9802 VSS.n9219 VSS.n9216 0.00299305
R9803 VSS.n9228 VSS.n9227 0.00299305
R9804 VSS.n9225 VSS.n9224 0.00299305
R9805 VSS.n9194 VSS.n9193 0.00299305
R9806 VSS.n9202 VSS.n9201 0.00299305
R9807 VSS.n9205 VSS.n9204 0.00299305
R9808 VSS.n9211 VSS.n9210 0.00299305
R9809 VSS.n7839 VSS.n7816 0.00299305
R9810 VSS.n7842 VSS.n7817 0.00299305
R9811 VSS.n8957 VSS.n8956 0.00299305
R9812 VSS.n7826 VSS.n7812 0.00299305
R9813 VSS.n7825 VSS.n7824 0.00299305
R9814 VSS.n8959 VSS.n7813 0.00299305
R9815 VSS.n8946 VSS.n8945 0.00299305
R9816 VSS.n7858 VSS.n7855 0.00299305
R9817 VSS.n7867 VSS.n7866 0.00299305
R9818 VSS.n7864 VSS.n7863 0.00299305
R9819 VSS.n7900 VSS.n7897 0.00299305
R9820 VSS.n7905 VSS.n7904 0.00299305
R9821 VSS.n7914 VSS.n7913 0.00299305
R9822 VSS.n7911 VSS.n7910 0.00299305
R9823 VSS.n7790 VSS.n7784 0.00299305
R9824 VSS.n7798 VSS.n7797 0.00299305
R9825 VSS.n7800 VSS.n7799 0.00299305
R9826 VSS.n7740 VSS.n7739 0.00299305
R9827 VSS.n7746 VSS.n7745 0.00299305
R9828 VSS.n7749 VSS.n7748 0.00299305
R9829 VSS.n7633 VSS.n7630 0.00299305
R9830 VSS.n8979 VSS.n7629 0.00299305
R9831 VSS.n8969 VSS.n7628 0.00299305
R9832 VSS.n8973 VSS.n7627 0.00299305
R9833 VSS.n7620 VSS.n7619 0.00299305
R9834 VSS.n7621 VSS.n7618 0.00299305
R9835 VSS.n8987 VSS.n8986 0.00299305
R9836 VSS.n7634 VSS.n7617 0.00299305
R9837 VSS.n7711 VSS.n7705 0.00299305
R9838 VSS.n7719 VSS.n7718 0.00299305
R9839 VSS.n7721 VSS.n7720 0.00299305
R9840 VSS.n7692 VSS.n7678 0.00299305
R9841 VSS.n7683 VSS.n7682 0.00299305
R9842 VSS.n7690 VSS.n7689 0.00299305
R9843 VSS.n7668 VSS.n7665 0.00299305
R9844 VSS.n7769 VSS.n7664 0.00299305
R9845 VSS.n7759 VSS.n7663 0.00299305
R9846 VSS.n7763 VSS.n7662 0.00299305
R9847 VSS.n7655 VSS.n7654 0.00299305
R9848 VSS.n7656 VSS.n7653 0.00299305
R9849 VSS.n7777 VSS.n7776 0.00299305
R9850 VSS.n7669 VSS.n7652 0.00299305
R9851 VSS.n9883 VSS.n7143 0.00299305
R9852 VSS.n9894 VSS.n9893 0.00299305
R9853 VSS.n7074 VSS.n7073 0.00299305
R9854 VSS.n7080 VSS.n7075 0.00299305
R9855 VSS.n7086 VSS.n7085 0.00299305
R9856 VSS.n7120 VSS.n7094 0.00299305
R9857 VSS.n7119 VSS.n7118 0.00299305
R9858 VSS.n7129 VSS.n7117 0.00299305
R9859 VSS.n7103 VSS.n7095 0.00299305
R9860 VSS.n7098 VSS.n7097 0.00299305
R9861 VSS.n7115 VSS.n7092 0.00299305
R9862 VSS.n7108 VSS.n7096 0.00299305
R9863 VSS.n9874 VSS.n9868 0.00299305
R9864 VSS.n9882 VSS.n9881 0.00299305
R9865 VSS.n7929 VSS.n7889 0.00299305
R9866 VSS.n7933 VSS.n7890 0.00299305
R9867 VSS.n7937 VSS.n7891 0.00299305
R9868 VSS.n8921 VSS.n8920 0.00299305
R9869 VSS.n8904 VSS.n7945 0.00299305
R9870 VSS.n8912 VSS.n8911 0.00299305
R9871 VSS.n8906 VSS.n8905 0.00299305
R9872 VSS.n7995 VSS.n7994 0.00299305
R9873 VSS.n7992 VSS.n7991 0.00299305
R9874 VSS.n7981 VSS.n7979 0.00299305
R9875 VSS.n6853 VSS.n6632 0.00299305
R9876 VSS.n6642 VSS.n6641 0.00299305
R9877 VSS.n6652 VSS.n6640 0.00299305
R9878 VSS.n6649 VSS.n6639 0.00299305
R9879 VSS.n6797 VSS.n6637 0.00299305
R9880 VSS.n6801 VSS.n6636 0.00299305
R9881 VSS.n6808 VSS.n6635 0.00299305
R9882 VSS.n6805 VSS.n6634 0.00299305
R9883 VSS.n6889 VSS.n6883 0.00299305
R9884 VSS.n6909 VSS.n6908 0.00299305
R9885 VSS.n6625 VSS.n6612 0.00299305
R9886 VSS.n6615 VSS.n6614 0.00299305
R9887 VSS.n6619 VSS.n6613 0.00299305
R9888 VSS.n6899 VSS.n6898 0.00299305
R9889 VSS.n6897 VSS.n6896 0.00299305
R9890 VSS.n6920 VSS.n6584 0.00299305
R9891 VSS.n6594 VSS.n6593 0.00299305
R9892 VSS.n6604 VSS.n6592 0.00299305
R9893 VSS.n6601 VSS.n6591 0.00299305
R9894 VSS.n6865 VSS.n6589 0.00299305
R9895 VSS.n6869 VSS.n6588 0.00299305
R9896 VSS.n6876 VSS.n6587 0.00299305
R9897 VSS.n6873 VSS.n6586 0.00299305
R9898 VSS.n6962 VSS.n6956 0.00299305
R9899 VSS.n6982 VSS.n6981 0.00299305
R9900 VSS.n6577 VSS.n6564 0.00299305
R9901 VSS.n6567 VSS.n6566 0.00299305
R9902 VSS.n6571 VSS.n6565 0.00299305
R9903 VSS.n6972 VSS.n6971 0.00299305
R9904 VSS.n6970 VSS.n6969 0.00299305
R9905 VSS.n7010 VSS.n6518 0.00299305
R9906 VSS.n7008 VSS.n6519 0.00299305
R9907 VSS.n7039 VSS.n7038 0.00299305
R9908 VSS.n6528 VSS.n6514 0.00299305
R9909 VSS.n6527 VSS.n6526 0.00299305
R9910 VSS.n7041 VSS.n6515 0.00299305
R9911 VSS.n6994 VSS.n6993 0.00299305
R9912 VSS.n6547 VSS.n6544 0.00299305
R9913 VSS.n6556 VSS.n6555 0.00299305
R9914 VSS.n6553 VSS.n6552 0.00299305
R9915 VSS.n6935 VSS.n6932 0.00299305
R9916 VSS.n6940 VSS.n6939 0.00299305
R9917 VSS.n6949 VSS.n6948 0.00299305
R9918 VSS.n6946 VSS.n6945 0.00299305
R9919 VSS.n6277 VSS.n6276 0.00299305
R9920 VSS.n6288 VSS.n6287 0.00299305
R9921 VSS.n7062 VSS.n6274 0.00299305
R9922 VSS.n6477 VSS.n6476 0.00299305
R9923 VSS.n6469 VSS.n6468 0.00299305
R9924 VSS.n6466 VSS.n6465 0.00299305
R9925 VSS.n7052 VSS.n6486 0.00299305
R9926 VSS.n6496 VSS.n6495 0.00299305
R9927 VSS.n6506 VSS.n6494 0.00299305
R9928 VSS.n6503 VSS.n6493 0.00299305
R9929 VSS.n7018 VSS.n6491 0.00299305
R9930 VSS.n7022 VSS.n6490 0.00299305
R9931 VSS.n7029 VSS.n6489 0.00299305
R9932 VSS.n7026 VSS.n6488 0.00299305
R9933 VSS.n6445 VSS.n6427 0.00299305
R9934 VSS.n6456 VSS.n6455 0.00299305
R9935 VSS.n6301 VSS.n6300 0.00299305
R9936 VSS.n6307 VSS.n6302 0.00299305
R9937 VSS.n6313 VSS.n6312 0.00299305
R9938 VSS.n6330 VSS.n6321 0.00299305
R9939 VSS.n6329 VSS.n6328 0.00299305
R9940 VSS.n6413 VSS.n6327 0.00299305
R9941 VSS.n6375 VSS.n6322 0.00299305
R9942 VSS.n6371 VSS.n6324 0.00299305
R9943 VSS.n6325 VSS.n6319 0.00299305
R9944 VSS.n6379 VSS.n6323 0.00299305
R9945 VSS.n6436 VSS.n6430 0.00299305
R9946 VSS.n6444 VSS.n6443 0.00299305
R9947 VSS.n6830 VSS.n6829 0.00299305
R9948 VSS.n6785 VSS.n6679 0.00299305
R9949 VSS.n6688 VSS.n6687 0.00299305
R9950 VSS.n6777 VSS.n6686 0.00299305
R9951 VSS.n6773 VSS.n6685 0.00299305
R9952 VSS.n6731 VSS.n6683 0.00299305
R9953 VSS.n6733 VSS.n6682 0.00299305
R9954 VSS.n6727 VSS.n6681 0.00299305
R9955 VSS.n6039 VSS.n6038 0.00299305
R9956 VSS.n6032 VSS.n6031 0.00299305
R9957 VSS.n6026 VSS.n6025 0.00299305
R9958 VSS.n6020 VSS.n6019 0.00299305
R9959 VSS.n6014 VSS.n6013 0.00299305
R9960 VSS.n6008 VSS.n6007 0.00299305
R9961 VSS.n6043 VSS.n5992 0.00299305
R9962 VSS.n6002 VSS.n6001 0.00299305
R9963 VSS.n5866 VSS.n5865 0.00299305
R9964 VSS.n5898 VSS.n5897 0.00299305
R9965 VSS.n5882 VSS.n5881 0.00299305
R9966 VSS.n5876 VSS.n5875 0.00299305
R9967 VSS.n5870 VSS.n5869 0.00299305
R9968 VSS.n5854 VSS.n5791 0.00299305
R9969 VSS.n5860 VSS.n5856 0.00299305
R9970 VSS.n5841 VSS.n5840 0.00299305
R9971 VSS.n5834 VSS.n5833 0.00299305
R9972 VSS.n5828 VSS.n5827 0.00299305
R9973 VSS.n5822 VSS.n5821 0.00299305
R9974 VSS.n5816 VSS.n5815 0.00299305
R9975 VSS.n5810 VSS.n5809 0.00299305
R9976 VSS.n5845 VSS.n5794 0.00299305
R9977 VSS.n5804 VSS.n5803 0.00299305
R9978 VSS.n5685 VSS.n5684 0.00299305
R9979 VSS.n5717 VSS.n5716 0.00299305
R9980 VSS.n5701 VSS.n5700 0.00299305
R9981 VSS.n5695 VSS.n5694 0.00299305
R9982 VSS.n5689 VSS.n5688 0.00299305
R9983 VSS.n5673 VSS.n5610 0.00299305
R9984 VSS.n5679 VSS.n5675 0.00299305
R9985 VSS.n5660 VSS.n5659 0.00299305
R9986 VSS.n5653 VSS.n5652 0.00299305
R9987 VSS.n5647 VSS.n5646 0.00299305
R9988 VSS.n5641 VSS.n5640 0.00299305
R9989 VSS.n5635 VSS.n5634 0.00299305
R9990 VSS.n5629 VSS.n5628 0.00299305
R9991 VSS.n5664 VSS.n5613 0.00299305
R9992 VSS.n5623 VSS.n5622 0.00299305
R9993 VSS.n5505 VSS.n5504 0.00299305
R9994 VSS.n5537 VSS.n5536 0.00299305
R9995 VSS.n5521 VSS.n5520 0.00299305
R9996 VSS.n5515 VSS.n5514 0.00299305
R9997 VSS.n5509 VSS.n5508 0.00299305
R9998 VSS.n5493 VSS.n5430 0.00299305
R9999 VSS.n5499 VSS.n5495 0.00299305
R10000 VSS.n5480 VSS.n5479 0.00299305
R10001 VSS.n5473 VSS.n5472 0.00299305
R10002 VSS.n5467 VSS.n5466 0.00299305
R10003 VSS.n5461 VSS.n5460 0.00299305
R10004 VSS.n5455 VSS.n5454 0.00299305
R10005 VSS.n5449 VSS.n5448 0.00299305
R10006 VSS.n5484 VSS.n5433 0.00299305
R10007 VSS.n5443 VSS.n5442 0.00299305
R10008 VSS.n5325 VSS.n5324 0.00299305
R10009 VSS.n5357 VSS.n5356 0.00299305
R10010 VSS.n5341 VSS.n5340 0.00299305
R10011 VSS.n5335 VSS.n5334 0.00299305
R10012 VSS.n5329 VSS.n5328 0.00299305
R10013 VSS.n5313 VSS.n5250 0.00299305
R10014 VSS.n5319 VSS.n5315 0.00299305
R10015 VSS.n5300 VSS.n5299 0.00299305
R10016 VSS.n5293 VSS.n5292 0.00299305
R10017 VSS.n5287 VSS.n5286 0.00299305
R10018 VSS.n5281 VSS.n5280 0.00299305
R10019 VSS.n5275 VSS.n5274 0.00299305
R10020 VSS.n5269 VSS.n5268 0.00299305
R10021 VSS.n5304 VSS.n5253 0.00299305
R10022 VSS.n5263 VSS.n5262 0.00299305
R10023 VSS.n10059 VSS.n10058 0.00299305
R10024 VSS.n10091 VSS.n10090 0.00299305
R10025 VSS.n10075 VSS.n10074 0.00299305
R10026 VSS.n10069 VSS.n10068 0.00299305
R10027 VSS.n10063 VSS.n10062 0.00299305
R10028 VSS.n10047 VSS.n4577 0.00299305
R10029 VSS.n10053 VSS.n10049 0.00299305
R10030 VSS.n4627 VSS.n4626 0.00299305
R10031 VSS.n4586 VSS.n4585 0.00299305
R10032 VSS.n4592 VSS.n4591 0.00299305
R10033 VSS.n4598 VSS.n4597 0.00299305
R10034 VSS.n4602 VSS.n4601 0.00299305
R10035 VSS.n3765 VSS.n3764 0.00299305
R10036 VSS.n3808 VSS.n3807 0.00299305
R10037 VSS.n3802 VSS.n3801 0.00299305
R10038 VSS.n3769 VSS.n3768 0.00299305
R10039 VSS.n3781 VSS.n3780 0.00299305
R10040 VSS.n3790 VSS.n3789 0.00299305
R10041 VSS.n3775 VSS.n3774 0.00299305
R10042 VSS.n4617 VSS.n4613 0.00299305
R10043 VSS.n4623 VSS.n4619 0.00299305
R10044 VSS.n6061 VSS.n6060 0.00299305
R10045 VSS.n6055 VSS.n6054 0.00299305
R10046 VSS.n6072 VSS.n6071 0.00299305
R10047 VSS.n6067 VSS.n6063 0.00299305
R10048 VSS.n6080 VSS.n5972 0.00299305
R10049 VSS.n5986 VSS.n5982 0.00299305
R10050 VSS.n5980 VSS.n5976 0.00299305
R10051 VSS.n6166 VSS.n6165 0.00299305
R10052 VSS.n6161 VSS.n6160 0.00299305
R10053 VSS.n6176 VSS.n6175 0.00299305
R10054 VSS.n6170 VSS.n6169 0.00299305
R10055 VSS.n11094 VSS.n11093 0.00299305
R10056 VSS.n11106 VSS.n11105 0.00299305
R10057 VSS.n11088 VSS.n11087 0.00299305
R10058 VSS.n11100 VSS.n11099 0.00299305
R10059 VSS.n3747 VSS.n3743 0.00299305
R10060 VSS.n3753 VSS.n3749 0.00299305
R10061 VSS.n11130 VSS.n3755 0.00299305
R10062 VSS.n11056 VSS.n11055 0.00299305
R10063 VSS.n11108 VSS.n11051 0.00299305
R10064 VSS.n11066 VSS.n11065 0.00299305
R10065 VSS.n6343 VSS.n6342 0.00299305
R10066 VSS.n6401 VSS.n6400 0.00299305
R10067 VSS.n6398 VSS.n6397 0.00299305
R10068 VSS.n11021 VSS.n3831 0.00299305
R10069 VSS.n11019 VSS.n3832 0.00299305
R10070 VSS.n11009 VSS.n3834 0.00299305
R10071 VSS.n10969 VSS.n3874 0.00299305
R10072 VSS.n10980 VSS.n3875 0.00299305
R10073 VSS.n3878 VSS.n3876 0.00299305
R10074 VSS.n10949 VSS.n10948 0.00299305
R10075 VSS.n10915 VSS.n10914 0.00299305
R10076 VSS.n10908 VSS.n10902 0.00299305
R10077 VSS.n7289 VSS.n7288 0.00299305
R10078 VSS.n7347 VSS.n7346 0.00299305
R10079 VSS.n7344 VSS.n7343 0.00299305
R10080 VSS.n10870 VSS.n3899 0.00299305
R10081 VSS.n10868 VSS.n3900 0.00299305
R10082 VSS.n10858 VSS.n3902 0.00299305
R10083 VSS.n4007 VSS.n4003 0.00299305
R10084 VSS.n4013 VSS.n4009 0.00299305
R10085 VSS.n4020 VSS.n3971 0.00299305
R10086 VSS.n4039 VSS.n4038 0.00299305
R10087 VSS.n4084 VSS.n4034 0.00299305
R10088 VSS.n4049 VSS.n4048 0.00299305
R10089 VSS.n4416 VSS.n4115 0.00299305
R10090 VSS.n4429 VSS.n4116 0.00299305
R10091 VSS.n4426 VSS.n4117 0.00299305
R10092 VSS.n4421 VSS.n4118 0.00299305
R10093 VSS.n4393 VSS.n4191 0.00299305
R10094 VSS.n4397 VSS.n4192 0.00299305
R10095 VSS.n4198 VSS.n4193 0.00299305
R10096 VSS.n4221 VSS.n4194 0.00299305
R10097 VSS.n4215 VSS.n4189 0.00299305
R10098 VSS.n4142 VSS.n4141 0.00299305
R10099 VSS.n4140 VSS.n4136 0.00299305
R10100 VSS.n4448 VSS.n4447 0.00299305
R10101 VSS.n4148 VSS.n4147 0.00299305
R10102 VSS.n4361 VSS.n4183 0.00299305
R10103 VSS.n4373 VSS.n4182 0.00299305
R10104 VSS.n4363 VSS.n4185 0.00299305
R10105 VSS.n4367 VSS.n4184 0.00299305
R10106 VSS.n4305 VSS.n4304 0.00299305
R10107 VSS.n4320 VSS.n4319 0.00299305
R10108 VSS.n4317 VSS.n4308 0.00299305
R10109 VSS.n4312 VSS.n4311 0.00299305
R10110 VSS.n4335 VSS.n4252 0.00299305
R10111 VSS.n4343 VSS.n4342 0.00299305
R10112 VSS.n4264 VSS.n4250 0.00299305
R10113 VSS.n4257 VSS.n4253 0.00299305
R10114 VSS.n4285 VSS.n4279 0.00299305
R10115 VSS.n4293 VSS.n4292 0.00299305
R10116 VSS.n4294 VSS.n4272 0.00299305
R10117 VSS.n4346 VSS.n4345 0.00299305
R10118 VSS.n4239 VSS.n4235 0.00299305
R10119 VSS.n4238 VSS.n4237 0.00299305
R10120 VSS.n4219 VSS.n4196 0.00299305
R10121 VSS.n4169 VSS.n4168 0.00299305
R10122 VSS.n4175 VSS.n4167 0.00299305
R10123 VSS.n4172 VSS.n4166 0.00299305
R10124 VSS.n4407 VSS.n4406 0.00299305
R10125 VSS.n4126 VSS.n4120 0.00299305
R10126 VSS.n10778 VSS.n10777 0.00299305
R10127 VSS.n4129 VSS.n4127 0.00299305
R10128 VSS.n10766 VSS.n10765 0.00299305
R10129 VSS.n10764 VSS.n10763 0.00299305
R10130 VSS.n10756 VSS.n10750 0.00299305
R10131 VSS.n1295 VSS.n1294 0.00299305
R10132 VSS.n1264 VSS.n1263 0.00299305
R10133 VSS.n1258 VSS.n1257 0.00299305
R10134 VSS.n1252 VSS.n1251 0.00299305
R10135 VSS.n1284 VSS.n1280 0.00299305
R10136 VSS.n1278 VSS.n1274 0.00299305
R10137 VSS.n1297 VSS.n1248 0.00299305
R10138 VSS.n786 VSS.n785 0.00299305
R10139 VSS.n780 VSS.n779 0.00299305
R10140 VSS.n664 VSS.n663 0.00299305
R10141 VSS.n791 VSS.n654 0.00299305
R10142 VSS.n680 VSS.n679 0.00299305
R10143 VSS.n674 VSS.n673 0.00299305
R10144 VSS.n668 VSS.n667 0.00299305
R10145 VSS.n1348 VSS.n1347 0.00299305
R10146 VSS.n1212 VSS.n1211 0.00299305
R10147 VSS.n1206 VSS.n1205 0.00299305
R10148 VSS.n1200 VSS.n1199 0.00299305
R10149 VSS.n1222 VSS.n1218 0.00299305
R10150 VSS.n1228 VSS.n1224 0.00299305
R10151 VSS.n1336 VSS.n1230 0.00299305
R10152 VSS.n1044 VSS.n1043 0.00299305
R10153 VSS.n1037 VSS.n1036 0.00299305
R10154 VSS.n1031 VSS.n1030 0.00299305
R10155 VSS.n1025 VSS.n1024 0.00299305
R10156 VSS.n1019 VSS.n1018 0.00299305
R10157 VSS.n1013 VSS.n1012 0.00299305
R10158 VSS.n1048 VSS.n997 0.00299305
R10159 VSS.n1007 VSS.n1006 0.00299305
R10160 VSS.n14177 VSS.n14176 0.00299305
R10161 VSS.n14193 VSS.n14192 0.00299305
R10162 VSS.n14190 VSS.n14180 0.00299305
R10163 VSS.n14186 VSS.n14185 0.00299305
R10164 VSS.n1109 VSS.n1108 0.00299305
R10165 VSS.n1092 VSS.n1091 0.00299305
R10166 VSS.n1098 VSS.n1097 0.00299305
R10167 VSS.n1102 VSS.n1101 0.00299305
R10168 VSS.n970 VSS.n966 0.00299305
R10169 VSS.n976 VSS.n972 0.00299305
R10170 VSS.n1086 VSS.n978 0.00299305
R10171 VSS.n14318 VSS.n14317 0.00299305
R10172 VSS.n14313 VSS.n14312 0.00299305
R10173 VSS.n14328 VSS.n14327 0.00299305
R10174 VSS.n14322 VSS.n14321 0.00299305
R10175 VSS.n14217 VSS.n573 0.00299305
R10176 VSS.n14221 VSS.n574 0.00299305
R10177 VSS.n580 VSS.n575 0.00299305
R10178 VSS.n14169 VSS.n576 0.00299305
R10179 VSS.n14163 VSS.n571 0.00299305
R10180 VSS.n14231 VSS.n14230 0.00299305
R10181 VSS.n559 VSS.n548 0.00299305
R10182 VSS.n558 VSS.n557 0.00299305
R10183 VSS.n10703 VSS.n10702 0.00299305
R10184 VSS.n10670 VSS.n10669 0.00299305
R10185 VSS.n10664 VSS.n10663 0.00299305
R10186 VSS.n10658 VSS.n10657 0.00299305
R10187 VSS.n10692 VSS.n10689 0.00299305
R10188 VSS.n10705 VSS.n10654 0.00299305
R10189 VSS.n10687 VSS.n10683 0.00299305
R10190 VSS.n10681 VSS.n10677 0.00299305
R10191 VSS.n14271 VSS.n14270 0.00299305
R10192 VSS.n14276 VSS.n509 0.00299305
R10193 VSS.n519 VSS.n518 0.00299305
R10194 VSS.n14259 VSS.n14258 0.00299305
R10195 VSS.n535 VSS.n534 0.00299305
R10196 VSS.n529 VSS.n528 0.00299305
R10197 VSS.n523 VSS.n522 0.00299305
R10198 VSS.n14203 VSS.n14202 0.00299305
R10199 VSS.n591 VSS.n587 0.00299305
R10200 VSS.n601 VSS.n590 0.00299305
R10201 VSS.n592 VSS.n589 0.00299305
R10202 VSS.n1137 VSS.n916 0.00299305
R10203 VSS.n1145 VSS.n931 0.00299305
R10204 VSS.n933 VSS.n932 0.00299305
R10205 VSS.n1141 VSS.n930 0.00299305
R10206 VSS.n928 VSS.n913 0.00299305
R10207 VSS.n1153 VSS.n1152 0.00299305
R10208 VSS.n927 VSS.n926 0.00299305
R10209 VSS.n920 VSS.n917 0.00299305
R10210 VSS.n13115 VSS.n13109 0.00299305
R10211 VSS.n13123 VSS.n13122 0.00299305
R10212 VSS.n13124 VSS.n2348 0.00299305
R10213 VSS.n13135 VSS.n13134 0.00299305
R10214 VSS.n1915 VSS.n1914 0.00299305
R10215 VSS.n1921 VSS.n1916 0.00299305
R10216 VSS.n1927 VSS.n1926 0.00299305
R10217 VSS.n2467 VSS.n2466 0.00299305
R10218 VSS.n2477 VSS.n2464 0.00299305
R10219 VSS.n13055 VSS.n13054 0.00299305
R10220 VSS.n12416 VSS.n12415 0.00299305
R10221 VSS.n12413 VSS.n12412 0.00299305
R10222 VSS.n12406 VSS.n12400 0.00299305
R10223 VSS.n12405 VSS.n12404 0.00299305
R10224 VSS.n12450 VSS.n12449 0.00299305
R10225 VSS.n12444 VSS.n12443 0.00299305
R10226 VSS.n12438 VSS.n12437 0.00299305
R10227 VSS.n12394 VSS.n12393 0.00299305
R10228 VSS.n2496 VSS.n2487 0.00299305
R10229 VSS.n2495 VSS.n2494 0.00299305
R10230 VSS.n13037 VSS.n2493 0.00299305
R10231 VSS.n2540 VSS.n2488 0.00299305
R10232 VSS.n2536 VSS.n2490 0.00299305
R10233 VSS.n2491 VSS.n2485 0.00299305
R10234 VSS.n2544 VSS.n2489 0.00299305
R10235 VSS.n13071 VSS.n13070 0.00299305
R10236 VSS.n13087 VSS.n13086 0.00299305
R10237 VSS.n13084 VSS.n13074 0.00299305
R10238 VSS.n13080 VSS.n13079 0.00299305
R10239 VSS.n2451 VSS.n2450 0.00299305
R10240 VSS.n2442 VSS.n2441 0.00299305
R10241 VSS.n2440 VSS.n2439 0.00299305
R10242 VSS.n2435 VSS.n2432 0.00299305
R10243 VSS.n2371 VSS.n2358 0.00299305
R10244 VSS.n13102 VSS.n2355 0.00299305
R10245 VSS.n2370 VSS.n2354 0.00299305
R10246 VSS.n2379 VSS.n2359 0.00299305
R10247 VSS.n2387 VSS.n2361 0.00299305
R10248 VSS.n2373 VSS.n2362 0.00299305
R10249 VSS.n2384 VSS.n2360 0.00299305
R10250 VSS.n2328 VSS.n1935 0.00299305
R10251 VSS.n2336 VSS.n1941 0.00299305
R10252 VSS.n1943 VSS.n1942 0.00299305
R10253 VSS.n2332 VSS.n1940 0.00299305
R10254 VSS.n1939 VSS.n1933 0.00299305
R10255 VSS.n2293 VSS.n1938 0.00299305
R10256 VSS.n2289 VSS.n1937 0.00299305
R10257 VSS.n2285 VSS.n1936 0.00299305
R10258 VSS.n14167 VSS.n578 0.00299305
R10259 VSS.n2405 VSS.n551 0.00299305
R10260 VSS.n2416 VSS.n550 0.00299305
R10261 VSS.n2413 VSS.n553 0.00299305
R10262 VSS.n2410 VSS.n552 0.00299305
R10263 VSS.n1164 VSS.n885 0.00299305
R10264 VSS.n895 VSS.n894 0.00299305
R10265 VSS.n905 VSS.n893 0.00299305
R10266 VSS.n902 VSS.n892 0.00299305
R10267 VSS.n938 VSS.n890 0.00299305
R10268 VSS.n944 VSS.n889 0.00299305
R10269 VSS.n948 VSS.n888 0.00299305
R10270 VSS.n951 VSS.n887 0.00299305
R10271 VSS.n1384 VSS.n1383 0.00299305
R10272 VSS.n1387 VSS.n1386 0.00299305
R10273 VSS.n1397 VSS.n1396 0.00299305
R10274 VSS.n866 VSS.n865 0.00299305
R10275 VSS.n872 VSS.n867 0.00299305
R10276 VSS.n878 VSS.n877 0.00299305
R10277 VSS.n1376 VSS.n1375 0.00299305
R10278 VSS.n14299 VSS.n14298 0.00299305
R10279 VSS.n14293 VSS.n14292 0.00299305
R10280 VSS.n14333 VSS.n14282 0.00299305
R10281 VSS.n14287 VSS.n14286 0.00299305
R10282 VSS.n1566 VSS.n1565 0.00299305
R10283 VSS.n1559 VSS.n1558 0.00299305
R10284 VSS.n1553 VSS.n1552 0.00299305
R10285 VSS.n1547 VSS.n1546 0.00299305
R10286 VSS.n1541 VSS.n1540 0.00299305
R10287 VSS.n1535 VSS.n1534 0.00299305
R10288 VSS.n1570 VSS.n1519 0.00299305
R10289 VSS.n1529 VSS.n1528 0.00299305
R10290 VSS.n13741 VSS.n13740 0.00299305
R10291 VSS.n13850 VSS.n13849 0.00299305
R10292 VSS.n13856 VSS.n13855 0.00299305
R10293 VSS.n13725 VSS.n13724 0.00299305
R10294 VSS.n13731 VSS.n13730 0.00299305
R10295 VSS.n13735 VSS.n13734 0.00299305
R10296 VSS.n13711 VSS.n13707 0.00299305
R10297 VSS.n13806 VSS.n13805 0.00299305
R10298 VSS.n13799 VSS.n13798 0.00299305
R10299 VSS.n13793 VSS.n13792 0.00299305
R10300 VSS.n13787 VSS.n13786 0.00299305
R10301 VSS.n13781 VSS.n13780 0.00299305
R10302 VSS.n13775 VSS.n13774 0.00299305
R10303 VSS.n13810 VSS.n13759 0.00299305
R10304 VSS.n13769 VSS.n13768 0.00299305
R10305 VSS.n13278 VSS.n13277 0.00299305
R10306 VSS.n13385 VSS.n13384 0.00299305
R10307 VSS.n13391 VSS.n13390 0.00299305
R10308 VSS.n13262 VSS.n13261 0.00299305
R10309 VSS.n13268 VSS.n13267 0.00299305
R10310 VSS.n13272 VSS.n13271 0.00299305
R10311 VSS.n13248 VSS.n13244 0.00299305
R10312 VSS.n1491 VSS.n1487 0.00299305
R10313 VSS.n1497 VSS.n1493 0.00299305
R10314 VSS.n1607 VSS.n1499 0.00299305
R10315 VSS.n759 VSS.n758 0.00299305
R10316 VSS.n752 VSS.n751 0.00299305
R10317 VSS.n746 VSS.n745 0.00299305
R10318 VSS.n740 VSS.n739 0.00299305
R10319 VSS.n734 VSS.n733 0.00299305
R10320 VSS.n728 VSS.n727 0.00299305
R10321 VSS.n763 VSS.n712 0.00299305
R10322 VSS.n722 VSS.n721 0.00299305
R10323 VSS.n14113 VSS.n649 0.00299305
R10324 VSS.n14117 VSS.n14116 0.00299305
R10325 VSS.n648 VSS.n647 0.00299305
R10326 VSS.n641 VSS.n639 0.00299305
R10327 VSS.n1444 VSS.n637 0.00299305
R10328 VSS.n1446 VSS.n636 0.00299305
R10329 VSS.n1453 VSS.n635 0.00299305
R10330 VSS.n1455 VSS.n634 0.00299305
R10331 VSS.n14101 VSS.n14100 0.00299305
R10332 VSS.n14104 VSS.n14103 0.00299305
R10333 VSS.n1689 VSS.n1688 0.00299305
R10334 VSS.n1692 VSS.n1691 0.00299305
R10335 VSS.n1683 VSS.n1682 0.00299305
R10336 VSS.n1677 VSS.n1676 0.00299305
R10337 VSS.n14093 VSS.n14092 0.00299305
R10338 VSS.n13660 VSS.n13654 0.00299305
R10339 VSS.n13667 VSS.n13666 0.00299305
R10340 VSS.n13699 VSS.n13669 0.00299305
R10341 VSS.n13690 VSS.n13689 0.00299305
R10342 VSS.n13682 VSS.n13681 0.00299305
R10343 VSS.n13679 VSS.n13678 0.00299305
R10344 VSS.n1663 VSS.n1660 0.00299305
R10345 VSS.n14073 VSS.n1659 0.00299305
R10346 VSS.n14063 VSS.n1658 0.00299305
R10347 VSS.n14067 VSS.n1657 0.00299305
R10348 VSS.n1650 VSS.n1649 0.00299305
R10349 VSS.n1651 VSS.n1648 0.00299305
R10350 VSS.n14081 VSS.n14080 0.00299305
R10351 VSS.n1664 VSS.n1647 0.00299305
R10352 VSS.n13894 VSS.n13649 0.00299305
R10353 VSS.n13905 VSS.n13904 0.00299305
R10354 VSS.n13208 VSS.n13207 0.00299305
R10355 VSS.n13214 VSS.n13209 0.00299305
R10356 VSS.n13220 VSS.n13219 0.00299305
R10357 VSS.n13237 VSS.n13228 0.00299305
R10358 VSS.n13236 VSS.n13235 0.00299305
R10359 VSS.n13635 VSS.n13234 0.00299305
R10360 VSS.n13539 VSS.n13229 0.00299305
R10361 VSS.n13535 VSS.n13231 0.00299305
R10362 VSS.n13232 VSS.n13226 0.00299305
R10363 VSS.n13543 VSS.n13230 0.00299305
R10364 VSS.n13885 VSS.n13879 0.00299305
R10365 VSS.n13893 VSS.n13892 0.00299305
R10366 VSS.n824 VSS.n823 0.00299305
R10367 VSS.n834 VSS.n816 0.00299305
R10368 VSS.n1436 VSS.n817 0.00299305
R10369 VSS.n1409 VSS.n1408 0.00299305
R10370 VSS.n848 VSS.n845 0.00299305
R10371 VSS.n857 VSS.n856 0.00299305
R10372 VSS.n854 VSS.n853 0.00299305
R10373 VSS.n1182 VSS.n1181 0.00299305
R10374 VSS.n1184 VSS.n1175 0.00299305
R10375 VSS.n1189 VSS.n1188 0.00299305
R10376 VSS.n1192 VSS.n1191 0.00299305
R10377 VSS.n2224 VSS.n2218 0.00299305
R10378 VSS.n2232 VSS.n2231 0.00299305
R10379 VSS.n2234 VSS.n2233 0.00299305
R10380 VSS.n2192 VSS.n2191 0.00299305
R10381 VSS.n2198 VSS.n2197 0.00299305
R10382 VSS.n2201 VSS.n2200 0.00299305
R10383 VSS.n2243 VSS.n2004 0.00299305
R10384 VSS.n2247 VSS.n2246 0.00299305
R10385 VSS.n2003 VSS.n2002 0.00299305
R10386 VSS.n1996 VSS.n1994 0.00299305
R10387 VSS.n2038 VSS.n1992 0.00299305
R10388 VSS.n2040 VSS.n1991 0.00299305
R10389 VSS.n2047 VSS.n1990 0.00299305
R10390 VSS.n2049 VSS.n1989 0.00299305
R10391 VSS.n2159 VSS.n2153 0.00299305
R10392 VSS.n2167 VSS.n2166 0.00299305
R10393 VSS.n2169 VSS.n2168 0.00299305
R10394 VSS.n2120 VSS.n2106 0.00299305
R10395 VSS.n2111 VSS.n2110 0.00299305
R10396 VSS.n2118 VSS.n2117 0.00299305
R10397 VSS.n2178 VSS.n2079 0.00299305
R10398 VSS.n2182 VSS.n2181 0.00299305
R10399 VSS.n2078 VSS.n2077 0.00299305
R10400 VSS.n2071 VSS.n2069 0.00299305
R10401 VSS.n2087 VSS.n2067 0.00299305
R10402 VSS.n2089 VSS.n2066 0.00299305
R10403 VSS.n2096 VSS.n2065 0.00299305
R10404 VSS.n2098 VSS.n2064 0.00299305
R10405 VSS.n1837 VSS.n1836 0.00299305
R10406 VSS.n1848 VSS.n1847 0.00299305
R10407 VSS.n13197 VSS.n1834 0.00299305
R10408 VSS.n12655 VSS.n12654 0.00299305
R10409 VSS.n12661 VSS.n12660 0.00299305
R10410 VSS.n12664 VSS.n12663 0.00299305
R10411 VSS.n13187 VSS.n1856 0.00299305
R10412 VSS.n1866 VSS.n1865 0.00299305
R10413 VSS.n1876 VSS.n1864 0.00299305
R10414 VSS.n1873 VSS.n1863 0.00299305
R10415 VSS.n2135 VSS.n1861 0.00299305
R10416 VSS.n2139 VSS.n1860 0.00299305
R10417 VSS.n2146 VSS.n1859 0.00299305
R10418 VSS.n2143 VSS.n1858 0.00299305
R10419 VSS.n13922 VSS.n13921 0.00299305
R10420 VSS.n12689 VSS.n12688 0.00299305
R10421 VSS.n12685 VSS.n12684 0.00299305
R10422 VSS.n12678 VSS.n12672 0.00299305
R10423 VSS.n12677 VSS.n12676 0.00299305
R10424 VSS.n1792 VSS.n1779 0.00299305
R10425 VSS.n13936 VSS.n1776 0.00299305
R10426 VSS.n1791 VSS.n1775 0.00299305
R10427 VSS.n1800 VSS.n1780 0.00299305
R10428 VSS.n1808 VSS.n1782 0.00299305
R10429 VSS.n1794 VSS.n1783 0.00299305
R10430 VSS.n1805 VSS.n1781 0.00299305
R10431 VSS.n1826 VSS.n1825 0.00299305
R10432 VSS.n1819 VSS.n1817 0.00299305
R10433 VSS.n2026 VSS.n2025 0.00299305
R10434 VSS.n1974 VSS.n1971 0.00299305
R10435 VSS.n2313 VSS.n1970 0.00299305
R10436 VSS.n2309 VSS.n1969 0.00299305
R10437 VSS.n2304 VSS.n1968 0.00299305
R10438 VSS.n2320 VSS.n1952 0.00299305
R10439 VSS.n1966 VSS.n1951 0.00299305
R10440 VSS.n1956 VSS.n1955 0.00299305
R10441 VSS.n12983 VSS.n2583 0.00299305
R10442 VSS.n12987 VSS.n12986 0.00299305
R10443 VSS.n2582 VSS.n2581 0.00299305
R10444 VSS.n2575 VSS.n2573 0.00299305
R10445 VSS.n2645 VSS.n2571 0.00299305
R10446 VSS.n2647 VSS.n2570 0.00299305
R10447 VSS.n2654 VSS.n2569 0.00299305
R10448 VSS.n2656 VSS.n2568 0.00299305
R10449 VSS.n12964 VSS.n12958 0.00299305
R10450 VSS.n2719 VSS.n2718 0.00299305
R10451 VSS.n2715 VSS.n2714 0.00299305
R10452 VSS.n2708 VSS.n2702 0.00299305
R10453 VSS.n2707 VSS.n2706 0.00299305
R10454 VSS.n12974 VSS.n12973 0.00299305
R10455 VSS.n12972 VSS.n12971 0.00299305
R10456 VSS.n2690 VSS.n2687 0.00299305
R10457 VSS.n12943 VSS.n2686 0.00299305
R10458 VSS.n12933 VSS.n2685 0.00299305
R10459 VSS.n12937 VSS.n2684 0.00299305
R10460 VSS.n2677 VSS.n2676 0.00299305
R10461 VSS.n2678 VSS.n2675 0.00299305
R10462 VSS.n12951 VSS.n12950 0.00299305
R10463 VSS.n2691 VSS.n2674 0.00299305
R10464 VSS.n2774 VSS.n2772 0.00299305
R10465 VSS.n2809 VSS.n2808 0.00299305
R10466 VSS.n2791 VSS.n2790 0.00299305
R10467 VSS.n2799 VSS.n2798 0.00299305
R10468 VSS.n2797 VSS.n2796 0.00299305
R10469 VSS.n2817 VSS.n2816 0.00299305
R10470 VSS.n2785 VSS.n2784 0.00299305
R10471 VSS.n12906 VSS.n2764 0.00299305
R10472 VSS.n12910 VSS.n12909 0.00299305
R10473 VSS.n2763 VSS.n2762 0.00299305
R10474 VSS.n2756 VSS.n2754 0.00299305
R10475 VSS.n2826 VSS.n2752 0.00299305
R10476 VSS.n2828 VSS.n2751 0.00299305
R10477 VSS.n2835 VSS.n2750 0.00299305
R10478 VSS.n2837 VSS.n2749 0.00299305
R10479 VSS.n12887 VSS.n12881 0.00299305
R10480 VSS.n2899 VSS.n2898 0.00299305
R10481 VSS.n2895 VSS.n2894 0.00299305
R10482 VSS.n2888 VSS.n2882 0.00299305
R10483 VSS.n2887 VSS.n2886 0.00299305
R10484 VSS.n12897 VSS.n12896 0.00299305
R10485 VSS.n12895 VSS.n12894 0.00299305
R10486 VSS.n3044 VSS.n3038 0.00299305
R10487 VSS.n3051 VSS.n3050 0.00299305
R10488 VSS.n12640 VSS.n3053 0.00299305
R10489 VSS.n12631 VSS.n12630 0.00299305
R10490 VSS.n12623 VSS.n12622 0.00299305
R10491 VSS.n12620 VSS.n12619 0.00299305
R10492 VSS.n2870 VSS.n2867 0.00299305
R10493 VSS.n12866 VSS.n2866 0.00299305
R10494 VSS.n12856 VSS.n2865 0.00299305
R10495 VSS.n12860 VSS.n2864 0.00299305
R10496 VSS.n2857 VSS.n2856 0.00299305
R10497 VSS.n2858 VSS.n2855 0.00299305
R10498 VSS.n12874 VSS.n12873 0.00299305
R10499 VSS.n2871 VSS.n2854 0.00299305
R10500 VSS.n12717 VSS.n12716 0.00299305
R10501 VSS.n3080 VSS.n3079 0.00299305
R10502 VSS.n3076 VSS.n3075 0.00299305
R10503 VSS.n3069 VSS.n3063 0.00299305
R10504 VSS.n3068 VSS.n3067 0.00299305
R10505 VSS.n2970 VSS.n2957 0.00299305
R10506 VSS.n12731 VSS.n2954 0.00299305
R10507 VSS.n2969 VSS.n2953 0.00299305
R10508 VSS.n3005 VSS.n2958 0.00299305
R10509 VSS.n3013 VSS.n2960 0.00299305
R10510 VSS.n2972 VSS.n2961 0.00299305
R10511 VSS.n3010 VSS.n2959 0.00299305
R10512 VSS.n3031 VSS.n3030 0.00299305
R10513 VSS.n3024 VSS.n3022 0.00299305
R10514 VSS.n2606 VSS.n2605 0.00299305
R10515 VSS.n2526 VSS.n2523 0.00299305
R10516 VSS.n13018 VSS.n2522 0.00299305
R10517 VSS.n13014 VSS.n2521 0.00299305
R10518 VSS.n13009 VSS.n2520 0.00299305
R10519 VSS.n13025 VSS.n2504 0.00299305
R10520 VSS.n2518 VSS.n2503 0.00299305
R10521 VSS.n2508 VSS.n2507 0.00299305
R10522 VSS.n11677 VSS.n11571 0.00299305
R10523 VSS.n11673 VSS.n11672 0.00299305
R10524 VSS.n11667 VSS.n11666 0.00299305
R10525 VSS.n11661 VSS.n11660 0.00299305
R10526 VSS.n11655 VSS.n11654 0.00299305
R10527 VSS.n11649 VSS.n11648 0.00299305
R10528 VSS.n11643 VSS.n11642 0.00299305
R10529 VSS.n11581 VSS.n11580 0.00299305
R10530 VSS.n12227 VSS.n12226 0.00299305
R10531 VSS.n12259 VSS.n12258 0.00299305
R10532 VSS.n12243 VSS.n12242 0.00299305
R10533 VSS.n12237 VSS.n12236 0.00299305
R10534 VSS.n12231 VSS.n12230 0.00299305
R10535 VSS.n12215 VSS.n12210 0.00299305
R10536 VSS.n12221 VSS.n12217 0.00299305
R10537 VSS.n11746 VSS.n11695 0.00299305
R10538 VSS.n11742 VSS.n11741 0.00299305
R10539 VSS.n11736 VSS.n11735 0.00299305
R10540 VSS.n11730 VSS.n11729 0.00299305
R10541 VSS.n11724 VSS.n11723 0.00299305
R10542 VSS.n11718 VSS.n11717 0.00299305
R10543 VSS.n11712 VSS.n11711 0.00299305
R10544 VSS.n11705 VSS.n11704 0.00299305
R10545 VSS.n12120 VSS.n12119 0.00299305
R10546 VSS.n12152 VSS.n12151 0.00299305
R10547 VSS.n12136 VSS.n12135 0.00299305
R10548 VSS.n12130 VSS.n12129 0.00299305
R10549 VSS.n12124 VSS.n12123 0.00299305
R10550 VSS.n12108 VSS.n12046 0.00299305
R10551 VSS.n12114 VSS.n12110 0.00299305
R10552 VSS.n12095 VSS.n12094 0.00299305
R10553 VSS.n12088 VSS.n12087 0.00299305
R10554 VSS.n12082 VSS.n12081 0.00299305
R10555 VSS.n12076 VSS.n12075 0.00299305
R10556 VSS.n12070 VSS.n12069 0.00299305
R10557 VSS.n12064 VSS.n12063 0.00299305
R10558 VSS.n12099 VSS.n12048 0.00299305
R10559 VSS.n12058 VSS.n12057 0.00299305
R10560 VSS.n11952 VSS.n11951 0.00299305
R10561 VSS.n11984 VSS.n11983 0.00299305
R10562 VSS.n11968 VSS.n11967 0.00299305
R10563 VSS.n11962 VSS.n11961 0.00299305
R10564 VSS.n11956 VSS.n11955 0.00299305
R10565 VSS.n11940 VSS.n11935 0.00299305
R10566 VSS.n11946 VSS.n11942 0.00299305
R10567 VSS.n11878 VSS.n11827 0.00299305
R10568 VSS.n11874 VSS.n11873 0.00299305
R10569 VSS.n11868 VSS.n11867 0.00299305
R10570 VSS.n11862 VSS.n11861 0.00299305
R10571 VSS.n11856 VSS.n11855 0.00299305
R10572 VSS.n11850 VSS.n11849 0.00299305
R10573 VSS.n11844 VSS.n11843 0.00299305
R10574 VSS.n11837 VSS.n11836 0.00299305
R10575 VSS.n3524 VSS.n3523 0.00299305
R10576 VSS.n3556 VSS.n3555 0.00299305
R10577 VSS.n3540 VSS.n3539 0.00299305
R10578 VSS.n3534 VSS.n3533 0.00299305
R10579 VSS.n3528 VSS.n3527 0.00299305
R10580 VSS.n3512 VSS.n3450 0.00299305
R10581 VSS.n3518 VSS.n3514 0.00299305
R10582 VSS.n3499 VSS.n3498 0.00299305
R10583 VSS.n3492 VSS.n3491 0.00299305
R10584 VSS.n3486 VSS.n3485 0.00299305
R10585 VSS.n3480 VSS.n3479 0.00299305
R10586 VSS.n3474 VSS.n3473 0.00299305
R10587 VSS.n3468 VSS.n3467 0.00299305
R10588 VSS.n3503 VSS.n3452 0.00299305
R10589 VSS.n3462 VSS.n3461 0.00299305
R10590 VSS.n3099 VSS.n3098 0.00299305
R10591 VSS.n12592 VSS.n12591 0.00299305
R10592 VSS.n3115 VSS.n3114 0.00299305
R10593 VSS.n3109 VSS.n3108 0.00299305
R10594 VSS.n3103 VSS.n3102 0.00299305
R10595 VSS.n12606 VSS.n3087 0.00299305
R10596 VSS.n3093 VSS.n3089 0.00299305
R10597 VSS.n3163 VSS.n3162 0.00299305
R10598 VSS.n3167 VSS.n3166 0.00299305
R10599 VSS.n3126 VSS.n3125 0.00299305
R10600 VSS.n3132 VSS.n3131 0.00299305
R10601 VSS.n3136 VSS.n3135 0.00299305
R10602 VSS.n3227 VSS.n3226 0.00299305
R10603 VSS.n3258 VSS.n3257 0.00299305
R10604 VSS.n3264 VSS.n3263 0.00299305
R10605 VSS.n3268 VSS.n3217 0.00299305
R10606 VSS.n3250 VSS.n3249 0.00299305
R10607 VSS.n3243 VSS.n3242 0.00299305
R10608 VSS.n3237 VSS.n3236 0.00299305
R10609 VSS.n3231 VSS.n3230 0.00299305
R10610 VSS.n3151 VSS.n3147 0.00299305
R10611 VSS.n3157 VSS.n3153 0.00299305
R10612 VSS.n11611 VSS.n11610 0.00299305
R10613 VSS.n11632 VSS.n11631 0.00299305
R10614 VSS.n11622 VSS.n11621 0.00299305
R10615 VSS.n11617 VSS.n11613 0.00299305
R10616 VSS.n11601 VSS.n11597 0.00299305
R10617 VSS.n11595 VSS.n11591 0.00299305
R10618 VSS.n11589 VSS.n11585 0.00299305
R10619 VSS.n12371 VSS.n12370 0.00299305
R10620 VSS.n12454 VSS.n12366 0.00299305
R10621 VSS.n12381 VSS.n12380 0.00299305
R10622 VSS.n12375 VSS.n12374 0.00299305
R10623 VSS.n12745 VSS.n12744 0.00299305
R10624 VSS.n12746 VSS.n2947 0.00299305
R10625 VSS.n12755 VSS.n12754 0.00299305
R10626 VSS.n12775 VSS.n2936 0.00299305
R10627 VSS.n12773 VSS.n2937 0.00299305
R10628 VSS.n12763 VSS.n2939 0.00299305
R10629 VSS.n13950 VSS.n13944 0.00299305
R10630 VSS.n13958 VSS.n13957 0.00299305
R10631 VSS.n13959 VSS.n1769 0.00299305
R10632 VSS.n14018 VSS.n14017 0.00299305
R10633 VSS.n1725 VSS.n1721 0.00299305
R10634 VSS.n1724 VSS.n1723 0.00299305
R10635 VSS.n13567 VSS.n13566 0.00299305
R10636 VSS.n13560 VSS.n13558 0.00299305
R10637 VSS.n13578 VSS.n13577 0.00299305
R10638 VSS.n13605 VSS.n13604 0.00299305
R10639 VSS.n13490 VSS.n13486 0.00299305
R10640 VSS.n13489 VSS.n13488 0.00299305
R10641 VSS.n13334 VSS.n13330 0.00299305
R10642 VSS.n13340 VSS.n13336 0.00299305
R10643 VSS.n13345 VSS.n13296 0.00299305
R10644 VSS.n13409 VSS.n13408 0.00299305
R10645 VSS.n13436 VSS.n13435 0.00299305
R10646 VSS.n13446 VSS.n13445 0.00299305
R10647 VSS.n828 VSS.n822 0.00299304
R10648 VSS.n1485 VSS.n1484 0.00299304
R10649 VSS.n7924 VSS.n7888 0.00299304
R10650 VSS.n9175 VSS.n9169 0.00299304
R10651 VSS.n9339 VSS.n9338 0.00299304
R10652 VSS.n9682 VSS.n9680 0.00299304
R10653 VSS.n9052 VSS.n9051 0.00299304
R10654 VSS.n8351 VSS.n8350 0.00299304
R10655 VSS.n8694 VSS.n8692 0.00299304
R10656 VSS.n9624 VSS.n9623 0.00299304
R10657 VSS.n8305 VSS.n8304 0.00299304
R10658 VSS.n8249 VSS.n8248 0.00299304
R10659 VSS.n8853 VSS.n8851 0.00299304
R10660 VSS.n9958 VSS.n9957 0.00299304
R10661 VSS.n6193 VSS.n6192 0.00299304
R10662 VSS.n8449 VSS.n8448 0.00299304
R10663 VSS.n9816 VSS.n9815 0.00299304
R10664 VSS.n7355 VSS.n7272 0.00299304
R10665 VSS.n7199 VSS.n7194 0.00299304
R10666 VSS.n7834 VSS.n7815 0.00299304
R10667 VSS.n7789 VSS.n7788 0.00299304
R10668 VSS.n7710 VSS.n7709 0.00299304
R10669 VSS.n7124 VSS.n7116 0.00299304
R10670 VSS.n9873 VSS.n9872 0.00299304
R10671 VSS.n7984 VSS.n7983 0.00299304
R10672 VSS.n6888 VSS.n6887 0.00299304
R10673 VSS.n6961 VSS.n6960 0.00299304
R10674 VSS.n7004 VSS.n6517 0.00299304
R10675 VSS.n6281 VSS.n6275 0.00299304
R10676 VSS.n6409 VSS.n6326 0.00299304
R10677 VSS.n6435 VSS.n6434 0.00299304
R10678 VSS.n6821 VSS.n6820 0.00299304
R10679 VSS.n6721 VSS.n6680 0.00299304
R10680 VSS.n5894 VSS.n5892 0.00299304
R10681 VSS.n5713 VSS.n5711 0.00299304
R10682 VSS.n5533 VSS.n5531 0.00299304
R10683 VSS.n5353 VSS.n5351 0.00299304
R10684 VSS.n10087 VSS.n10085 0.00299304
R10685 VSS.n3796 VSS.n3795 0.00299304
R10686 VSS.n4611 VSS.n4609 0.00299304
R10687 VSS.n5990 VSS.n5988 0.00299304
R10688 VSS.n3741 VSS.n3739 0.00299304
R10689 VSS.n11060 VSS.n11059 0.00299304
R10690 VSS.n6337 VSS.n6336 0.00299304
R10691 VSS.n11013 VSS.n3833 0.00299304
R10692 VSS.n10973 VSS.n3873 0.00299304
R10693 VSS.n10907 VSS.n10906 0.00299304
R10694 VSS.n7283 VSS.n7282 0.00299304
R10695 VSS.n10862 VSS.n3901 0.00299304
R10696 VSS.n4001 VSS.n3999 0.00299304
R10697 VSS.n4043 VSS.n4042 0.00299304
R10698 VSS.n4388 VSS.n4190 0.00299304
R10699 VSS.n4284 VSS.n4283 0.00299304
R10700 VSS.n4243 VSS.n4236 0.00299304
R10701 VSS.n4121 VSS.n4119 0.00299304
R10702 VSS.n10755 VSS.n10754 0.00299304
R10703 VSS.n1288 VSS.n1286 0.00299304
R10704 VSS.n686 VSS.n685 0.00299304
R10705 VSS.n1216 VSS.n1215 0.00299304
R10706 VSS.n964 VSS.n963 0.00299304
R10707 VSS.n14212 VSS.n572 0.00299304
R10708 VSS.n561 VSS.n556 0.00299304
R10709 VSS.n14265 VSS.n14264 0.00299304
R10710 VSS.n13114 VSS.n13113 0.00299304
R10711 VSS.n2469 VSS.n2465 0.00299304
R10712 VSS.n13033 VSS.n2492 0.00299304
R10713 VSS.n2365 VSS.n2364 0.00299304
R10714 VSS.n13659 VSS.n13658 0.00299304
R10715 VSS.n13631 VSS.n13233 0.00299304
R10716 VSS.n13884 VSS.n13883 0.00299304
R10717 VSS.n2223 VSS.n2222 0.00299304
R10718 VSS.n2158 VSS.n2157 0.00299304
R10719 VSS.n1841 VSS.n1835 0.00299304
R10720 VSS.n1786 VSS.n1785 0.00299304
R10721 VSS.n1824 VSS.n1823 0.00299304
R10722 VSS.n2018 VSS.n2017 0.00299304
R10723 VSS.n1958 VSS.n1954 0.00299304
R10724 VSS.n12963 VSS.n12962 0.00299304
R10725 VSS.n2777 VSS.n2776 0.00299304
R10726 VSS.n12886 VSS.n12885 0.00299304
R10727 VSS.n3043 VSS.n3042 0.00299304
R10728 VSS.n2964 VSS.n2963 0.00299304
R10729 VSS.n3029 VSS.n3028 0.00299304
R10730 VSS.n2598 VSS.n2597 0.00299304
R10731 VSS.n2510 VSS.n2506 0.00299304
R10732 VSS.n12255 VSS.n12253 0.00299304
R10733 VSS.n12148 VSS.n12146 0.00299304
R10734 VSS.n11980 VSS.n11978 0.00299304
R10735 VSS.n3552 VSS.n3550 0.00299304
R10736 VSS.n12604 VSS.n12602 0.00299304
R10737 VSS.n3145 VSS.n3143 0.00299304
R10738 VSS.n11605 VSS.n11603 0.00299304
R10739 VSS.n12739 VSS.n12738 0.00299304
R10740 VSS.n12767 VSS.n2938 0.00299304
R10741 VSS.n13949 VSS.n13948 0.00299304
R10742 VSS.n1729 VSS.n1722 0.00299304
R10743 VSS.n13565 VSS.n13564 0.00299304
R10744 VSS.n13494 VSS.n13487 0.00299304
R10745 VSS.n13328 VSS.n13326 0.00299304
R10746 VSS.n13440 VSS.n13439 0.00299304
R10747 VSS.n11511 VSS.n11507 0.00298917
R10748 VSS.n11318 VSS.n11317 0.00296757
R10749 VSS.n11317 VSS.n11316 0.00296757
R10750 VSS.n4488 VSS.n4487 0.00295776
R10751 VSS.n11525 VSS.n3614 0.00290614
R10752 VSS.n4501 VSS.n4478 0.00288062
R10753 VSS.n4501 VSS.n4500 0.00288062
R10754 VSS.n303 VSS.n301 0.00288044
R10755 VSS.n4515 VSS.n4467 0.00288031
R10756 VSS.n4515 VSS.n4514 0.00288031
R10757 VSS.n14393 VSS.n382 0.00288031
R10758 VSS.n14461 VSS.n37 0.00288031
R10759 VSS.n182 VSS.n180 0.00288031
R10760 VSS.n345 VSS.n344 0.00288031
R10761 VSS.n272 VSS.n271 0.00288031
R10762 VSS.n160 VSS.n159 0.00288031
R10763 VSS.n99 VSS.n98 0.00288031
R10764 VSS.n277 VSS.n276 0.00288014
R10765 VSS.n14444 VSS.n278 0.00288014
R10766 VSS.n306 VSS.n305 0.00288014
R10767 VSS.n14444 VSS.n290 0.00288014
R10768 VSS.n14394 VSS.n351 0.00288014
R10769 VSS.n14394 VSS.n367 0.00288014
R10770 VSS.n14381 VSS.n492 0.00288014
R10771 VSS.n14381 VSS.n482 0.00288014
R10772 VSS.n14381 VSS.n486 0.00288014
R10773 VSS.n14393 VSS.n14392 0.00288014
R10774 VSS.n14394 VSS.n371 0.00288014
R10775 VSS.n14455 VSS.n166 0.00288014
R10776 VSS.n188 VSS.n187 0.00288014
R10777 VSS.n14455 VSS.n170 0.00288014
R10778 VSS.n125 VSS.n124 0.00288014
R10779 VSS.n14455 VSS.n197 0.00288014
R10780 VSS.n182 VSS.n181 0.00288014
R10781 VSS.n303 VSS.n302 0.00288014
R10782 VSS.n14444 VSS.n307 0.00288014
R10783 VSS.n14444 VSS.n309 0.00288014
R10784 VSS.n14455 VSS.n185 0.00288014
R10785 VSS.n184 VSS.n183 0.00288014
R10786 VSS.n192 VSS.n191 0.00288014
R10787 VSS.n14443 VSS.n14442 0.00288014
R10788 VSS.n370 VSS.n369 0.00288014
R10789 VSS.n14394 VSS.n363 0.00288014
R10790 VSS.n366 VSS.n365 0.00288014
R10791 VSS.n14381 VSS.n478 0.00288014
R10792 VSS.n14381 VSS.n474 0.00288014
R10793 VSS.n14381 VSS.n447 0.00288014
R10794 VSS.n357 VSS.n356 0.00288014
R10795 VSS.n354 VSS.n353 0.00288014
R10796 VSS.n14394 VSS.n359 0.00288014
R10797 VSS.n14394 VSS.n355 0.00288014
R10798 VSS.n284 VSS.n283 0.00288014
R10799 VSS.n281 VSS.n280 0.00288014
R10800 VSS.n14444 VSS.n286 0.00288014
R10801 VSS.n14444 VSS.n282 0.00288014
R10802 VSS.n195 VSS.n194 0.00288014
R10803 VSS.n14455 VSS.n189 0.00288014
R10804 VSS.n14455 VSS.n193 0.00288014
R10805 VSS.n77 VSS.n66 0.00288014
R10806 VSS.n64 VSS.n63 0.00288014
R10807 VSS.n169 VSS.n168 0.00288014
R10808 VSS.n163 VSS.n162 0.00288014
R10809 VSS.n288 VSS.n287 0.00288014
R10810 VSS.n361 VSS.n360 0.00288014
R10811 VSS.n350 VSS.n349 0.00288014
R10812 VSS.n14381 VSS.n501 0.00288014
R10813 VSS.n14394 VSS.n346 0.00288014
R10814 VSS.n14444 VSS.n273 0.00288014
R10815 VSS.n14455 VSS.n161 0.00288014
R10816 VSS.n45 VSS.n44 0.00288014
R10817 VSS.n51 VSS.n50 0.00288014
R10818 VSS.n45 VSS.n43 0.00288014
R10819 VSS.n45 VSS.n39 0.00288014
R10820 VSS.n112 VSS.n111 0.00288014
R10821 VSS.n45 VSS.n40 0.00288014
R10822 VSS.n45 VSS.n42 0.00288014
R10823 VSS.n138 VSS.n137 0.00288014
R10824 VSS.n45 VSS.n41 0.00288014
R10825 VSS.n14461 VSS.n48 0.00288014
R10826 VSS.n47 VSS.n46 0.00288014
R10827 VSS.n5067 VSS.n4764 0.00258771
R10828 VSS.n5075 VSS.n4757 0.00258771
R10829 VSS.n5084 VSS.n4749 0.00258771
R10830 VSS.n5091 VSS.n4747 0.00258771
R10831 VSS.n10493 VSS.n10254 0.00258771
R10832 VSS.n10338 VSS.n10320 0.00258771
R10833 VSS.n10305 VSS.n10304 0.00258771
R10834 VSS.n5197 VSS.n5196 0.00258351
R10835 VSS.n12348 VSS.n12347 0.00257469
R10836 VSS.n11341 VSS.n11340 0.00253147
R10837 VSS.n11328 VSS.n11327 0.00253147
R10838 VSS.n11328 VSS.n11197 0.00250667
R10839 VSS.n11340 VSS.n11339 0.00250667
R10840 VSS.n13459 VSS.n13458 0.00249311
R10841 VSS.n13471 VSS.n13470 0.00249311
R10842 VSS.n13404 VSS.n13403 0.00249311
R10843 VSS.n13465 VSS.n13464 0.00249311
R10844 VSS.n13595 VSS.n13594 0.00249311
R10845 VSS.n13601 VSS.n13600 0.00249311
R10846 VSS.n13588 VSS.n13587 0.00249311
R10847 VSS.n13509 VSS.n13508 0.00249311
R10848 VSS.n14008 VSS.n14007 0.00249311
R10849 VSS.n14014 VSS.n14013 0.00249311
R10850 VSS.n1762 VSS.n1761 0.00249311
R10851 VSS.n1744 VSS.n1743 0.00249311
R10852 VSS.n12789 VSS.n12788 0.00249311
R10853 VSS.n12799 VSS.n12798 0.00249311
R10854 VSS.n12784 VSS.n2931 0.00249311
R10855 VSS.n12794 VSS.n12793 0.00249311
R10856 VSS.n4069 VSS.n4068 0.00249311
R10857 VSS.n4081 VSS.n4080 0.00249311
R10858 VSS.n4063 VSS.n4062 0.00249311
R10859 VSS.n4075 VSS.n4074 0.00249311
R10860 VSS.n10884 VSS.n10883 0.00249311
R10861 VSS.n10894 VSS.n10893 0.00249311
R10862 VSS.n10879 VSS.n3894 0.00249311
R10863 VSS.n10889 VSS.n10888 0.00249311
R10864 VSS.n10927 VSS.n10926 0.00249311
R10865 VSS.n10939 VSS.n10938 0.00249311
R10866 VSS.n10920 VSS.n10918 0.00249311
R10867 VSS.n10935 VSS.n10925 0.00249311
R10868 VSS.n11035 VSS.n11034 0.00249311
R10869 VSS.n11045 VSS.n11044 0.00249311
R10870 VSS.n11030 VSS.n3826 0.00249311
R10871 VSS.n11040 VSS.n11039 0.00249311
R10872 VSS.n9680 VSS.n9679 0.00249311
R10873 VSS.n9674 VSS.n9673 0.00249311
R10874 VSS.n9668 VSS.n9667 0.00249311
R10875 VSS.n9642 VSS.n9641 0.00249311
R10876 VSS.n9051 VSS.n9050 0.00249311
R10877 VSS.n9132 VSS.n9131 0.00249311
R10878 VSS.n9126 VSS.n9125 0.00249311
R10879 VSS.n9029 VSS.n9028 0.00249311
R10880 VSS.n9020 VSS.n9019 0.00249311
R10881 VSS.n9045 VSS.n9044 0.00249311
R10882 VSS.n9039 VSS.n9038 0.00249311
R10883 VSS.n9033 VSS.n9032 0.00249311
R10884 VSS.n9688 VSS.n9687 0.00249311
R10885 VSS.n9657 VSS.n9656 0.00249311
R10886 VSS.n9651 VSS.n9650 0.00249311
R10887 VSS.n9645 VSS.n9644 0.00249311
R10888 VSS.n8350 VSS.n8349 0.00249311
R10889 VSS.n8353 VSS.n8352 0.00249311
R10890 VSS.n8359 VSS.n8358 0.00249311
R10891 VSS.n8344 VSS.n8343 0.00249311
R10892 VSS.n8467 VSS.n8466 0.00249311
R10893 VSS.n8413 VSS.n8412 0.00249311
R10894 VSS.n8477 VSS.n8476 0.00249311
R10895 VSS.n8471 VSS.n8470 0.00249311
R10896 VSS.n8505 VSS.n8504 0.00249311
R10897 VSS.n8503 VSS.n8502 0.00249311
R10898 VSS.n8499 VSS.n8498 0.00249311
R10899 VSS.n8493 VSS.n8492 0.00249311
R10900 VSS.n8385 VSS.n8367 0.00249311
R10901 VSS.n8378 VSS.n8377 0.00249311
R10902 VSS.n8374 VSS.n8373 0.00249311
R10903 VSS.n8381 VSS.n8366 0.00249311
R10904 VSS.n8404 VSS.n8403 0.00249311
R10905 VSS.n8402 VSS.n8401 0.00249311
R10906 VSS.n8398 VSS.n8397 0.00249311
R10907 VSS.n8392 VSS.n8391 0.00249311
R10908 VSS.n8692 VSS.n8691 0.00249311
R10909 VSS.n8686 VSS.n8685 0.00249311
R10910 VSS.n8680 VSS.n8679 0.00249311
R10911 VSS.n8654 VSS.n8653 0.00249311
R10912 VSS.n9623 VSS.n9622 0.00249311
R10913 VSS.n9629 VSS.n9628 0.00249311
R10914 VSS.n7521 VSS.n7520 0.00249311
R10915 VSS.n7530 VSS.n7529 0.00249311
R10916 VSS.n9617 VSS.n9616 0.00249311
R10917 VSS.n7546 VSS.n7545 0.00249311
R10918 VSS.n7540 VSS.n7539 0.00249311
R10919 VSS.n7534 VSS.n7533 0.00249311
R10920 VSS.n8700 VSS.n8699 0.00249311
R10921 VSS.n8669 VSS.n8668 0.00249311
R10922 VSS.n8663 VSS.n8662 0.00249311
R10923 VSS.n8657 VSS.n8656 0.00249311
R10924 VSS.n8304 VSS.n8303 0.00249311
R10925 VSS.n8307 VSS.n8306 0.00249311
R10926 VSS.n8313 VSS.n8312 0.00249311
R10927 VSS.n8319 VSS.n8318 0.00249311
R10928 VSS.n8611 VSS.n8610 0.00249311
R10929 VSS.n8604 VSS.n8603 0.00249311
R10930 VSS.n8598 VSS.n8597 0.00249311
R10931 VSS.n8592 VSS.n8591 0.00249311
R10932 VSS.n8586 VSS.n8585 0.00249311
R10933 VSS.n8580 VSS.n8579 0.00249311
R10934 VSS.n8565 VSS.n8564 0.00249311
R10935 VSS.n8574 VSS.n8573 0.00249311
R10936 VSS.n8749 VSS.n8748 0.00249311
R10937 VSS.n8300 VSS.n8299 0.00249311
R10938 VSS.n8294 VSS.n8293 0.00249311
R10939 VSS.n8288 VSS.n8287 0.00249311
R10940 VSS.n8251 VSS.n8248 0.00249311
R10941 VSS.n8254 VSS.n8247 0.00249311
R10942 VSS.n8257 VSS.n8245 0.00249311
R10943 VSS.n8775 VSS.n8774 0.00249311
R10944 VSS.n8241 VSS.n8220 0.00249311
R10945 VSS.n8236 VSS.n8221 0.00249311
R10946 VSS.n8233 VSS.n8222 0.00249311
R10947 VSS.n8226 VSS.n8225 0.00249311
R10948 VSS.n8786 VSS.n8195 0.00249311
R10949 VSS.n8791 VSS.n8790 0.00249311
R10950 VSS.n8207 VSS.n8206 0.00249311
R10951 VSS.n8202 VSS.n8201 0.00249311
R10952 VSS.n6188 VSS.n6187 0.00249311
R10953 VSS.n4662 VSS.n4661 0.00249311
R10954 VSS.n6198 VSS.n6197 0.00249311
R10955 VSS.n6192 VSS.n6191 0.00249311
R10956 VSS.n9978 VSS.n6214 0.00249311
R10957 VSS.n6216 VSS.n6215 0.00249311
R10958 VSS.n6224 VSS.n6223 0.00249311
R10959 VSS.n6228 VSS.n6227 0.00249311
R10960 VSS.n6747 VSS.n6718 0.00249311
R10961 VSS.n6755 VSS.n6754 0.00249311
R10962 VSS.n6716 VSS.n6715 0.00249311
R10963 VSS.n6751 VSS.n6750 0.00249311
R10964 VSS.n6710 VSS.n6693 0.00249311
R10965 VSS.n6763 VSS.n6694 0.00249311
R10966 VSS.n6708 VSS.n6707 0.00249311
R10967 VSS.n6703 VSS.n6702 0.00249311
R10968 VSS.n6233 VSS.n6232 0.00249311
R10969 VSS.n9967 VSS.n9952 0.00249311
R10970 VSS.n9954 VSS.n9953 0.00249311
R10971 VSS.n9958 VSS.n9956 0.00249311
R10972 VSS.n8153 VSS.n8018 0.00249311
R10973 VSS.n8023 VSS.n8017 0.00249311
R10974 VSS.n8030 VSS.n8022 0.00249311
R10975 VSS.n8025 VSS.n8024 0.00249311
R10976 VSS.n8100 VSS.n8098 0.00249311
R10977 VSS.n8108 VSS.n8107 0.00249311
R10978 VSS.n8096 VSS.n8095 0.00249311
R10979 VSS.n8104 VSS.n8103 0.00249311
R10980 VSS.n8047 VSS.n8040 0.00249311
R10981 VSS.n8048 VSS.n8046 0.00249311
R10982 VSS.n8083 VSS.n8082 0.00249311
R10983 VSS.n8079 VSS.n8078 0.00249311
R10984 VSS.n8126 VSS.n8119 0.00249311
R10985 VSS.n8144 VSS.n8143 0.00249311
R10986 VSS.n8140 VSS.n8139 0.00249311
R10987 VSS.n8136 VSS.n8131 0.00249311
R10988 VSS.n8069 VSS.n8051 0.00249311
R10989 VSS.n8066 VSS.n8052 0.00249311
R10990 VSS.n8062 VSS.n8053 0.00249311
R10991 VSS.n8058 VSS.n8054 0.00249311
R10992 VSS.n8879 VSS.n7975 0.00249311
R10993 VSS.n8887 VSS.n8886 0.00249311
R10994 VSS.n7973 VSS.n7972 0.00249311
R10995 VSS.n8883 VSS.n8882 0.00249311
R10996 VSS.n7967 VSS.n7949 0.00249311
R10997 VSS.n8895 VSS.n7950 0.00249311
R10998 VSS.n7965 VSS.n7964 0.00249311
R10999 VSS.n7960 VSS.n7959 0.00249311
R11000 VSS.n8867 VSS.n8003 0.00249311
R11001 VSS.n8863 VSS.n8005 0.00249311
R11002 VSS.n8859 VSS.n8006 0.00249311
R11003 VSS.n8852 VSS.n8851 0.00249311
R11004 VSS.n8815 VSS.n8190 0.00249311
R11005 VSS.n8192 VSS.n8191 0.00249311
R11006 VSS.n8806 VSS.n8797 0.00249311
R11007 VSS.n8802 VSS.n8799 0.00249311
R11008 VSS.n8824 VSS.n8163 0.00249311
R11009 VSS.n8829 VSS.n8828 0.00249311
R11010 VSS.n8175 VSS.n8174 0.00249311
R11011 VSS.n8170 VSS.n8169 0.00249311
R11012 VSS.n9553 VSS.n7571 0.00249311
R11013 VSS.n7573 VSS.n7572 0.00249311
R11014 VSS.n7585 VSS.n7584 0.00249311
R11015 VSS.n7581 VSS.n7578 0.00249311
R11016 VSS.n8270 VSS.n8269 0.00249311
R11017 VSS.n8274 VSS.n8273 0.00249311
R11018 VSS.n8277 VSS.n8262 0.00249311
R11019 VSS.n8281 VSS.n8263 0.00249311
R11020 VSS.n9560 VSS.n7566 0.00249311
R11021 VSS.n9567 VSS.n9566 0.00249311
R11022 VSS.n9568 VSS.n7564 0.00249311
R11023 VSS.n9575 VSS.n9574 0.00249311
R11024 VSS.n9582 VSS.n9580 0.00249311
R11025 VSS.n9588 VSS.n9587 0.00249311
R11026 VSS.n9591 VSS.n7552 0.00249311
R11027 VSS.n7554 VSS.n7553 0.00249311
R11028 VSS.n9577 VSS.n7554 0.00249311
R11029 VSS.n8534 VSS.n8533 0.00249311
R11030 VSS.n8540 VSS.n8539 0.00249311
R11031 VSS.n8546 VSS.n8545 0.00249311
R11032 VSS.n8550 VSS.n8549 0.00249311
R11033 VSS.n8444 VSS.n8443 0.00249311
R11034 VSS.n8439 VSS.n8438 0.00249311
R11035 VSS.n8454 VSS.n8453 0.00249311
R11036 VSS.n8448 VSS.n8447 0.00249311
R11037 VSS.n9411 VSS.n9410 0.00249311
R11038 VSS.n9404 VSS.n9403 0.00249311
R11039 VSS.n9398 VSS.n9397 0.00249311
R11040 VSS.n9392 VSS.n9391 0.00249311
R11041 VSS.n9386 VSS.n9385 0.00249311
R11042 VSS.n9380 VSS.n9379 0.00249311
R11043 VSS.n9365 VSS.n9364 0.00249311
R11044 VSS.n9374 VSS.n9373 0.00249311
R11045 VSS.n9787 VSS.n9786 0.00249311
R11046 VSS.n7401 VSS.n7400 0.00249311
R11047 VSS.n7407 VSS.n7406 0.00249311
R11048 VSS.n7411 VSS.n7410 0.00249311
R11049 VSS.n7384 VSS.n7383 0.00249311
R11050 VSS.n7417 VSS.n7416 0.00249311
R11051 VSS.n9781 VSS.n9780 0.00249311
R11052 VSS.n7382 VSS.n7381 0.00249311
R11053 VSS.n9785 VSS.n7382 0.00249311
R11054 VSS.n7468 VSS.n7467 0.00249311
R11055 VSS.n7461 VSS.n7460 0.00249311
R11056 VSS.n7455 VSS.n7454 0.00249311
R11057 VSS.n7449 VSS.n7448 0.00249311
R11058 VSS.n7443 VSS.n7442 0.00249311
R11059 VSS.n7437 VSS.n7436 0.00249311
R11060 VSS.n7422 VSS.n7421 0.00249311
R11061 VSS.n7431 VSS.n7430 0.00249311
R11062 VSS.n10834 VSS.n10833 0.00249311
R11063 VSS.n3937 VSS.n3936 0.00249311
R11064 VSS.n3943 VSS.n3942 0.00249311
R11065 VSS.n3947 VSS.n3946 0.00249311
R11066 VSS.n3920 VSS.n3919 0.00249311
R11067 VSS.n3953 VSS.n3952 0.00249311
R11068 VSS.n10828 VSS.n10827 0.00249311
R11069 VSS.n3918 VSS.n3917 0.00249311
R11070 VSS.n10832 VSS.n3918 0.00249311
R11071 VSS.n9338 VSS.n9337 0.00249311
R11072 VSS.n9341 VSS.n9340 0.00249311
R11073 VSS.n9347 VSS.n9346 0.00249311
R11074 VSS.n9353 VSS.n9352 0.00249311
R11075 VSS.n9105 VSS.n9104 0.00249311
R11076 VSS.n9098 VSS.n9097 0.00249311
R11077 VSS.n9092 VSS.n9091 0.00249311
R11078 VSS.n9086 VSS.n9085 0.00249311
R11079 VSS.n9080 VSS.n9079 0.00249311
R11080 VSS.n9074 VSS.n9073 0.00249311
R11081 VSS.n9059 VSS.n9058 0.00249311
R11082 VSS.n9068 VSS.n9067 0.00249311
R11083 VSS.n9446 VSS.n9445 0.00249311
R11084 VSS.n9334 VSS.n9333 0.00249311
R11085 VSS.n9328 VSS.n9327 0.00249311
R11086 VSS.n9322 VSS.n9321 0.00249311
R11087 VSS.n9514 VSS.n8995 0.00249311
R11088 VSS.n9519 VSS.n9518 0.00249311
R11089 VSS.n9013 VSS.n9012 0.00249311
R11090 VSS.n9008 VSS.n9007 0.00249311
R11091 VSS.n9275 VSS.n9274 0.00249311
R11092 VSS.n9276 VSS.n9272 0.00249311
R11093 VSS.n9284 VSS.n9283 0.00249311
R11094 VSS.n9285 VSS.n9018 0.00249311
R11095 VSS.n9313 VSS.n9312 0.00249311
R11096 VSS.n9309 VSS.n9293 0.00249311
R11097 VSS.n9296 VSS.n9295 0.00249311
R11098 VSS.n9300 VSS.n9298 0.00249311
R11099 VSS.n9494 VSS.n9492 0.00249311
R11100 VSS.n9501 VSS.n9500 0.00249311
R11101 VSS.n9504 VSS.n9488 0.00249311
R11102 VSS.n9489 VSS.n9317 0.00249311
R11103 VSS.n9489 VSS.n9016 0.00249311
R11104 VSS.n7232 VSS.n7231 0.00249311
R11105 VSS.n7227 VSS.n7218 0.00249311
R11106 VSS.n7223 VSS.n7222 0.00249311
R11107 VSS.n7222 VSS.n7180 0.00249311
R11108 VSS.n7235 VSS.n7219 0.00249311
R11109 VSS.n9836 VSS.n7159 0.00249311
R11110 VSS.n9841 VSS.n9840 0.00249311
R11111 VSS.n7177 VSS.n7176 0.00249311
R11112 VSS.n7172 VSS.n7171 0.00249311
R11113 VSS.n9472 VSS.n9471 0.00249311
R11114 VSS.n9476 VSS.n9475 0.00249311
R11115 VSS.n9483 VSS.n9482 0.00249311
R11116 VSS.n9480 VSS.n9479 0.00249311
R11117 VSS.n9826 VSS.n7186 0.00249311
R11118 VSS.n9825 VSS.n9810 0.00249311
R11119 VSS.n9812 VSS.n9811 0.00249311
R11120 VSS.n9816 VSS.n9814 0.00249311
R11121 VSS.n7258 VSS.n7210 0.00249311
R11122 VSS.n7254 VSS.n7212 0.00249311
R11123 VSS.n7247 VSS.n7215 0.00249311
R11124 VSS.n7246 VSS.n7244 0.00249311
R11125 VSS.n7278 VSS.n7276 0.00249311
R11126 VSS.n7277 VSS.n7275 0.00249311
R11127 VSS.n7359 VSS.n7358 0.00249311
R11128 VSS.n7355 VSS.n7354 0.00249311
R11129 VSS.n7322 VSS.n7321 0.00249311
R11130 VSS.n7318 VSS.n7317 0.00249311
R11131 VSS.n7314 VSS.n7265 0.00249311
R11132 VSS.n7325 VSS.n7324 0.00249311
R11133 VSS.n7199 VSS.n7198 0.00249311
R11134 VSS.n7204 VSS.n7197 0.00249311
R11135 VSS.n7196 VSS.n7191 0.00249311
R11136 VSS.n7377 VSS.n7376 0.00249311
R11137 VSS.n9175 VSS.n9172 0.00249311
R11138 VSS.n9178 VSS.n9171 0.00249311
R11139 VSS.n9163 VSS.n9161 0.00249311
R11140 VSS.n9164 VSS.n9162 0.00249311
R11141 VSS.n9239 VSS.n9215 0.00249311
R11142 VSS.n9217 VSS.n9216 0.00249311
R11143 VSS.n9229 VSS.n9228 0.00249311
R11144 VSS.n9225 VSS.n9222 0.00249311
R11145 VSS.n9194 VSS.n9192 0.00249311
R11146 VSS.n9201 VSS.n9200 0.00249311
R11147 VSS.n9206 VSS.n9205 0.00249311
R11148 VSS.n9210 VSS.n9209 0.00249311
R11149 VSS.n9263 VSS.n9262 0.00249311
R11150 VSS.n9259 VSS.n9258 0.00249311
R11151 VSS.n9255 VSS.n9247 0.00249311
R11152 VSS.n9250 VSS.n9249 0.00249311
R11153 VSS.n7824 VSS.n7823 0.00249311
R11154 VSS.n7812 VSS.n7810 0.00249311
R11155 VSS.n7847 VSS.n7827 0.00249311
R11156 VSS.n8958 VSS.n7827 0.00249311
R11157 VSS.n7813 VSS.n7811 0.00249311
R11158 VSS.n8946 VSS.n7854 0.00249311
R11159 VSS.n7856 VSS.n7855 0.00249311
R11160 VSS.n7868 VSS.n7867 0.00249311
R11161 VSS.n7864 VSS.n7861 0.00249311
R11162 VSS.n7901 VSS.n7900 0.00249311
R11163 VSS.n7904 VSS.n7896 0.00249311
R11164 VSS.n7915 VSS.n7914 0.00249311
R11165 VSS.n7911 VSS.n7908 0.00249311
R11166 VSS.n8956 VSS.n8955 0.00249311
R11167 VSS.n7843 VSS.n7842 0.00249311
R11168 VSS.n7839 VSS.n7831 0.00249311
R11169 VSS.n7834 VSS.n7833 0.00249311
R11170 VSS.n7745 VSS.n7744 0.00249311
R11171 VSS.n7740 VSS.n7731 0.00249311
R11172 VSS.n7736 VSS.n7735 0.00249311
R11173 VSS.n7735 VSS.n7631 0.00249311
R11174 VSS.n7748 VSS.n7732 0.00249311
R11175 VSS.n7807 VSS.n7633 0.00249311
R11176 VSS.n8980 VSS.n8979 0.00249311
R11177 VSS.n8970 VSS.n8969 0.00249311
R11178 VSS.n8974 VSS.n8973 0.00249311
R11179 VSS.n7624 VSS.n7620 0.00249311
R11180 VSS.n7621 VSS.n7612 0.00249311
R11181 VSS.n8988 VSS.n8987 0.00249311
R11182 VSS.n7635 VSS.n7634 0.00249311
R11183 VSS.n7799 VSS.n7642 0.00249311
R11184 VSS.n7798 VSS.n7783 0.00249311
R11185 VSS.n7785 VSS.n7784 0.00249311
R11186 VSS.n7789 VSS.n7787 0.00249311
R11187 VSS.n7683 VSS.n7680 0.00249311
R11188 VSS.n7693 VSS.n7692 0.00249311
R11189 VSS.n7697 VSS.n7696 0.00249311
R11190 VSS.n7697 VSS.n7666 0.00249311
R11191 VSS.n7689 VSS.n7688 0.00249311
R11192 VSS.n7728 VSS.n7668 0.00249311
R11193 VSS.n7770 VSS.n7769 0.00249311
R11194 VSS.n7760 VSS.n7759 0.00249311
R11195 VSS.n7764 VSS.n7763 0.00249311
R11196 VSS.n7659 VSS.n7655 0.00249311
R11197 VSS.n7656 VSS.n7647 0.00249311
R11198 VSS.n7778 VSS.n7777 0.00249311
R11199 VSS.n7670 VSS.n7669 0.00249311
R11200 VSS.n7720 VSS.n7701 0.00249311
R11201 VSS.n7719 VSS.n7704 0.00249311
R11202 VSS.n7706 VSS.n7705 0.00249311
R11203 VSS.n7710 VSS.n7708 0.00249311
R11204 VSS.n9893 VSS.n7071 0.00249311
R11205 VSS.n7073 VSS.n7072 0.00249311
R11206 VSS.n7081 VSS.n7080 0.00249311
R11207 VSS.n7085 VSS.n7084 0.00249311
R11208 VSS.n7133 VSS.n7120 0.00249311
R11209 VSS.n7132 VSS.n7119 0.00249311
R11210 VSS.n7129 VSS.n7121 0.00249311
R11211 VSS.n7124 VSS.n7123 0.00249311
R11212 VSS.n7104 VSS.n7103 0.00249311
R11213 VSS.n7111 VSS.n7098 0.00249311
R11214 VSS.n7099 VSS.n7092 0.00249311
R11215 VSS.n7108 VSS.n7100 0.00249311
R11216 VSS.n9873 VSS.n9871 0.00249311
R11217 VSS.n9869 VSS.n9868 0.00249311
R11218 VSS.n9882 VSS.n9867 0.00249311
R11219 VSS.n7144 VSS.n7143 0.00249311
R11220 VSS.n7924 VSS.n7923 0.00249311
R11221 VSS.n7929 VSS.n7921 0.00249311
R11222 VSS.n7933 VSS.n7932 0.00249311
R11223 VSS.n7937 VSS.n7893 0.00249311
R11224 VSS.n8921 VSS.n7944 0.00249311
R11225 VSS.n7946 VSS.n7945 0.00249311
R11226 VSS.n8912 VSS.n8903 0.00249311
R11227 VSS.n8908 VSS.n8905 0.00249311
R11228 VSS.n7994 VSS.n7978 0.00249311
R11229 VSS.n7992 VSS.n7977 0.00249311
R11230 VSS.n7988 VSS.n7979 0.00249311
R11231 VSS.n7983 VSS.n7980 0.00249311
R11232 VSS.n8930 VSS.n7873 0.00249311
R11233 VSS.n8935 VSS.n8934 0.00249311
R11234 VSS.n7886 VSS.n7885 0.00249311
R11235 VSS.n7881 VSS.n7880 0.00249311
R11236 VSS.n6643 VSS.n6632 0.00249311
R11237 VSS.n6644 VSS.n6642 0.00249311
R11238 VSS.n6653 VSS.n6652 0.00249311
R11239 VSS.n6650 VSS.n6649 0.00249311
R11240 VSS.n6798 VSS.n6797 0.00249311
R11241 VSS.n6802 VSS.n6801 0.00249311
R11242 VSS.n6809 VSS.n6808 0.00249311
R11243 VSS.n6806 VSS.n6805 0.00249311
R11244 VSS.n6908 VSS.n6610 0.00249311
R11245 VSS.n6612 VSS.n6611 0.00249311
R11246 VSS.n6622 VSS.n6615 0.00249311
R11247 VSS.n6619 VSS.n6616 0.00249311
R11248 VSS.n6898 VSS.n6859 0.00249311
R11249 VSS.n6884 VSS.n6883 0.00249311
R11250 VSS.n6888 VSS.n6886 0.00249311
R11251 VSS.n6897 VSS.n6882 0.00249311
R11252 VSS.n6595 VSS.n6584 0.00249311
R11253 VSS.n6596 VSS.n6594 0.00249311
R11254 VSS.n6605 VSS.n6604 0.00249311
R11255 VSS.n6602 VSS.n6601 0.00249311
R11256 VSS.n6866 VSS.n6865 0.00249311
R11257 VSS.n6870 VSS.n6869 0.00249311
R11258 VSS.n6877 VSS.n6876 0.00249311
R11259 VSS.n6874 VSS.n6873 0.00249311
R11260 VSS.n6981 VSS.n6562 0.00249311
R11261 VSS.n6564 VSS.n6563 0.00249311
R11262 VSS.n6574 VSS.n6567 0.00249311
R11263 VSS.n6571 VSS.n6568 0.00249311
R11264 VSS.n6971 VSS.n6926 0.00249311
R11265 VSS.n6957 VSS.n6956 0.00249311
R11266 VSS.n6961 VSS.n6959 0.00249311
R11267 VSS.n6970 VSS.n6955 0.00249311
R11268 VSS.n6526 VSS.n6525 0.00249311
R11269 VSS.n6514 VSS.n6512 0.00249311
R11270 VSS.n6536 VSS.n6529 0.00249311
R11271 VSS.n7040 VSS.n6529 0.00249311
R11272 VSS.n6515 VSS.n6513 0.00249311
R11273 VSS.n6994 VSS.n6543 0.00249311
R11274 VSS.n6545 VSS.n6544 0.00249311
R11275 VSS.n6557 VSS.n6556 0.00249311
R11276 VSS.n6553 VSS.n6550 0.00249311
R11277 VSS.n6936 VSS.n6935 0.00249311
R11278 VSS.n6939 VSS.n6931 0.00249311
R11279 VSS.n6950 VSS.n6949 0.00249311
R11280 VSS.n6946 VSS.n6943 0.00249311
R11281 VSS.n7038 VSS.n7037 0.00249311
R11282 VSS.n7009 VSS.n7008 0.00249311
R11283 VSS.n7010 VSS.n7007 0.00249311
R11284 VSS.n7004 VSS.n7003 0.00249311
R11285 VSS.n6468 VSS.n6464 0.00249311
R11286 VSS.n6476 VSS.n6475 0.00249311
R11287 VSS.n6479 VSS.n6291 0.00249311
R11288 VSS.n6479 VSS.n6289 0.00249311
R11289 VSS.n6466 VSS.n6295 0.00249311
R11290 VSS.n6497 VSS.n6486 0.00249311
R11291 VSS.n6498 VSS.n6496 0.00249311
R11292 VSS.n6507 VSS.n6506 0.00249311
R11293 VSS.n6504 VSS.n6503 0.00249311
R11294 VSS.n7019 VSS.n7018 0.00249311
R11295 VSS.n7023 VSS.n7022 0.00249311
R11296 VSS.n7030 VSS.n7029 0.00249311
R11297 VSS.n7027 VSS.n7026 0.00249311
R11298 VSS.n7063 VSS.n7062 0.00249311
R11299 VSS.n6287 VSS.n6272 0.00249311
R11300 VSS.n6284 VSS.n6277 0.00249311
R11301 VSS.n6281 VSS.n6278 0.00249311
R11302 VSS.n6455 VSS.n6298 0.00249311
R11303 VSS.n6300 VSS.n6299 0.00249311
R11304 VSS.n6308 VSS.n6307 0.00249311
R11305 VSS.n6312 VSS.n6311 0.00249311
R11306 VSS.n6332 VSS.n6330 0.00249311
R11307 VSS.n6331 VSS.n6329 0.00249311
R11308 VSS.n6413 VSS.n6412 0.00249311
R11309 VSS.n6409 VSS.n6408 0.00249311
R11310 VSS.n6376 VSS.n6375 0.00249311
R11311 VSS.n6372 VSS.n6371 0.00249311
R11312 VSS.n6368 VSS.n6319 0.00249311
R11313 VSS.n6379 VSS.n6378 0.00249311
R11314 VSS.n6435 VSS.n6433 0.00249311
R11315 VSS.n6431 VSS.n6430 0.00249311
R11316 VSS.n6444 VSS.n6429 0.00249311
R11317 VSS.n6428 VSS.n6427 0.00249311
R11318 VSS.n6793 VSS.n6792 0.00249311
R11319 VSS.n6817 VSS.n6816 0.00249311
R11320 VSS.n6821 VSS.n6819 0.00249311
R11321 VSS.n6830 VSS.n6815 0.00249311
R11322 VSS.n6689 VSS.n6679 0.00249311
R11323 VSS.n6690 VSS.n6688 0.00249311
R11324 VSS.n6777 VSS.n6776 0.00249311
R11325 VSS.n6773 VSS.n6772 0.00249311
R11326 VSS.n6732 VSS.n6731 0.00249311
R11327 VSS.n6733 VSS.n6730 0.00249311
R11328 VSS.n6727 VSS.n6726 0.00249311
R11329 VSS.n6721 VSS.n6720 0.00249311
R11330 VSS.n6841 VSS.n6658 0.00249311
R11331 VSS.n6660 VSS.n6659 0.00249311
R11332 VSS.n6670 VSS.n6663 0.00249311
R11333 VSS.n6667 VSS.n6664 0.00249311
R11334 VSS.n6038 VSS.n6037 0.00249311
R11335 VSS.n6031 VSS.n6030 0.00249311
R11336 VSS.n6025 VSS.n6024 0.00249311
R11337 VSS.n6019 VSS.n6018 0.00249311
R11338 VSS.n6013 VSS.n6012 0.00249311
R11339 VSS.n6007 VSS.n6006 0.00249311
R11340 VSS.n5992 VSS.n5991 0.00249311
R11341 VSS.n6001 VSS.n6000 0.00249311
R11342 VSS.n5897 VSS.n5896 0.00249311
R11343 VSS.n5881 VSS.n5880 0.00249311
R11344 VSS.n5875 VSS.n5874 0.00249311
R11345 VSS.n5869 VSS.n5868 0.00249311
R11346 VSS.n5791 VSS.n5790 0.00249311
R11347 VSS.n5865 VSS.n5864 0.00249311
R11348 VSS.n5892 VSS.n5891 0.00249311
R11349 VSS.n5856 VSS.n5855 0.00249311
R11350 VSS.n5840 VSS.n5839 0.00249311
R11351 VSS.n5833 VSS.n5832 0.00249311
R11352 VSS.n5827 VSS.n5826 0.00249311
R11353 VSS.n5821 VSS.n5820 0.00249311
R11354 VSS.n5815 VSS.n5814 0.00249311
R11355 VSS.n5809 VSS.n5808 0.00249311
R11356 VSS.n5794 VSS.n5793 0.00249311
R11357 VSS.n5803 VSS.n5802 0.00249311
R11358 VSS.n5716 VSS.n5715 0.00249311
R11359 VSS.n5700 VSS.n5699 0.00249311
R11360 VSS.n5694 VSS.n5693 0.00249311
R11361 VSS.n5688 VSS.n5687 0.00249311
R11362 VSS.n5610 VSS.n5609 0.00249311
R11363 VSS.n5684 VSS.n5683 0.00249311
R11364 VSS.n5711 VSS.n5710 0.00249311
R11365 VSS.n5675 VSS.n5674 0.00249311
R11366 VSS.n5659 VSS.n5658 0.00249311
R11367 VSS.n5652 VSS.n5651 0.00249311
R11368 VSS.n5646 VSS.n5645 0.00249311
R11369 VSS.n5640 VSS.n5639 0.00249311
R11370 VSS.n5634 VSS.n5633 0.00249311
R11371 VSS.n5628 VSS.n5627 0.00249311
R11372 VSS.n5613 VSS.n5612 0.00249311
R11373 VSS.n5622 VSS.n5621 0.00249311
R11374 VSS.n5536 VSS.n5535 0.00249311
R11375 VSS.n5520 VSS.n5519 0.00249311
R11376 VSS.n5514 VSS.n5513 0.00249311
R11377 VSS.n5508 VSS.n5507 0.00249311
R11378 VSS.n5430 VSS.n5429 0.00249311
R11379 VSS.n5504 VSS.n5503 0.00249311
R11380 VSS.n5531 VSS.n5530 0.00249311
R11381 VSS.n5495 VSS.n5494 0.00249311
R11382 VSS.n5479 VSS.n5478 0.00249311
R11383 VSS.n5472 VSS.n5471 0.00249311
R11384 VSS.n5466 VSS.n5465 0.00249311
R11385 VSS.n5460 VSS.n5459 0.00249311
R11386 VSS.n5454 VSS.n5453 0.00249311
R11387 VSS.n5448 VSS.n5447 0.00249311
R11388 VSS.n5433 VSS.n5432 0.00249311
R11389 VSS.n5442 VSS.n5441 0.00249311
R11390 VSS.n5356 VSS.n5355 0.00249311
R11391 VSS.n5340 VSS.n5339 0.00249311
R11392 VSS.n5334 VSS.n5333 0.00249311
R11393 VSS.n5328 VSS.n5327 0.00249311
R11394 VSS.n5250 VSS.n5249 0.00249311
R11395 VSS.n5324 VSS.n5323 0.00249311
R11396 VSS.n5351 VSS.n5350 0.00249311
R11397 VSS.n5315 VSS.n5314 0.00249311
R11398 VSS.n5299 VSS.n5298 0.00249311
R11399 VSS.n5292 VSS.n5291 0.00249311
R11400 VSS.n5286 VSS.n5285 0.00249311
R11401 VSS.n5280 VSS.n5279 0.00249311
R11402 VSS.n5274 VSS.n5273 0.00249311
R11403 VSS.n5268 VSS.n5267 0.00249311
R11404 VSS.n5253 VSS.n5252 0.00249311
R11405 VSS.n5262 VSS.n5261 0.00249311
R11406 VSS.n10090 VSS.n10089 0.00249311
R11407 VSS.n10074 VSS.n10073 0.00249311
R11408 VSS.n10068 VSS.n10067 0.00249311
R11409 VSS.n10062 VSS.n10061 0.00249311
R11410 VSS.n4577 VSS.n4576 0.00249311
R11411 VSS.n10058 VSS.n10057 0.00249311
R11412 VSS.n10085 VSS.n10084 0.00249311
R11413 VSS.n10049 VSS.n10048 0.00249311
R11414 VSS.n4585 VSS.n4584 0.00249311
R11415 VSS.n4591 VSS.n4590 0.00249311
R11416 VSS.n4597 VSS.n4596 0.00249311
R11417 VSS.n4601 VSS.n4600 0.00249311
R11418 VSS.n3764 VSS.n3763 0.00249311
R11419 VSS.n3807 VSS.n3806 0.00249311
R11420 VSS.n3801 VSS.n3800 0.00249311
R11421 VSS.n3795 VSS.n3794 0.00249311
R11422 VSS.n3768 VSS.n3767 0.00249311
R11423 VSS.n3780 VSS.n3779 0.00249311
R11424 VSS.n3789 VSS.n3788 0.00249311
R11425 VSS.n3774 VSS.n3773 0.00249311
R11426 VSS.n4609 VSS.n4608 0.00249311
R11427 VSS.n4613 VSS.n4612 0.00249311
R11428 VSS.n4619 VSS.n4618 0.00249311
R11429 VSS.n4626 VSS.n4625 0.00249311
R11430 VSS.n6054 VSS.n6053 0.00249311
R11431 VSS.n6060 VSS.n6059 0.00249311
R11432 VSS.n5988 VSS.n5987 0.00249311
R11433 VSS.n6063 VSS.n6062 0.00249311
R11434 VSS.n6071 VSS.n6070 0.00249311
R11435 VSS.n5972 VSS.n5971 0.00249311
R11436 VSS.n5982 VSS.n5981 0.00249311
R11437 VSS.n5976 VSS.n5975 0.00249311
R11438 VSS.n6165 VSS.n6164 0.00249311
R11439 VSS.n6160 VSS.n6159 0.00249311
R11440 VSS.n6175 VSS.n6174 0.00249311
R11441 VSS.n6169 VSS.n6168 0.00249311
R11442 VSS.n11093 VSS.n11092 0.00249311
R11443 VSS.n11105 VSS.n11104 0.00249311
R11444 VSS.n11087 VSS.n11086 0.00249311
R11445 VSS.n11099 VSS.n11098 0.00249311
R11446 VSS.n11136 VSS.n11135 0.00249311
R11447 VSS.n3726 VSS.n3725 0.00249311
R11448 VSS.n3732 VSS.n3731 0.00249311
R11449 VSS.n3736 VSS.n3735 0.00249311
R11450 VSS.n3739 VSS.n3738 0.00249311
R11451 VSS.n3743 VSS.n3742 0.00249311
R11452 VSS.n3749 VSS.n3748 0.00249311
R11453 VSS.n3755 VSS.n3754 0.00249311
R11454 VSS.n11055 VSS.n11054 0.00249311
R11455 VSS.n11051 VSS.n11050 0.00249311
R11456 VSS.n11065 VSS.n11064 0.00249311
R11457 VSS.n11059 VSS.n11058 0.00249311
R11458 VSS.n6389 VSS.n6388 0.00249311
R11459 VSS.n6352 VSS.n6350 0.00249311
R11460 VSS.n6363 VSS.n6362 0.00249311
R11461 VSS.n6359 VSS.n6358 0.00249311
R11462 VSS.n6339 VSS.n6336 0.00249311
R11463 VSS.n6343 VSS.n6335 0.00249311
R11464 VSS.n6402 VSS.n6401 0.00249311
R11465 VSS.n6397 VSS.n6396 0.00249311
R11466 VSS.n11021 VSS.n3839 0.00249311
R11467 VSS.n11020 VSS.n11019 0.00249311
R11468 VSS.n11010 VSS.n11009 0.00249311
R11469 VSS.n11013 VSS.n11012 0.00249311
R11470 VSS.n3861 VSS.n3854 0.00249311
R11471 VSS.n10990 VSS.n10989 0.00249311
R11472 VSS.n3867 VSS.n3866 0.00249311
R11473 VSS.n3871 VSS.n3870 0.00249311
R11474 VSS.n10973 VSS.n10972 0.00249311
R11475 VSS.n10969 VSS.n10968 0.00249311
R11476 VSS.n10980 VSS.n10979 0.00249311
R11477 VSS.n3879 VSS.n3878 0.00249311
R11478 VSS.n10950 VSS.n10949 0.00249311
R11479 VSS.n10914 VSS.n10901 0.00249311
R11480 VSS.n10911 VSS.n10902 0.00249311
R11481 VSS.n10907 VSS.n10903 0.00249311
R11482 VSS.n7335 VSS.n7334 0.00249311
R11483 VSS.n7298 VSS.n7296 0.00249311
R11484 VSS.n7309 VSS.n7308 0.00249311
R11485 VSS.n7305 VSS.n7304 0.00249311
R11486 VSS.n7285 VSS.n7282 0.00249311
R11487 VSS.n7289 VSS.n7281 0.00249311
R11488 VSS.n7348 VSS.n7347 0.00249311
R11489 VSS.n7343 VSS.n7342 0.00249311
R11490 VSS.n10870 VSS.n3907 0.00249311
R11491 VSS.n10869 VSS.n10868 0.00249311
R11492 VSS.n10859 VSS.n10858 0.00249311
R11493 VSS.n10862 VSS.n10861 0.00249311
R11494 VSS.n3980 VSS.n3979 0.00249311
R11495 VSS.n3986 VSS.n3985 0.00249311
R11496 VSS.n3992 VSS.n3991 0.00249311
R11497 VSS.n3996 VSS.n3995 0.00249311
R11498 VSS.n3999 VSS.n3998 0.00249311
R11499 VSS.n4003 VSS.n4002 0.00249311
R11500 VSS.n4009 VSS.n4008 0.00249311
R11501 VSS.n3971 VSS.n3970 0.00249311
R11502 VSS.n4038 VSS.n4037 0.00249311
R11503 VSS.n4034 VSS.n4033 0.00249311
R11504 VSS.n4048 VSS.n4047 0.00249311
R11505 VSS.n4042 VSS.n4041 0.00249311
R11506 VSS.n4144 VSS.n4141 0.00249311
R11507 VSS.n4137 VSS.n4136 0.00249311
R11508 VSS.n4448 VSS.n4135 0.00249311
R11509 VSS.n4148 VSS.n4139 0.00249311
R11510 VSS.n4199 VSS.n4198 0.00249311
R11511 VSS.n4397 VSS.n4396 0.00249311
R11512 VSS.n4393 VSS.n4385 0.00249311
R11513 VSS.n4388 VSS.n4387 0.00249311
R11514 VSS.n4361 VSS.n4202 0.00249311
R11515 VSS.n4374 VSS.n4373 0.00249311
R11516 VSS.n4364 VSS.n4363 0.00249311
R11517 VSS.n4368 VSS.n4367 0.00249311
R11518 VSS.n4336 VSS.n4335 0.00249311
R11519 VSS.n4342 VSS.n4341 0.00249311
R11520 VSS.n4265 VSS.n4264 0.00249311
R11521 VSS.n4258 VSS.n4257 0.00249311
R11522 VSS.n4304 VSS.n4263 0.00249311
R11523 VSS.n4321 VSS.n4320 0.00249311
R11524 VSS.n4317 VSS.n4316 0.00249311
R11525 VSS.n4311 VSS.n4310 0.00249311
R11526 VSS.n4284 VSS.n4282 0.00249311
R11527 VSS.n4280 VSS.n4279 0.00249311
R11528 VSS.n4293 VSS.n4278 0.00249311
R11529 VSS.n4273 VSS.n4272 0.00249311
R11530 VSS.n4347 VSS.n4346 0.00249311
R11531 VSS.n4239 VSS.n4231 0.00249311
R11532 VSS.n4246 VSS.n4238 0.00249311
R11533 VSS.n4243 VSS.n4240 0.00249311
R11534 VSS.n4216 VSS.n4215 0.00249311
R11535 VSS.n4221 VSS.n4213 0.00249311
R11536 VSS.n4210 VSS.n4195 0.00249311
R11537 VSS.n4404 VSS.n4195 0.00249311
R11538 VSS.n4220 VSS.n4219 0.00249311
R11539 VSS.n4170 VSS.n4169 0.00249311
R11540 VSS.n4176 VSS.n4175 0.00249311
R11541 VSS.n4172 VSS.n4163 0.00249311
R11542 VSS.n4408 VSS.n4407 0.00249311
R11543 VSS.n4417 VSS.n4416 0.00249311
R11544 VSS.n4430 VSS.n4429 0.00249311
R11545 VSS.n4427 VSS.n4426 0.00249311
R11546 VSS.n4422 VSS.n4421 0.00249311
R11547 VSS.n4123 VSS.n4121 0.00249311
R11548 VSS.n4120 VSS.n4109 0.00249311
R11549 VSS.n10779 VSS.n10778 0.00249311
R11550 VSS.n4130 VSS.n4129 0.00249311
R11551 VSS.n10766 VSS.n4134 0.00249311
R11552 VSS.n10763 VSS.n10749 0.00249311
R11553 VSS.n10751 VSS.n10750 0.00249311
R11554 VSS.n10755 VSS.n10753 0.00249311
R11555 VSS.n1286 VSS.n1285 0.00249311
R11556 VSS.n1280 VSS.n1279 0.00249311
R11557 VSS.n1274 VSS.n1273 0.00249311
R11558 VSS.n1248 VSS.n1247 0.00249311
R11559 VSS.n685 VSS.n684 0.00249311
R11560 VSS.n785 VSS.n784 0.00249311
R11561 VSS.n779 VSS.n778 0.00249311
R11562 VSS.n663 VSS.n662 0.00249311
R11563 VSS.n654 VSS.n653 0.00249311
R11564 VSS.n679 VSS.n678 0.00249311
R11565 VSS.n673 VSS.n672 0.00249311
R11566 VSS.n667 VSS.n666 0.00249311
R11567 VSS.n1294 VSS.n1293 0.00249311
R11568 VSS.n1263 VSS.n1262 0.00249311
R11569 VSS.n1257 VSS.n1256 0.00249311
R11570 VSS.n1251 VSS.n1250 0.00249311
R11571 VSS.n1215 VSS.n1214 0.00249311
R11572 VSS.n1218 VSS.n1217 0.00249311
R11573 VSS.n1224 VSS.n1223 0.00249311
R11574 VSS.n1230 VSS.n1229 0.00249311
R11575 VSS.n1043 VSS.n1042 0.00249311
R11576 VSS.n1036 VSS.n1035 0.00249311
R11577 VSS.n1030 VSS.n1029 0.00249311
R11578 VSS.n1024 VSS.n1023 0.00249311
R11579 VSS.n1018 VSS.n1017 0.00249311
R11580 VSS.n1012 VSS.n1011 0.00249311
R11581 VSS.n997 VSS.n996 0.00249311
R11582 VSS.n1006 VSS.n1005 0.00249311
R11583 VSS.n1347 VSS.n1346 0.00249311
R11584 VSS.n1211 VSS.n1210 0.00249311
R11585 VSS.n1205 VSS.n1204 0.00249311
R11586 VSS.n1199 VSS.n1198 0.00249311
R11587 VSS.n963 VSS.n962 0.00249311
R11588 VSS.n966 VSS.n965 0.00249311
R11589 VSS.n972 VSS.n971 0.00249311
R11590 VSS.n978 VSS.n977 0.00249311
R11591 VSS.n14317 VSS.n14316 0.00249311
R11592 VSS.n14312 VSS.n14311 0.00249311
R11593 VSS.n14327 VSS.n14326 0.00249311
R11594 VSS.n14321 VSS.n14320 0.00249311
R11595 VSS.n581 VSS.n580 0.00249311
R11596 VSS.n14221 VSS.n14220 0.00249311
R11597 VSS.n14217 VSS.n14209 0.00249311
R11598 VSS.n14212 VSS.n14211 0.00249311
R11599 VSS.n14231 VSS.n547 0.00249311
R11600 VSS.n559 VSS.n546 0.00249311
R11601 VSS.n566 VSS.n558 0.00249311
R11602 VSS.n561 VSS.n560 0.00249311
R11603 VSS.n10689 VSS.n10688 0.00249311
R11604 VSS.n10654 VSS.n10653 0.00249311
R11605 VSS.n10683 VSS.n10682 0.00249311
R11606 VSS.n10677 VSS.n10676 0.00249311
R11607 VSS.n14264 VSS.n14263 0.00249311
R11608 VSS.n14270 VSS.n14269 0.00249311
R11609 VSS.n509 VSS.n508 0.00249311
R11610 VSS.n518 VSS.n517 0.00249311
R11611 VSS.n14258 VSS.n14257 0.00249311
R11612 VSS.n534 VSS.n533 0.00249311
R11613 VSS.n528 VSS.n527 0.00249311
R11614 VSS.n522 VSS.n521 0.00249311
R11615 VSS.n10702 VSS.n10701 0.00249311
R11616 VSS.n10669 VSS.n10668 0.00249311
R11617 VSS.n10663 VSS.n10662 0.00249311
R11618 VSS.n10657 VSS.n10656 0.00249311
R11619 VSS.n14203 VSS.n586 0.00249311
R11620 VSS.n591 VSS.n585 0.00249311
R11621 VSS.n598 VSS.n590 0.00249311
R11622 VSS.n593 VSS.n592 0.00249311
R11623 VSS.n1137 VSS.n936 0.00249311
R11624 VSS.n1145 VSS.n1144 0.00249311
R11625 VSS.n934 VSS.n933 0.00249311
R11626 VSS.n1141 VSS.n1140 0.00249311
R11627 VSS.n928 VSS.n911 0.00249311
R11628 VSS.n1153 VSS.n912 0.00249311
R11629 VSS.n926 VSS.n925 0.00249311
R11630 VSS.n921 VSS.n920 0.00249311
R11631 VSS.n14176 VSS.n605 0.00249311
R11632 VSS.n14194 VSS.n14193 0.00249311
R11633 VSS.n14190 VSS.n14189 0.00249311
R11634 VSS.n14186 VSS.n14181 0.00249311
R11635 VSS.n12449 VSS.n12448 0.00249311
R11636 VSS.n12443 VSS.n12442 0.00249311
R11637 VSS.n12437 VSS.n12436 0.00249311
R11638 VSS.n12393 VSS.n12392 0.00249311
R11639 VSS.n12415 VSS.n12398 0.00249311
R11640 VSS.n12413 VSS.n12399 0.00249311
R11641 VSS.n12409 VSS.n12400 0.00249311
R11642 VSS.n12405 VSS.n12401 0.00249311
R11643 VSS.n2498 VSS.n2496 0.00249311
R11644 VSS.n2497 VSS.n2495 0.00249311
R11645 VSS.n13037 VSS.n13036 0.00249311
R11646 VSS.n13033 VSS.n13032 0.00249311
R11647 VSS.n2541 VSS.n2540 0.00249311
R11648 VSS.n2537 VSS.n2536 0.00249311
R11649 VSS.n2533 VSS.n2485 0.00249311
R11650 VSS.n2544 VSS.n2543 0.00249311
R11651 VSS.n13054 VSS.n2463 0.00249311
R11652 VSS.n2464 VSS.n2462 0.00249311
R11653 VSS.n2474 VSS.n2467 0.00249311
R11654 VSS.n2469 VSS.n2468 0.00249311
R11655 VSS.n2450 VSS.n2449 0.00249311
R11656 VSS.n2442 VSS.n2394 0.00249311
R11657 VSS.n2439 VSS.n2431 0.00249311
R11658 VSS.n2436 VSS.n2435 0.00249311
R11659 VSS.n13098 VSS.n2371 0.00249311
R11660 VSS.n2355 VSS.n2353 0.00249311
R11661 VSS.n2354 VSS.n2352 0.00249311
R11662 VSS.n2367 VSS.n2365 0.00249311
R11663 VSS.n2380 VSS.n2379 0.00249311
R11664 VSS.n2388 VSS.n2387 0.00249311
R11665 VSS.n2374 VSS.n2373 0.00249311
R11666 VSS.n2384 VSS.n2376 0.00249311
R11667 VSS.n13070 VSS.n2455 0.00249311
R11668 VSS.n13088 VSS.n13087 0.00249311
R11669 VSS.n13084 VSS.n13083 0.00249311
R11670 VSS.n13080 VSS.n13075 0.00249311
R11671 VSS.n13134 VSS.n1912 0.00249311
R11672 VSS.n1914 VSS.n1913 0.00249311
R11673 VSS.n1922 VSS.n1921 0.00249311
R11674 VSS.n1926 VSS.n1925 0.00249311
R11675 VSS.n2328 VSS.n1946 0.00249311
R11676 VSS.n2336 VSS.n2335 0.00249311
R11677 VSS.n1944 VSS.n1943 0.00249311
R11678 VSS.n2332 VSS.n2331 0.00249311
R11679 VSS.n2281 VSS.n1933 0.00249311
R11680 VSS.n2293 VSS.n2292 0.00249311
R11681 VSS.n2289 VSS.n2288 0.00249311
R11682 VSS.n2285 VSS.n2282 0.00249311
R11683 VSS.n2349 VSS.n2348 0.00249311
R11684 VSS.n13123 VSS.n13108 0.00249311
R11685 VSS.n13110 VSS.n13109 0.00249311
R11686 VSS.n13114 VSS.n13112 0.00249311
R11687 VSS.n14164 VSS.n14163 0.00249311
R11688 VSS.n14169 VSS.n14161 0.00249311
R11689 VSS.n14158 VSS.n577 0.00249311
R11690 VSS.n14228 VSS.n577 0.00249311
R11691 VSS.n14168 VSS.n14167 0.00249311
R11692 VSS.n2405 VSS.n2404 0.00249311
R11693 VSS.n2417 VSS.n2416 0.00249311
R11694 VSS.n2414 VSS.n2413 0.00249311
R11695 VSS.n2410 VSS.n2407 0.00249311
R11696 VSS.n896 VSS.n885 0.00249311
R11697 VSS.n897 VSS.n895 0.00249311
R11698 VSS.n906 VSS.n905 0.00249311
R11699 VSS.n903 VSS.n902 0.00249311
R11700 VSS.n939 VSS.n938 0.00249311
R11701 VSS.n945 VSS.n944 0.00249311
R11702 VSS.n949 VSS.n948 0.00249311
R11703 VSS.n951 VSS.n950 0.00249311
R11704 VSS.n1396 VSS.n863 0.00249311
R11705 VSS.n865 VSS.n864 0.00249311
R11706 VSS.n873 VSS.n872 0.00249311
R11707 VSS.n877 VSS.n876 0.00249311
R11708 VSS.n1376 VSS.n1374 0.00249311
R11709 VSS.n1383 VSS.n1382 0.00249311
R11710 VSS.n1386 VSS.n1370 0.00249311
R11711 VSS.n1371 VSS.n1170 0.00249311
R11712 VSS.n1371 VSS.n879 0.00249311
R11713 VSS.n1108 VSS.n1107 0.00249311
R11714 VSS.n1091 VSS.n1090 0.00249311
R11715 VSS.n1097 VSS.n1096 0.00249311
R11716 VSS.n1101 VSS.n1100 0.00249311
R11717 VSS.n14298 VSS.n14297 0.00249311
R11718 VSS.n14292 VSS.n14291 0.00249311
R11719 VSS.n14282 VSS.n14281 0.00249311
R11720 VSS.n14286 VSS.n14285 0.00249311
R11721 VSS.n1565 VSS.n1564 0.00249311
R11722 VSS.n1558 VSS.n1557 0.00249311
R11723 VSS.n1552 VSS.n1551 0.00249311
R11724 VSS.n1546 VSS.n1545 0.00249311
R11725 VSS.n1540 VSS.n1539 0.00249311
R11726 VSS.n1534 VSS.n1533 0.00249311
R11727 VSS.n1519 VSS.n1518 0.00249311
R11728 VSS.n1528 VSS.n1527 0.00249311
R11729 VSS.n13855 VSS.n13854 0.00249311
R11730 VSS.n13724 VSS.n13723 0.00249311
R11731 VSS.n13730 VSS.n13729 0.00249311
R11732 VSS.n13734 VSS.n13733 0.00249311
R11733 VSS.n13707 VSS.n13706 0.00249311
R11734 VSS.n13740 VSS.n13739 0.00249311
R11735 VSS.n13849 VSS.n13848 0.00249311
R11736 VSS.n13705 VSS.n13704 0.00249311
R11737 VSS.n13853 VSS.n13705 0.00249311
R11738 VSS.n13805 VSS.n13804 0.00249311
R11739 VSS.n13798 VSS.n13797 0.00249311
R11740 VSS.n13792 VSS.n13791 0.00249311
R11741 VSS.n13786 VSS.n13785 0.00249311
R11742 VSS.n13780 VSS.n13779 0.00249311
R11743 VSS.n13774 VSS.n13773 0.00249311
R11744 VSS.n13759 VSS.n13758 0.00249311
R11745 VSS.n13768 VSS.n13767 0.00249311
R11746 VSS.n13390 VSS.n13389 0.00249311
R11747 VSS.n13261 VSS.n13260 0.00249311
R11748 VSS.n13267 VSS.n13266 0.00249311
R11749 VSS.n13271 VSS.n13270 0.00249311
R11750 VSS.n13244 VSS.n13243 0.00249311
R11751 VSS.n13277 VSS.n13276 0.00249311
R11752 VSS.n13384 VSS.n13383 0.00249311
R11753 VSS.n13242 VSS.n13241 0.00249311
R11754 VSS.n13388 VSS.n13242 0.00249311
R11755 VSS.n1484 VSS.n1483 0.00249311
R11756 VSS.n1487 VSS.n1486 0.00249311
R11757 VSS.n1493 VSS.n1492 0.00249311
R11758 VSS.n1499 VSS.n1498 0.00249311
R11759 VSS.n758 VSS.n757 0.00249311
R11760 VSS.n751 VSS.n750 0.00249311
R11761 VSS.n745 VSS.n744 0.00249311
R11762 VSS.n739 VSS.n738 0.00249311
R11763 VSS.n733 VSS.n732 0.00249311
R11764 VSS.n727 VSS.n726 0.00249311
R11765 VSS.n712 VSS.n711 0.00249311
R11766 VSS.n721 VSS.n720 0.00249311
R11767 VSS.n1618 VSS.n1617 0.00249311
R11768 VSS.n1480 VSS.n1479 0.00249311
R11769 VSS.n1474 VSS.n1473 0.00249311
R11770 VSS.n1468 VSS.n1467 0.00249311
R11771 VSS.n14113 VSS.n629 0.00249311
R11772 VSS.n14118 VSS.n14117 0.00249311
R11773 VSS.n647 VSS.n646 0.00249311
R11774 VSS.n642 VSS.n641 0.00249311
R11775 VSS.n1445 VSS.n1444 0.00249311
R11776 VSS.n1446 VSS.n1442 0.00249311
R11777 VSS.n1454 VSS.n1453 0.00249311
R11778 VSS.n1455 VSS.n652 0.00249311
R11779 VSS.n1688 VSS.n1687 0.00249311
R11780 VSS.n1691 VSS.n1674 0.00249311
R11781 VSS.n1683 VSS.n1675 0.00249311
R11782 VSS.n1679 VSS.n1676 0.00249311
R11783 VSS.n14093 VSS.n14091 0.00249311
R11784 VSS.n14100 VSS.n14099 0.00249311
R11785 VSS.n14103 VSS.n14087 0.00249311
R11786 VSS.n14088 VSS.n1463 0.00249311
R11787 VSS.n14088 VSS.n650 0.00249311
R11788 VSS.n13681 VSS.n13677 0.00249311
R11789 VSS.n13689 VSS.n13688 0.00249311
R11790 VSS.n13692 VSS.n13671 0.00249311
R11791 VSS.n13692 VSS.n1661 0.00249311
R11792 VSS.n13679 VSS.n13675 0.00249311
R11793 VSS.n1671 VSS.n1663 0.00249311
R11794 VSS.n14074 VSS.n14073 0.00249311
R11795 VSS.n14064 VSS.n14063 0.00249311
R11796 VSS.n14068 VSS.n14067 0.00249311
R11797 VSS.n1654 VSS.n1650 0.00249311
R11798 VSS.n1651 VSS.n1642 0.00249311
R11799 VSS.n14082 VSS.n14081 0.00249311
R11800 VSS.n1665 VSS.n1664 0.00249311
R11801 VSS.n13700 VSS.n13699 0.00249311
R11802 VSS.n13667 VSS.n13653 0.00249311
R11803 VSS.n13663 VSS.n13654 0.00249311
R11804 VSS.n13659 VSS.n13655 0.00249311
R11805 VSS.n13904 VSS.n13205 0.00249311
R11806 VSS.n13207 VSS.n13206 0.00249311
R11807 VSS.n13215 VSS.n13214 0.00249311
R11808 VSS.n13219 VSS.n13218 0.00249311
R11809 VSS.n13239 VSS.n13237 0.00249311
R11810 VSS.n13238 VSS.n13236 0.00249311
R11811 VSS.n13635 VSS.n13634 0.00249311
R11812 VSS.n13631 VSS.n13630 0.00249311
R11813 VSS.n13540 VSS.n13539 0.00249311
R11814 VSS.n13536 VSS.n13535 0.00249311
R11815 VSS.n13532 VSS.n13226 0.00249311
R11816 VSS.n13543 VSS.n13542 0.00249311
R11817 VSS.n13884 VSS.n13882 0.00249311
R11818 VSS.n13880 VSS.n13879 0.00249311
R11819 VSS.n13893 VSS.n13878 0.00249311
R11820 VSS.n13650 VSS.n13649 0.00249311
R11821 VSS.n828 VSS.n825 0.00249311
R11822 VSS.n831 VSS.n824 0.00249311
R11823 VSS.n816 VSS.n814 0.00249311
R11824 VSS.n817 VSS.n815 0.00249311
R11825 VSS.n1409 VSS.n844 0.00249311
R11826 VSS.n846 VSS.n845 0.00249311
R11827 VSS.n858 VSS.n857 0.00249311
R11828 VSS.n854 VSS.n851 0.00249311
R11829 VSS.n1181 VSS.n1180 0.00249311
R11830 VSS.n1185 VSS.n1184 0.00249311
R11831 VSS.n1188 VSS.n1173 0.00249311
R11832 VSS.n1192 VSS.n1174 0.00249311
R11833 VSS.n1433 VSS.n1432 0.00249311
R11834 VSS.n1429 VSS.n1428 0.00249311
R11835 VSS.n1425 VSS.n1417 0.00249311
R11836 VSS.n1420 VSS.n1419 0.00249311
R11837 VSS.n2197 VSS.n2196 0.00249311
R11838 VSS.n2192 VSS.n2056 0.00249311
R11839 VSS.n2209 VSS.n2208 0.00249311
R11840 VSS.n2209 VSS.n2005 0.00249311
R11841 VSS.n2200 VSS.n2190 0.00249311
R11842 VSS.n2243 VSS.n1984 0.00249311
R11843 VSS.n2248 VSS.n2247 0.00249311
R11844 VSS.n2002 VSS.n2001 0.00249311
R11845 VSS.n1997 VSS.n1996 0.00249311
R11846 VSS.n2039 VSS.n2038 0.00249311
R11847 VSS.n2040 VSS.n2036 0.00249311
R11848 VSS.n2048 VSS.n2047 0.00249311
R11849 VSS.n2049 VSS.n2007 0.00249311
R11850 VSS.n2233 VSS.n2213 0.00249311
R11851 VSS.n2232 VSS.n2217 0.00249311
R11852 VSS.n2219 VSS.n2218 0.00249311
R11853 VSS.n2223 VSS.n2221 0.00249311
R11854 VSS.n2111 VSS.n2108 0.00249311
R11855 VSS.n2121 VSS.n2120 0.00249311
R11856 VSS.n2125 VSS.n2124 0.00249311
R11857 VSS.n2125 VSS.n2080 0.00249311
R11858 VSS.n2117 VSS.n2116 0.00249311
R11859 VSS.n2178 VSS.n2059 0.00249311
R11860 VSS.n2183 VSS.n2182 0.00249311
R11861 VSS.n2077 VSS.n2076 0.00249311
R11862 VSS.n2072 VSS.n2071 0.00249311
R11863 VSS.n2088 VSS.n2087 0.00249311
R11864 VSS.n2089 VSS.n2085 0.00249311
R11865 VSS.n2097 VSS.n2096 0.00249311
R11866 VSS.n2098 VSS.n2082 0.00249311
R11867 VSS.n2168 VSS.n2129 0.00249311
R11868 VSS.n2167 VSS.n2152 0.00249311
R11869 VSS.n2154 VSS.n2153 0.00249311
R11870 VSS.n2158 VSS.n2156 0.00249311
R11871 VSS.n12660 VSS.n12659 0.00249311
R11872 VSS.n12655 VSS.n12647 0.00249311
R11873 VSS.n12651 VSS.n12650 0.00249311
R11874 VSS.n12650 VSS.n1849 0.00249311
R11875 VSS.n12663 VSS.n12648 0.00249311
R11876 VSS.n1867 VSS.n1856 0.00249311
R11877 VSS.n1868 VSS.n1866 0.00249311
R11878 VSS.n1877 VSS.n1876 0.00249311
R11879 VSS.n1874 VSS.n1873 0.00249311
R11880 VSS.n2136 VSS.n2135 0.00249311
R11881 VSS.n2140 VSS.n2139 0.00249311
R11882 VSS.n2147 VSS.n2146 0.00249311
R11883 VSS.n2144 VSS.n2143 0.00249311
R11884 VSS.n13198 VSS.n13197 0.00249311
R11885 VSS.n1847 VSS.n1832 0.00249311
R11886 VSS.n1844 VSS.n1837 0.00249311
R11887 VSS.n1841 VSS.n1838 0.00249311
R11888 VSS.n12688 VSS.n12670 0.00249311
R11889 VSS.n12685 VSS.n12671 0.00249311
R11890 VSS.n12681 VSS.n12672 0.00249311
R11891 VSS.n12677 VSS.n12673 0.00249311
R11892 VSS.n13932 VSS.n1792 0.00249311
R11893 VSS.n1776 VSS.n1774 0.00249311
R11894 VSS.n1775 VSS.n1773 0.00249311
R11895 VSS.n1788 VSS.n1786 0.00249311
R11896 VSS.n1801 VSS.n1800 0.00249311
R11897 VSS.n1809 VSS.n1808 0.00249311
R11898 VSS.n1795 VSS.n1794 0.00249311
R11899 VSS.n1805 VSS.n1797 0.00249311
R11900 VSS.n1824 VSS.n1822 0.00249311
R11901 VSS.n1825 VSS.n1818 0.00249311
R11902 VSS.n13918 VSS.n1817 0.00249311
R11903 VSS.n13922 VSS.n1815 0.00249311
R11904 VSS.n2029 VSS.n2012 0.00249311
R11905 VSS.n2022 VSS.n2013 0.00249311
R11906 VSS.n2018 VSS.n2014 0.00249311
R11907 VSS.n2026 VSS.n2011 0.00249311
R11908 VSS.n2279 VSS.n1974 0.00249311
R11909 VSS.n2313 VSS.n2312 0.00249311
R11910 VSS.n2309 VSS.n2301 0.00249311
R11911 VSS.n2304 VSS.n2303 0.00249311
R11912 VSS.n1952 VSS.n1950 0.00249311
R11913 VSS.n1951 VSS.n1949 0.00249311
R11914 VSS.n1963 VSS.n1956 0.00249311
R11915 VSS.n1958 VSS.n1957 0.00249311
R11916 VSS.n2271 VSS.n1981 0.00249311
R11917 VSS.n2270 VSS.n2255 0.00249311
R11918 VSS.n2257 VSS.n2256 0.00249311
R11919 VSS.n2261 VSS.n2259 0.00249311
R11920 VSS.n12983 VSS.n2563 0.00249311
R11921 VSS.n12988 VSS.n12987 0.00249311
R11922 VSS.n2581 VSS.n2580 0.00249311
R11923 VSS.n2576 VSS.n2575 0.00249311
R11924 VSS.n2646 VSS.n2645 0.00249311
R11925 VSS.n2647 VSS.n2643 0.00249311
R11926 VSS.n2655 VSS.n2654 0.00249311
R11927 VSS.n2656 VSS.n2586 0.00249311
R11928 VSS.n2718 VSS.n2700 0.00249311
R11929 VSS.n2715 VSS.n2701 0.00249311
R11930 VSS.n2711 VSS.n2702 0.00249311
R11931 VSS.n2707 VSS.n2703 0.00249311
R11932 VSS.n12973 VSS.n2663 0.00249311
R11933 VSS.n12959 VSS.n12958 0.00249311
R11934 VSS.n12963 VSS.n12961 0.00249311
R11935 VSS.n12972 VSS.n12957 0.00249311
R11936 VSS.n2698 VSS.n2690 0.00249311
R11937 VSS.n12944 VSS.n12943 0.00249311
R11938 VSS.n12934 VSS.n12933 0.00249311
R11939 VSS.n12938 VSS.n12937 0.00249311
R11940 VSS.n2681 VSS.n2677 0.00249311
R11941 VSS.n2678 VSS.n2669 0.00249311
R11942 VSS.n12952 VSS.n12951 0.00249311
R11943 VSS.n2692 VSS.n2691 0.00249311
R11944 VSS.n2809 VSS.n2788 0.00249311
R11945 VSS.n2805 VSS.n2790 0.00249311
R11946 VSS.n2798 VSS.n2793 0.00249311
R11947 VSS.n2797 VSS.n2795 0.00249311
R11948 VSS.n2818 VSS.n2817 0.00249311
R11949 VSS.n2781 VSS.n2772 0.00249311
R11950 VSS.n2776 VSS.n2773 0.00249311
R11951 VSS.n2785 VSS.n2771 0.00249311
R11952 VSS.n12906 VSS.n2744 0.00249311
R11953 VSS.n12911 VSS.n12910 0.00249311
R11954 VSS.n2762 VSS.n2761 0.00249311
R11955 VSS.n2757 VSS.n2756 0.00249311
R11956 VSS.n2827 VSS.n2826 0.00249311
R11957 VSS.n2828 VSS.n2824 0.00249311
R11958 VSS.n2836 VSS.n2835 0.00249311
R11959 VSS.n2837 VSS.n2767 0.00249311
R11960 VSS.n2898 VSS.n2880 0.00249311
R11961 VSS.n2895 VSS.n2881 0.00249311
R11962 VSS.n2891 VSS.n2882 0.00249311
R11963 VSS.n2887 VSS.n2883 0.00249311
R11964 VSS.n12896 VSS.n2844 0.00249311
R11965 VSS.n12882 VSS.n12881 0.00249311
R11966 VSS.n12886 VSS.n12884 0.00249311
R11967 VSS.n12895 VSS.n12880 0.00249311
R11968 VSS.n12622 VSS.n12618 0.00249311
R11969 VSS.n12630 VSS.n12629 0.00249311
R11970 VSS.n12633 VSS.n3055 0.00249311
R11971 VSS.n12633 VSS.n2868 0.00249311
R11972 VSS.n12620 VSS.n3059 0.00249311
R11973 VSS.n2878 VSS.n2870 0.00249311
R11974 VSS.n12867 VSS.n12866 0.00249311
R11975 VSS.n12857 VSS.n12856 0.00249311
R11976 VSS.n12861 VSS.n12860 0.00249311
R11977 VSS.n2861 VSS.n2857 0.00249311
R11978 VSS.n2858 VSS.n2849 0.00249311
R11979 VSS.n12875 VSS.n12874 0.00249311
R11980 VSS.n2872 VSS.n2871 0.00249311
R11981 VSS.n12641 VSS.n12640 0.00249311
R11982 VSS.n3051 VSS.n3037 0.00249311
R11983 VSS.n3047 VSS.n3038 0.00249311
R11984 VSS.n3043 VSS.n3039 0.00249311
R11985 VSS.n3079 VSS.n3061 0.00249311
R11986 VSS.n3076 VSS.n3062 0.00249311
R11987 VSS.n3072 VSS.n3063 0.00249311
R11988 VSS.n3068 VSS.n3064 0.00249311
R11989 VSS.n12727 VSS.n2970 0.00249311
R11990 VSS.n2954 VSS.n2952 0.00249311
R11991 VSS.n2953 VSS.n2951 0.00249311
R11992 VSS.n2966 VSS.n2964 0.00249311
R11993 VSS.n3006 VSS.n3005 0.00249311
R11994 VSS.n3014 VSS.n3013 0.00249311
R11995 VSS.n2973 VSS.n2972 0.00249311
R11996 VSS.n3010 VSS.n3002 0.00249311
R11997 VSS.n3029 VSS.n3027 0.00249311
R11998 VSS.n3030 VSS.n3023 0.00249311
R11999 VSS.n12713 VSS.n3022 0.00249311
R12000 VSS.n12717 VSS.n3020 0.00249311
R12001 VSS.n2636 VSS.n2592 0.00249311
R12002 VSS.n2602 VSS.n2593 0.00249311
R12003 VSS.n2598 VSS.n2594 0.00249311
R12004 VSS.n2606 VSS.n2591 0.00249311
R12005 VSS.n2530 VSS.n2526 0.00249311
R12006 VSS.n13018 VSS.n13017 0.00249311
R12007 VSS.n13014 VSS.n13006 0.00249311
R12008 VSS.n13009 VSS.n13008 0.00249311
R12009 VSS.n2504 VSS.n2502 0.00249311
R12010 VSS.n2503 VSS.n2501 0.00249311
R12011 VSS.n2515 VSS.n2508 0.00249311
R12012 VSS.n2510 VSS.n2509 0.00249311
R12013 VSS.n2626 VSS.n2609 0.00249311
R12014 VSS.n2625 VSS.n2610 0.00249311
R12015 VSS.n2612 VSS.n2611 0.00249311
R12016 VSS.n2616 VSS.n2614 0.00249311
R12017 VSS.n11571 VSS.n11570 0.00249311
R12018 VSS.n11672 VSS.n11671 0.00249311
R12019 VSS.n11666 VSS.n11665 0.00249311
R12020 VSS.n11660 VSS.n11659 0.00249311
R12021 VSS.n11654 VSS.n11653 0.00249311
R12022 VSS.n11648 VSS.n11647 0.00249311
R12023 VSS.n11642 VSS.n11641 0.00249311
R12024 VSS.n11580 VSS.n11579 0.00249311
R12025 VSS.n12258 VSS.n12257 0.00249311
R12026 VSS.n12242 VSS.n12241 0.00249311
R12027 VSS.n12236 VSS.n12235 0.00249311
R12028 VSS.n12230 VSS.n12229 0.00249311
R12029 VSS.n12210 VSS.n12209 0.00249311
R12030 VSS.n12226 VSS.n12225 0.00249311
R12031 VSS.n12253 VSS.n12252 0.00249311
R12032 VSS.n12217 VSS.n12216 0.00249311
R12033 VSS.n11695 VSS.n11694 0.00249311
R12034 VSS.n11741 VSS.n11740 0.00249311
R12035 VSS.n11735 VSS.n11734 0.00249311
R12036 VSS.n11729 VSS.n11728 0.00249311
R12037 VSS.n11723 VSS.n11722 0.00249311
R12038 VSS.n11717 VSS.n11716 0.00249311
R12039 VSS.n11711 VSS.n11710 0.00249311
R12040 VSS.n11704 VSS.n11703 0.00249311
R12041 VSS.n12151 VSS.n12150 0.00249311
R12042 VSS.n12135 VSS.n12134 0.00249311
R12043 VSS.n12129 VSS.n12128 0.00249311
R12044 VSS.n12123 VSS.n12122 0.00249311
R12045 VSS.n12046 VSS.n12045 0.00249311
R12046 VSS.n12119 VSS.n12118 0.00249311
R12047 VSS.n12146 VSS.n12145 0.00249311
R12048 VSS.n12110 VSS.n12109 0.00249311
R12049 VSS.n12094 VSS.n12093 0.00249311
R12050 VSS.n12087 VSS.n12086 0.00249311
R12051 VSS.n12081 VSS.n12080 0.00249311
R12052 VSS.n12075 VSS.n12074 0.00249311
R12053 VSS.n12069 VSS.n12068 0.00249311
R12054 VSS.n12063 VSS.n12062 0.00249311
R12055 VSS.n12048 VSS.n12047 0.00249311
R12056 VSS.n12057 VSS.n12056 0.00249311
R12057 VSS.n11983 VSS.n11982 0.00249311
R12058 VSS.n11967 VSS.n11966 0.00249311
R12059 VSS.n11961 VSS.n11960 0.00249311
R12060 VSS.n11955 VSS.n11954 0.00249311
R12061 VSS.n11935 VSS.n11934 0.00249311
R12062 VSS.n11951 VSS.n11950 0.00249311
R12063 VSS.n11978 VSS.n11977 0.00249311
R12064 VSS.n11942 VSS.n11941 0.00249311
R12065 VSS.n11827 VSS.n11826 0.00249311
R12066 VSS.n11873 VSS.n11872 0.00249311
R12067 VSS.n11867 VSS.n11866 0.00249311
R12068 VSS.n11861 VSS.n11860 0.00249311
R12069 VSS.n11855 VSS.n11854 0.00249311
R12070 VSS.n11849 VSS.n11848 0.00249311
R12071 VSS.n11843 VSS.n11842 0.00249311
R12072 VSS.n11836 VSS.n11835 0.00249311
R12073 VSS.n3555 VSS.n3554 0.00249311
R12074 VSS.n3539 VSS.n3538 0.00249311
R12075 VSS.n3533 VSS.n3532 0.00249311
R12076 VSS.n3527 VSS.n3526 0.00249311
R12077 VSS.n3450 VSS.n3449 0.00249311
R12078 VSS.n3523 VSS.n3522 0.00249311
R12079 VSS.n3550 VSS.n3549 0.00249311
R12080 VSS.n3514 VSS.n3513 0.00249311
R12081 VSS.n3498 VSS.n3497 0.00249311
R12082 VSS.n3491 VSS.n3490 0.00249311
R12083 VSS.n3485 VSS.n3484 0.00249311
R12084 VSS.n3479 VSS.n3478 0.00249311
R12085 VSS.n3473 VSS.n3472 0.00249311
R12086 VSS.n3467 VSS.n3466 0.00249311
R12087 VSS.n3452 VSS.n3451 0.00249311
R12088 VSS.n3461 VSS.n3460 0.00249311
R12089 VSS.n12591 VSS.n12590 0.00249311
R12090 VSS.n3114 VSS.n3113 0.00249311
R12091 VSS.n3108 VSS.n3107 0.00249311
R12092 VSS.n3102 VSS.n3101 0.00249311
R12093 VSS.n3087 VSS.n3086 0.00249311
R12094 VSS.n3098 VSS.n3097 0.00249311
R12095 VSS.n12602 VSS.n12601 0.00249311
R12096 VSS.n3089 VSS.n3088 0.00249311
R12097 VSS.n3166 VSS.n3165 0.00249311
R12098 VSS.n3125 VSS.n3124 0.00249311
R12099 VSS.n3131 VSS.n3130 0.00249311
R12100 VSS.n3135 VSS.n3134 0.00249311
R12101 VSS.n3226 VSS.n3225 0.00249311
R12102 VSS.n3257 VSS.n3256 0.00249311
R12103 VSS.n3263 VSS.n3262 0.00249311
R12104 VSS.n3217 VSS.n3216 0.00249311
R12105 VSS.n3249 VSS.n3248 0.00249311
R12106 VSS.n3242 VSS.n3241 0.00249311
R12107 VSS.n3236 VSS.n3235 0.00249311
R12108 VSS.n3230 VSS.n3229 0.00249311
R12109 VSS.n3143 VSS.n3142 0.00249311
R12110 VSS.n3147 VSS.n3146 0.00249311
R12111 VSS.n3153 VSS.n3152 0.00249311
R12112 VSS.n3162 VSS.n3161 0.00249311
R12113 VSS.n11631 VSS.n11630 0.00249311
R12114 VSS.n11610 VSS.n11609 0.00249311
R12115 VSS.n11603 VSS.n11602 0.00249311
R12116 VSS.n11613 VSS.n11612 0.00249311
R12117 VSS.n11621 VSS.n11620 0.00249311
R12118 VSS.n11597 VSS.n11596 0.00249311
R12119 VSS.n11591 VSS.n11590 0.00249311
R12120 VSS.n11585 VSS.n11584 0.00249311
R12121 VSS.n12370 VSS.n12369 0.00249311
R12122 VSS.n12366 VSS.n12365 0.00249311
R12123 VSS.n12380 VSS.n12379 0.00249311
R12124 VSS.n12374 VSS.n12373 0.00249311
R12125 VSS.n2978 VSS.n2976 0.00249311
R12126 VSS.n2995 VSS.n2994 0.00249311
R12127 VSS.n2991 VSS.n2990 0.00249311
R12128 VSS.n2985 VSS.n2984 0.00249311
R12129 VSS.n12741 VSS.n12738 0.00249311
R12130 VSS.n12745 VSS.n12737 0.00249311
R12131 VSS.n2948 VSS.n2947 0.00249311
R12132 VSS.n12755 VSS.n2946 0.00249311
R12133 VSS.n12775 VSS.n12761 0.00249311
R12134 VSS.n12774 VSS.n12773 0.00249311
R12135 VSS.n12764 VSS.n12763 0.00249311
R12136 VSS.n12767 VSS.n12766 0.00249311
R12137 VSS.n13969 VSS.n1760 0.00249311
R12138 VSS.n13986 VSS.n13985 0.00249311
R12139 VSS.n13982 VSS.n13981 0.00249311
R12140 VSS.n13976 VSS.n13975 0.00249311
R12141 VSS.n13949 VSS.n13947 0.00249311
R12142 VSS.n13945 VSS.n13944 0.00249311
R12143 VSS.n13958 VSS.n13943 0.00249311
R12144 VSS.n1770 VSS.n1769 0.00249311
R12145 VSS.n14019 VSS.n14018 0.00249311
R12146 VSS.n1725 VSS.n1717 0.00249311
R12147 VSS.n1732 VSS.n1724 0.00249311
R12148 VSS.n1729 VSS.n1726 0.00249311
R12149 VSS.n13554 VSS.n13553 0.00249311
R12150 VSS.n13516 VSS.n13514 0.00249311
R12151 VSS.n13527 VSS.n13526 0.00249311
R12152 VSS.n13523 VSS.n13522 0.00249311
R12153 VSS.n13565 VSS.n13563 0.00249311
R12154 VSS.n13566 VSS.n13559 0.00249311
R12155 VSS.n13573 VSS.n13558 0.00249311
R12156 VSS.n13578 VSS.n13557 0.00249311
R12157 VSS.n13606 VSS.n13605 0.00249311
R12158 VSS.n13490 VSS.n13482 0.00249311
R12159 VSS.n13497 VSS.n13489 0.00249311
R12160 VSS.n13494 VSS.n13491 0.00249311
R12161 VSS.n13307 VSS.n13306 0.00249311
R12162 VSS.n13313 VSS.n13312 0.00249311
R12163 VSS.n13319 VSS.n13318 0.00249311
R12164 VSS.n13323 VSS.n13322 0.00249311
R12165 VSS.n13326 VSS.n13325 0.00249311
R12166 VSS.n13330 VSS.n13329 0.00249311
R12167 VSS.n13336 VSS.n13335 0.00249311
R12168 VSS.n13296 VSS.n13295 0.00249311
R12169 VSS.n13408 VSS.n13407 0.00249311
R12170 VSS.n13435 VSS.n13434 0.00249311
R12171 VSS.n13445 VSS.n13444 0.00249311
R12172 VSS.n13439 VSS.n13438 0.00249311
R12173 VSS.n9429 VSS.n9428 0.00239617
R12174 VSS.n1601 VSS.n1600 0.00239617
R12175 VSS.n299 VSS.n298 0.00238
R12176 VSS.n4465 VSS.n4464 0.00238
R12177 VSS.n4476 VSS.n4475 0.00238
R12178 VSS.n4495 VSS.n4493 0.00238
R12179 VSS.n4509 VSS.n4507 0.00238
R12180 VSS.n380 VSS.n379 0.00238
R12181 VSS.n35 VSS.n34 0.00238
R12182 VSS.n178 VSS.n177 0.00238
R12183 VSS.n340 VSS.n337 0.00238
R12184 VSS.n267 VSS.n264 0.00238
R12185 VSS.n155 VSS.n152 0.00238
R12186 VSS.n94 VSS.n91 0.00238
R12187 VSS.n8630 VSS.n8563 0.00225009
R12188 VSS.n8733 VSS.n8732 0.00225009
R12189 VSS.n9705 VSS.n9640 0.00225009
R12190 VSS.n9120 VSS.n9119 0.00225009
R12191 VSS.n10822 VSS.n10821 0.00225009
R12192 VSS.n9775 VSS.n9774 0.00225009
R12193 VSS.n14367 VSS.n14366 0.00225009
R12194 VSS.n1081 VSS.n1080 0.00225009
R12195 VSS.n1331 VSS.n1330 0.00225009
R12196 VSS.n773 VSS.n772 0.00225009
R12197 VSS.n13378 VSS.n13377 0.00225009
R12198 VSS.n13843 VSS.n13842 0.00225009
R12199 VSS.n14348 VSS 0.00213006
R12200 VSS.n13824 VSS 0.00213006
R12201 VSS.n13361 VSS 0.00213006
R12202 VSS.n1584 VSS 0.00213006
R12203 VSS VSS.n469 0.00213006
R12204 VSS.n13419 VSS.n13417 0.00206853
R12205 VSS.n5607 VSS.n5605 0.0020625
R12206 VSS.n1062 VSS 0.00206214
R12207 VSS.n11511 VSS.n11510 0.00201061
R12208 VSS.n3285 VSS.n3284 0.00200697
R12209 VSS.n3278 VSS.n3276 0.00200697
R12210 VSS.n12818 VSS.n12817 0.00200683
R12211 VSS.n11295 VSS.n11294 0.002
R12212 VSS.n1312 VSS 0.00199422
R12213 VSS.n8629 VSS.n8628 0.00192045
R12214 VSS.n8708 VSS.n8320 0.00192045
R12215 VSS.n9704 VSS.n9703 0.00192045
R12216 VSS.n9115 VSS.n9053 0.00192045
R12217 VSS.n4025 VSS.n3955 0.00192045
R12218 VSS.n7478 VSS.n7420 0.00192045
R12219 VSS.n9428 VSS.n9427 0.00192045
R12220 VSS.n14364 VSS.n14363 0.00192045
R12221 VSS.n1078 VSS.n1077 0.00192045
R12222 VSS.n1328 VSS.n1327 0.00192045
R12223 VSS.n768 VSS.n687 0.00192045
R12224 VSS.n13375 VSS.n13374 0.00192045
R12225 VSS.n13840 VSS.n13839 0.00192045
R12226 VSS.n1600 VSS.n1599 0.00192045
R12227 VSS.n11475 VSS.n11472 0.00178939
R12228 VSS.n11220 VSS.n11211 0.00178939
R12229 VSS.n11208 VSS.n11205 0.00178939
R12230 VSS.n11268 VSS.n11265 0.00178939
R12231 VSS.n11273 VSS.n11270 0.00178939
R12232 VSS.n11419 VSS.n11418 0.00178939
R12233 VSS.n6242 VSS.n6241 0.00175017
R12234 VSS.n8843 VSS.n8840 0.00175017
R12235 VSS.n9542 VSS.n7594 0.00175017
R12236 VSS.n9861 VSS.n9856 0.00175017
R12237 VSS.n7604 VSS.n7600 0.00175017
R12238 VSS.n9532 VSS.n9530 0.00175017
R12239 VSS.n9908 VSS.n6268 0.00175017
R12240 VSS.n9927 VSS.n6251 0.00175017
R12241 VSS.n6249 VSS.n6244 0.00175017
R12242 VSS.n10038 VSS.n10033 0.00175017
R12243 VSS.n4641 VSS.n4638 0.00175017
R12244 VSS.n10021 VSS.n4643 0.00175017
R12245 VSS.n10012 VSS.n4647 0.00175017
R12246 VSS.n10003 VSS.n4651 0.00175017
R12247 VSS.n9994 VSS.n4655 0.00175017
R12248 VSS.n4441 VSS.n4154 0.00175017
R12249 VSS.n4354 VSS.n4207 0.00175017
R12250 VSS.n13145 VSS.n1903 0.00175017
R12251 VSS.n14148 VSS.n613 0.00175017
R12252 VSS.n14139 VSS.n615 0.00175017
R12253 VSS.n14041 VSS.n1705 0.00175017
R12254 VSS.n14047 VSS.n623 0.00175017
R12255 VSS.n14131 VSS.n14129 0.00175017
R12256 VSS.n12705 VSS.n12700 0.00175017
R12257 VSS.n1893 VSS.n1890 0.00175017
R12258 VSS.n13163 VSS.n1895 0.00175017
R12259 VSS.n13154 VSS.n1899 0.00175017
R12260 VSS.n12842 VSS.n2920 0.00175017
R12261 VSS.n12847 VSS.n2915 0.00175017
R12262 VSS.n2910 VSS.n2738 0.00175017
R12263 VSS.n12924 VSS.n2735 0.00175017
R12264 VSS.n2730 VSS.n2557 0.00175017
R12265 VSS.n12425 VSS.n2555 0.00175017
R12266 VSS.n3625 VSS.n3624 0.00173379
R12267 VSS.n3624 VSS.n3623 0.00173379
R12268 VSS.n11506 VSS.n11505 0.00152605
R12269 VSS.n11512 VSS.n11506 0.00151551
R12270 VSS.n13581 VSS.n13580 0.00151492
R12271 VSS.n13966 VSS.n13965 0.00151492
R12272 VSS.n12758 VSS.n12757 0.00151492
R12273 VSS.n2634 VSS.n2633 0.00151492
R12274 VSS.n2027 VSS.n1978 0.00151492
R12275 VSS.n4018 VSS.n4015 0.00151492
R12276 VSS.n7339 VSS.n7338 0.00151492
R12277 VSS.n10986 VSS.n3877 0.00151492
R12278 VSS.n6393 VSS.n6392 0.00151492
R12279 VSS.n6838 VSS.n6837 0.00151492
R12280 VSS.n9666 VSS.n9663 0.00151492
R12281 VSS.n8678 VSS.n8675 0.00151492
R12282 VSS.n8868 VSS.n8002 0.00151492
R12283 VSS.n9975 VSS.n9974 0.00151492
R12284 VSS.n9558 VSS.n7558 0.00151492
R12285 VSS.n8556 VSS.n8553 0.00151492
R12286 VSS.n7396 VSS.n7395 0.00151492
R12287 VSS.n3929 VSS.n3928 0.00151492
R12288 VSS.n9318 VSS.n9316 0.00151492
R12289 VSS.n7187 VSS.n7185 0.00151492
R12290 VSS.n7374 VSS.n7373 0.00151492
R12291 VSS.n9244 VSS.n9183 0.00151492
R12292 VSS.n8951 VSS.n7828 0.00151492
R12293 VSS.n7643 VSS.n7641 0.00151492
R12294 VSS.n7702 VSS.n7700 0.00151492
R12295 VSS.n9890 VSS.n9889 0.00151492
R12296 VSS.n8927 VSS.n7892 0.00151492
R12297 VSS.n6905 VSS.n6627 0.00151492
R12298 VSS.n6978 VSS.n6579 0.00151492
R12299 VSS.n6999 VSS.n6530 0.00151492
R12300 VSS.n7060 VSS.n7059 0.00151492
R12301 VSS.n6452 VSS.n6451 0.00151492
R12302 VSS.n5887 VSS.n5886 0.00151492
R12303 VSS.n5706 VSS.n5705 0.00151492
R12304 VSS.n5526 VSS.n5525 0.00151492
R12305 VSS.n5346 VSS.n5345 0.00151492
R12306 VSS.n10080 VSS.n10079 0.00151492
R12307 VSS.n4607 VSS.n4606 0.00151492
R12308 VSS.n10775 VSS.n4128 0.00151492
R12309 VSS.n4403 VSS.n4197 0.00151492
R12310 VSS.n4301 VSS.n4300 0.00151492
R12311 VSS.n1341 VSS.n1338 0.00151492
R12312 VSS.n14227 VSS.n579 0.00151492
R12313 VSS.n13131 VSS.n13130 0.00151492
R12314 VSS.n13052 VSS.n13051 0.00151492
R12315 VSS.n1393 VSS.n880 0.00151492
R12316 VSS.n1612 VSS.n1609 0.00151492
R12317 VSS.n1464 VSS.n1462 0.00151492
R12318 VSS.n13697 VSS.n13696 0.00151492
R12319 VSS.n13901 VSS.n13900 0.00151492
R12320 VSS.n1414 VSS.n836 0.00151492
R12321 VSS.n2214 VSS.n2212 0.00151492
R12322 VSS.n2130 VSS.n2128 0.00151492
R12323 VSS.n13195 VSS.n13194 0.00151492
R12324 VSS.n13923 VSS.n1814 0.00151492
R12325 VSS.n2664 VSS.n2662 0.00151492
R12326 VSS.n2814 VSS.n2813 0.00151492
R12327 VSS.n2845 VSS.n2843 0.00151492
R12328 VSS.n12638 VSS.n12637 0.00151492
R12329 VSS.n12718 VSS.n3019 0.00151492
R12330 VSS.n12248 VSS.n12247 0.00151492
R12331 VSS.n12141 VSS.n12140 0.00151492
R12332 VSS.n11973 VSS.n11972 0.00151492
R12333 VSS.n3545 VSS.n3544 0.00151492
R12334 VSS.n12597 VSS.n12596 0.00151492
R12335 VSS.n3141 VSS.n3140 0.00151492
R12336 VSS.n2633 VSS.n2607 0.00150769
R12337 VSS.n1979 VSS.n1978 0.00150769
R12338 VSS.n1414 VSS.n837 0.00150769
R12339 VSS.n6839 VSS.n6838 0.00150769
R12340 VSS.n8928 VSS.n8927 0.00150769
R12341 VSS.n9244 VSS.n9184 0.00150769
R12342 VSS.n9443 VSS.n9442 0.00150769
R12343 VSS.n8821 VSS.n8177 0.00150769
R12344 VSS.n8783 VSS.n8209 0.00150769
R12345 VSS.n8746 VSS.n8745 0.00150769
R12346 VSS.n9976 VSS.n9975 0.00150769
R12347 VSS.n8149 VSS.n8035 0.00150769
R12348 VSS.n8067 VSS.n8002 0.00150769
R12349 VSS.n9558 VSS.n7556 0.00150769
R12350 VSS.n9316 VSS.n9315 0.00150769
R12351 VSS.n7220 VSS.n7185 0.00150769
R12352 VSS.n7373 VSS.n7209 0.00150769
R12353 VSS.n8951 VSS.n7819 0.00150769
R12354 VSS.n7733 VSS.n7641 0.00150769
R12355 VSS.n7700 VSS.n7699 0.00150769
R12356 VSS.n9891 VSS.n9890 0.00150769
R12357 VSS.n6906 VSS.n6905 0.00150769
R12358 VSS.n6979 VSS.n6978 0.00150769
R12359 VSS.n6999 VSS.n6521 0.00150769
R12360 VSS.n7059 VSS.n6290 0.00150769
R12361 VSS.n6453 VSS.n6452 0.00150769
R12362 VSS.n3721 VSS.n3718 0.00150769
R12363 VSS.n6393 VSS.n6391 0.00150769
R12364 VSS.n3877 VSS.n3858 0.00150769
R12365 VSS.n7339 VSS.n7337 0.00150769
R12366 VSS.n4302 VSS.n4301 0.00150769
R12367 VSS.n4197 VSS.n4188 0.00150769
R12368 VSS.n4128 VSS.n4113 0.00150769
R12369 VSS.n1269 VSS.n1268 0.00150769
R12370 VSS.n14199 VSS.n603 0.00150769
R12371 VSS.n960 VSS.n957 0.00150769
R12372 VSS.n13051 VSS.n2479 0.00150769
R12373 VSS.n2456 VSS.n2454 0.00150769
R12374 VSS.n13132 VSS.n13131 0.00150769
R12375 VSS.n579 VSS.n570 0.00150769
R12376 VSS.n1394 VSS.n1393 0.00150769
R12377 VSS.n13716 VSS.n13715 0.00150769
R12378 VSS.n13256 VSS.n13255 0.00150769
R12379 VSS.n1685 VSS.n1462 0.00150769
R12380 VSS.n13696 VSS.n13670 0.00150769
R12381 VSS.n13902 VSS.n13901 0.00150769
R12382 VSS.n2212 VSS.n2211 0.00150769
R12383 VSS.n2128 VSS.n2127 0.00150769
R12384 VSS.n13194 VSS.n1850 0.00150769
R12385 VSS.n12686 VSS.n1814 0.00150769
R12386 VSS.n2716 VSS.n2662 0.00150769
R12387 VSS.n2813 VSS.n2787 0.00150769
R12388 VSS.n2896 VSS.n2843 0.00150769
R12389 VSS.n12637 VSS.n3054 0.00150769
R12390 VSS.n3077 VSS.n3019 0.00150769
R12391 VSS.n12758 VSS.n2945 0.00150769
R12392 VSS.n13967 VSS.n13966 0.00150769
R12393 VSS.n13581 VSS.n13556 0.00150769
R12394 VSS.n13301 VSS.n13298 0.00150769
R12395 VSS.n11329 VSS.n11328 0.00150431
R12396 VSS.n11340 VSS.n11336 0.00150431
R12397 VSS.n11305 VSS.n11304 0.0015
R12398 VSS.n11324 VSS.n11314 0.0015
R12399 VSS.n3282 VSS.n3280 0.00149516
R12400 VSS.n3282 VSS.n3215 0.00149516
R12401 VSS.n12819 VSS.n12804 0.00149516
R12402 VSS.n11490 VSS.n11489 0.00146193
R12403 VSS.n10791 VSS.n10790 0.00125069
R12404 VSS.n10736 VSS.n10735 0.00125069
R12405 VSS.n4331 VSS.n4330 0.0012504
R12406 VSS.n11200 VSS.n11199 0.00118497
R12407 VSS.n11199 VSS.n11198 0.00118497
R12408 VSS.n14462 VSS.n14461 0.00115542
R12409 VSS.n3303 VSS.n3297 0.00114286
R12410 VSS.n3339 VSS.n3335 0.00114286
R12411 VSS.n3393 VSS.n3389 0.00114286
R12412 VSS.n11822 VSS.n11818 0.00114286
R12413 VSS.n11805 VSS.n11801 0.00114286
R12414 VSS.n12278 VSS.n12272 0.00114286
R12415 VSS.n12357 VSS.n12355 0.00114286
R12416 VSS.n1511 VSS.n1509 0.00114286
R12417 VSS.n7489 VSS.n7485 0.00114286
R12418 VSS.n990 VSS.n988 0.00114286
R12419 VSS.n12332 VSS.n12331 0.00114286
R12420 VSS.n1320 VSS.n1319 0.00114286
R12421 VSS.n11924 VSS.n11923 0.00114286
R12422 VSS.n12037 VSS.n12032 0.00114286
R12423 VSS.n11758 VSS.n11757 0.00114286
R12424 VSS.n5601 VSS.n5600 0.00114281
R12425 VSS.n5421 VSS.n5420 0.00114281
R12426 VSS.n5241 VSS.n5240 0.00114281
R12427 VSS.n10104 VSS.n4569 0.00114281
R12428 VSS.n11147 VSS.n3711 0.00114281
R12429 VSS.n11522 VSS.n11518 0.00114266
R12430 VSS.n10724 VSS.n505 0.00114214
R12431 VSS.n10803 VSS.n10802 0.00114214
R12432 VSS.n13747 VSS.n13743 0.00114214
R12433 VSS.n13284 VSS.n13280 0.00114214
R12434 VSS.n13414 VSS.n13410 0.00114214
R12435 VSS.n5959 VSS.n5957 0.00114214
R12436 VSS.n5778 VSS.n5776 0.00114214
R12437 VSS.n6142 VSS.n6140 0.00114214
R12438 VSS.n19 VSS.n15 0.001142
R12439 VSS.n14479 VSS.n14475 0.001142
R12440 VSS.n4097 VSS.n4094 0.00106587
R12441 VSS.n14353 VSS.n14352 0.00106587
R12442 VSS.n1067 VSS.n1064 0.00106587
R12443 VSS.n1589 VSS.n1586 0.00106587
R12444 VSS.n13829 VSS.n13826 0.00106587
R12445 VSS.n461 VSS.n460 0.00106587
R12446 VSS.n696 VSS.n695 0.00106587
R12447 VSS.n3438 VSS.n3435 0.00106587
R12448 VSS.n11920 VSS.n11919 0.00106587
R12449 VSS.n12036 VSS.n12033 0.00106587
R12450 VSS.n10734 VSS.n10649 0.00106586
R12451 VSS.n1591 VSS.n1590 0.00106586
R12452 VSS.n13831 VSS.n13830 0.00106586
R12453 VSS.n11532 VSS.n11531 0.00106582
R12454 VSS.n10719 VSS.n10718 0.00106068
R12455 VSS.n8426 VSS.n8425 0.00106068
R12456 VSS.n11531 VSS.n11530 0.00106068
R12457 VSS.n10649 VSS.n10648 0.00106064
R12458 VSS.n1592 VSS.n1591 0.00106064
R12459 VSS.n13832 VSS.n13831 0.00106064
R12460 VSS.n14354 VSS.n14353 0.00106063
R12461 VSS.n1064 VSS.n1063 0.00106063
R12462 VSS.n1586 VSS.n1585 0.00106063
R12463 VSS.n13826 VSS.n13825 0.00106063
R12464 VSS.n468 VSS.n461 0.00106063
R12465 VSS.n697 VSS.n696 0.00106063
R12466 VSS.n1314 VSS.n1313 0.00106063
R12467 VSS.n11774 VSS.n11773 0.00106063
R12468 VSS.n11921 VSS.n11920 0.00106063
R12469 VSS.n3435 VSS.n3434 0.00106063
R12470 VSS.n11288 VSS.n11278 0.00105948
R12471 VSS.n11530 VSS.n11529 0.00104326
R12472 VSS.n8426 VSS.n8424 0.00104326
R12473 VSS.n10723 VSS.n10719 0.00104326
R12474 VSS.n4098 VSS.n4093 0.00104326
R12475 VSS.n6146 VSS.n6145 0.00104325
R12476 VSS.n5963 VSS.n5962 0.00104325
R12477 VSS.n5782 VSS.n5781 0.00104325
R12478 VSS.n10142 VSS.n10138 0.00104325
R12479 VSS.n5194 VSS.n5190 0.00104325
R12480 VSS.n5374 VSS.n5370 0.00104325
R12481 VSS.n5554 VSS.n5550 0.00104325
R12482 VSS.n5734 VSS.n5730 0.00104325
R12483 VSS.n5915 VSS.n5911 0.00104325
R12484 VSS.n6097 VSS.n6093 0.00104325
R12485 VSS.n11076 VSS.n3703 0.00104325
R12486 VSS.n14478 VSS.n14477 0.0010432
R12487 VSS.n14355 VSS.n14339 0.00104317
R12488 VSS.n702 VSS.n698 0.00104317
R12489 VSS.n1315 VSS.n1303 0.00104317
R12490 VSS.n12202 VSS.n11775 0.00104317
R12491 VSS.n12038 VSS.n11808 0.00104317
R12492 VSS.n11524 VSS.n11523 0.00104317
R12493 VSS.n11149 VSS.n11148 0.00104317
R12494 VSS.n5597 VSS.n5596 0.00104317
R12495 VSS.n5417 VSS.n5416 0.00104317
R12496 VSS.n5237 VSS.n5236 0.00104317
R12497 VSS.n10106 VSS.n10105 0.00104317
R12498 VSS.n11460 VSS.n11457 0.00103939
R12499 VSS.n11465 VSS.n11462 0.00103939
R12500 VSS.n11470 VSS.n11467 0.00103939
R12501 VSS.n11470 VSS.n11469 0.00103939
R12502 VSS.n11465 VSS.n11464 0.00103939
R12503 VSS.n11460 VSS.n11459 0.00103939
R12504 VSS.n11475 VSS.n11474 0.00103939
R12505 VSS.n11211 VSS.n11210 0.00103939
R12506 VSS.n11208 VSS.n11207 0.00103939
R12507 VSS.n11268 VSS.n11267 0.00103939
R12508 VSS.n11273 VSS.n11272 0.00103939
R12509 VSS.n11418 VSS.n11417 0.00103939
R12510 VSS.n11476 VSS.n11475 0.00103403
R12511 VSS.n11261 VSS.n11211 0.00103403
R12512 VSS.n11261 VSS.n11208 0.00103403
R12513 VSS.n11274 VSS.n11268 0.00103403
R12514 VSS.n11274 VSS.n11273 0.00103403
R12515 VSS.n11418 VSS.n11415 0.00103403
R12516 VSS.n7505 VSS.n7496 0.00103325
R12517 VSS.n7512 VSS.n7508 0.00103325
R12518 VSS.n8328 VSS.n8324 0.00103325
R12519 VSS.n8335 VSS.n8331 0.00103325
R12520 VSS.n3963 VSS.n3959 0.00103325
R12521 VSS.n7493 VSS.n7492 0.00103325
R12522 VSS.n4031 VSS.n3967 0.00103325
R12523 VSS.n9766 VSS.n7479 0.00103325
R12524 VSS.n7491 VSS.n7490 0.00103325
R12525 VSS.n7495 VSS.n7494 0.00103325
R12526 VSS.n7507 VSS.n7506 0.00103325
R12527 VSS.n8714 VSS.n8650 0.00103325
R12528 VSS.n8330 VSS.n8329 0.00103325
R12529 VSS.n13366 VSS.n13352 0.00103325
R12530 VSS.n13367 VSS.n13366 0.00103325
R12531 VSS.n4098 VSS.n4097 0.00103324
R12532 VSS.n10723 VSS.n10722 0.00103324
R12533 VSS.n8424 VSS.n8423 0.00103324
R12534 VSS.n11529 VSS.n11528 0.00103324
R12535 VSS.n10142 VSS.n10141 0.00103323
R12536 VSS.n5194 VSS.n5193 0.00103323
R12537 VSS.n5374 VSS.n5373 0.00103323
R12538 VSS.n5554 VSS.n5553 0.00103323
R12539 VSS.n5734 VSS.n5733 0.00103323
R12540 VSS.n5915 VSS.n5914 0.00103323
R12541 VSS.n6097 VSS.n6096 0.00103323
R12542 VSS.n3703 VSS.n3702 0.00103323
R12543 VSS.n507 VSS.n506 0.00103323
R12544 VSS.n1236 VSS.n1235 0.00103323
R12545 VSS.n13286 VSS.n13285 0.00103323
R12546 VSS.n13416 VSS.n13415 0.00103323
R12547 VSS.n5964 VSS.n5963 0.00103323
R12548 VSS.n5783 VSS.n5782 0.00103323
R12549 VSS.n6147 VSS.n6146 0.00103323
R12550 VSS.n14470 VSS.n14469 0.00103322
R12551 VSS.n14477 VSS.n14476 0.00103319
R12552 VSS.n14 VSS.n13 0.00103319
R12553 VSS.n8417 VSS.n8338 0.00103319
R12554 VSS.n8641 VSS.n8639 0.00103319
R12555 VSS.n8649 VSS.n8646 0.00103319
R12556 VSS.n8722 VSS.n8721 0.00103319
R12557 VSS.n8715 VSS.n7515 0.00103319
R12558 VSS.n9716 VSS.n9714 0.00103319
R12559 VSS.n9724 VSS.n9721 0.00103319
R12560 VSS.n9733 VSS.n9731 0.00103319
R12561 VSS.n9741 VSS.n9738 0.00103319
R12562 VSS.n9749 VSS.n9747 0.00103319
R12563 VSS.n9760 VSS.n9758 0.00103319
R12564 VSS.n9761 VSS.n3966 0.00103319
R12565 VSS.n10811 VSS.n10810 0.00103319
R12566 VSS.n10810 VSS.n10808 0.00103319
R12567 VSS.n10812 VSS.n3966 0.00103319
R12568 VSS.n9765 VSS.n9760 0.00103319
R12569 VSS.n9753 VSS.n9749 0.00103319
R12570 VSS.n9746 VSS.n9741 0.00103319
R12571 VSS.n9737 VSS.n9733 0.00103319
R12572 VSS.n9730 VSS.n9724 0.00103319
R12573 VSS.n9720 VSS.n9716 0.00103319
R12574 VSS.n9713 VSS.n7515 0.00103319
R12575 VSS.n8721 VSS.n8719 0.00103319
R12576 VSS.n8723 VSS.n8649 0.00103319
R12577 VSS.n8645 VSS.n8641 0.00103319
R12578 VSS.n8638 VSS.n8338 0.00103319
R12579 VSS.n13365 VSS.n13364 0.00103319
R12580 VSS.n13364 VSS.n13362 0.00103319
R12581 VSS.n12575 VSS.n3175 0.00103319
R12582 VSS.n12575 VSS.n12574 0.00103319
R12583 VSS.n14355 VSS.n14354 0.00103317
R12584 VSS.n468 VSS.n467 0.00103317
R12585 VSS.n1315 VSS.n1314 0.00103317
R12586 VSS.n698 VSS.n697 0.00103317
R12587 VSS.n11775 VSS.n11774 0.00103317
R12588 VSS.n11808 VSS.n11807 0.00103317
R12589 VSS.n11922 VSS.n11921 0.00103317
R12590 VSS.n3434 VSS.n3433 0.00103317
R12591 VSS.n14352 VSS.n14349 0.0010331
R12592 VSS.n7489 VSS.n7488 0.0010331
R12593 VSS.n988 VSS.n987 0.0010331
R12594 VSS.n1319 VSS.n1318 0.0010331
R12595 VSS.n460 VSS.n457 0.0010331
R12596 VSS.n11757 VSS.n11756 0.0010331
R12597 VSS.n12037 VSS.n12036 0.0010331
R12598 VSS.n3439 VSS.n3438 0.0010331
R12599 VSS.n1509 VSS.n1508 0.0010331
R12600 VSS.n3297 VSS.n3296 0.0010331
R12601 VSS.n3339 VSS.n3338 0.0010331
R12602 VSS.n3393 VSS.n3392 0.0010331
R12603 VSS.n11822 VSS.n11821 0.0010331
R12604 VSS.n11805 VSS.n11804 0.0010331
R12605 VSS.n12272 VSS.n12271 0.0010331
R12606 VSS.n12331 VSS.n12330 0.0010331
R12607 VSS.n12355 VSS.n12354 0.0010331
R12608 VSS.n5602 VSS.n5601 0.00103308
R12609 VSS.n5422 VSS.n5421 0.00103308
R12610 VSS.n5242 VSS.n5241 0.00103308
R12611 VSS.n10104 VSS.n10103 0.00103308
R12612 VSS.n11147 VSS.n11146 0.00103308
R12613 VSS.n11522 VSS.n11521 0.00103305
R12614 VSS.n10804 VSS.n10803 0.00103293
R12615 VSS.n14374 VSS.n505 0.00103293
R12616 VSS.n1239 VSS.n1234 0.00103293
R12617 VSS.n13751 VSS.n13747 0.00103293
R12618 VSS.n13289 VSS.n13284 0.00103293
R12619 VSS.n13421 VSS.n13414 0.00103293
R12620 VSS.n6140 VSS.n6139 0.00103293
R12621 VSS.n5957 VSS.n4668 0.00103293
R12622 VSS.n5776 VSS.n4677 0.00103293
R12623 VSS.n14480 VSS.n14479 0.0010329
R12624 VSS.n19 VSS.n18 0.0010329
R12625 VSS.n11329 VSS.n3699 0.00102396
R12626 VSS.n11336 VSS.n3697 0.00102396
R12627 VSS.n10150 VSS.n10149 0.00102352
R12628 VSS.n5202 VSS.n5201 0.00102352
R12629 VSS.n5382 VSS.n5381 0.00102352
R12630 VSS.n5562 VSS.n5561 0.00102352
R12631 VSS.n5742 VSS.n5741 0.00102352
R12632 VSS.n5923 VSS.n5922 0.00102352
R12633 VSS.n6105 VSS.n6104 0.00102352
R12634 VSS.n11191 VSS.n11183 0.00102352
R12635 VSS.n10727 VSS.n10726 0.00102352
R12636 VSS.n9756 VSS.n9755 0.00102352
R12637 VSS.n8419 VSS.n8418 0.00102352
R12638 VSS.n983 VSS.n982 0.00102352
R12639 VSS.n1504 VSS.n1503 0.00102352
R12640 VSS.n3306 VSS.n3305 0.00102352
R12641 VSS.n3361 VSS.n3360 0.00102352
R12642 VSS.n3568 VSS.n3567 0.00102352
R12643 VSS.n11997 VSS.n11996 0.00102352
R12644 VSS.n12164 VSS.n12163 0.00102352
R12645 VSS.n11688 VSS.n11687 0.00102352
R12646 VSS.n12336 VSS.n12335 0.00102352
R12647 VSS.n12350 VSS.n11567 0.00102352
R12648 VSS.n12466 VSS.n11533 0.00102352
R12649 VSS.n10733 VSS.n10732 0.00102351
R12650 VSS.n1069 VSS.n1068 0.0010235
R12651 VSS.n3307 VSS.n3304 0.0010235
R12652 VSS.n12165 VSS.n11776 0.0010235
R12653 VSS.n12280 VSS.n12279 0.0010235
R12654 VSS.n12334 VSS.n12333 0.0010235
R12655 VSS.n14503 VSS.n14502 0.0010235
R12656 VSS.n14472 VSS.n14471 0.0010235
R12657 VSS.n14473 VSS.n14463 0.00102105
R12658 VSS.n14500 VSS.n14497 0.00102105
R12659 VSS.n14496 VSS.n14495 0.00102105
R12660 VSS.n14506 VSS.n12 0.00102105
R12661 VSS.n3209 VSS.n3208 0.00102105
R12662 VSS.n3210 VSS.n3209 0.00102057
R12663 VSS.n14472 VSS.n14468 0.00102057
R12664 VSS.n14503 VSS.n14496 0.00102057
R12665 VSS.n6093 VSS.n4669 0.00101835
R12666 VSS.n5911 VSS.n4678 0.00101835
R12667 VSS.n5730 VSS.n4687 0.00101835
R12668 VSS.n5550 VSS.n4698 0.00101835
R12669 VSS.n5370 VSS.n4710 0.00101835
R12670 VSS.n5190 VSS.n5184 0.00101835
R12671 VSS.n10138 VSS.n10131 0.00101835
R12672 VSS.n11076 VSS.n11075 0.00101835
R12673 VSS.n14502 VSS.n14501 0.00101832
R12674 VSS.n14471 VSS.n14470 0.00101832
R12675 VSS.n7485 VSS.n7480 0.00101832
R12676 VSS.n990 VSS.n989 0.00101832
R12677 VSS.n1511 VSS.n1510 0.00101832
R12678 VSS.n3304 VSS.n3303 0.00101832
R12679 VSS.n3335 VSS.n3329 0.00101832
R12680 VSS.n3389 VSS.n3383 0.00101832
R12681 VSS.n11818 VSS.n11812 0.00101832
R12682 VSS.n11801 VSS.n11776 0.00101832
R12683 VSS.n12279 VSS.n12278 0.00101832
R12684 VSS.n12357 VSS.n12356 0.00101832
R12685 VSS.n12333 VSS.n12332 0.00101832
R12686 VSS.n1070 VSS.n1069 0.00101831
R12687 VSS.n10734 VSS.n10733 0.0010183
R12688 VSS.n10728 VSS.n10727 0.0010183
R12689 VSS.n9755 VSS.n9754 0.0010183
R12690 VSS.n982 VSS.n981 0.0010183
R12691 VSS.n1503 VSS.n1502 0.0010183
R12692 VSS.n3307 VSS.n3306 0.0010183
R12693 VSS.n3362 VSS.n3361 0.0010183
R12694 VSS.n3569 VSS.n3568 0.0010183
R12695 VSS.n11998 VSS.n11997 0.0010183
R12696 VSS.n12165 VSS.n12164 0.0010183
R12697 VSS.n11567 VSS.n11566 0.0010183
R12698 VSS.n12335 VSS.n12334 0.0010183
R12699 VSS.n11533 VSS.n11532 0.0010183
R12700 VSS.n6106 VSS.n6105 0.0010183
R12701 VSS.n5924 VSS.n5923 0.0010183
R12702 VSS.n5743 VSS.n5742 0.0010183
R12703 VSS.n5563 VSS.n5562 0.0010183
R12704 VSS.n5383 VSS.n5382 0.0010183
R12705 VSS.n5203 VSS.n5202 0.0010183
R12706 VSS.n10151 VSS.n10150 0.0010183
R12707 VSS.n11183 VSS.n11182 0.0010183
R12708 VSS.n11289 VSS.n11288 0.00101822
R12709 VSS.n13328 VSS.n13327 0.00101585
R12710 VSS.n13440 VSS.n13437 0.00101585
R12711 VSS.n13564 VSS.n13562 0.00101585
R12712 VSS.n13492 VSS.n13487 0.00101585
R12713 VSS.n13948 VSS.n13946 0.00101585
R12714 VSS.n1727 VSS.n1722 0.00101585
R12715 VSS.n12740 VSS.n12739 0.00101585
R12716 VSS.n12765 VSS.n2938 0.00101585
R12717 VSS.n2597 VSS.n2596 0.00101585
R12718 VSS.n2017 VSS.n2016 0.00101585
R12719 VSS.n4001 VSS.n4000 0.00101585
R12720 VSS.n4043 VSS.n4040 0.00101585
R12721 VSS.n7284 VSS.n7283 0.00101585
R12722 VSS.n10860 VSS.n3901 0.00101585
R12723 VSS.n10971 VSS.n3873 0.00101585
R12724 VSS.n10906 VSS.n10905 0.00101585
R12725 VSS.n6338 VSS.n6337 0.00101585
R12726 VSS.n11011 VSS.n3833 0.00101585
R12727 VSS.n3741 VSS.n3740 0.00101585
R12728 VSS.n6820 VSS.n6818 0.00101585
R12729 VSS.n9682 VSS.n9681 0.00101585
R12730 VSS.n9052 VSS.n9049 0.00101585
R12731 VSS.n8351 VSS.n8348 0.00101585
R12732 VSS.n8449 VSS.n8446 0.00101585
R12733 VSS.n8694 VSS.n8693 0.00101585
R12734 VSS.n9624 VSS.n9621 0.00101585
R12735 VSS.n8305 VSS.n8302 0.00101585
R12736 VSS.n8250 VSS.n8249 0.00101585
R12737 VSS.n6193 VSS.n6190 0.00101585
R12738 VSS.n9957 VSS.n9955 0.00101585
R12739 VSS.n8854 VSS.n8853 0.00101585
R12740 VSS.n9339 VSS.n9336 0.00101585
R12741 VSS.n9815 VSS.n9813 0.00101585
R12742 VSS.n7201 VSS.n7194 0.00101585
R12743 VSS.n7353 VSS.n7272 0.00101585
R12744 VSS.n9173 VSS.n9169 0.00101585
R12745 VSS.n7832 VSS.n7815 0.00101585
R12746 VSS.n7788 VSS.n7786 0.00101585
R12747 VSS.n7709 VSS.n7707 0.00101585
R12748 VSS.n9872 VSS.n9870 0.00101585
R12749 VSS.n7122 VSS.n7116 0.00101585
R12750 VSS.n7922 VSS.n7888 0.00101585
R12751 VSS.n7985 VSS.n7984 0.00101585
R12752 VSS.n6887 VSS.n6885 0.00101585
R12753 VSS.n6960 VSS.n6958 0.00101585
R12754 VSS.n7002 VSS.n6517 0.00101585
R12755 VSS.n6279 VSS.n6275 0.00101585
R12756 VSS.n6434 VSS.n6432 0.00101585
R12757 VSS.n6407 VSS.n6326 0.00101585
R12758 VSS.n6723 VSS.n6680 0.00101585
R12759 VSS.n5894 VSS.n5893 0.00101585
R12760 VSS.n5713 VSS.n5712 0.00101585
R12761 VSS.n5533 VSS.n5532 0.00101585
R12762 VSS.n5353 VSS.n5352 0.00101585
R12763 VSS.n10087 VSS.n10086 0.00101585
R12764 VSS.n4611 VSS.n4610 0.00101585
R12765 VSS.n3796 VSS.n3793 0.00101585
R12766 VSS.n5990 VSS.n5989 0.00101585
R12767 VSS.n11060 VSS.n11057 0.00101585
R12768 VSS.n4122 VSS.n4119 0.00101585
R12769 VSS.n10754 VSS.n10752 0.00101585
R12770 VSS.n4386 VSS.n4190 0.00101585
R12771 VSS.n4283 VSS.n4281 0.00101585
R12772 VSS.n4241 VSS.n4236 0.00101585
R12773 VSS.n1288 VSS.n1287 0.00101585
R12774 VSS.n686 VSS.n683 0.00101585
R12775 VSS.n1216 VSS.n1213 0.00101585
R12776 VSS.n964 VSS.n961 0.00101585
R12777 VSS.n14210 VSS.n572 0.00101585
R12778 VSS.n563 VSS.n556 0.00101585
R12779 VSS.n14265 VSS.n14262 0.00101585
R12780 VSS.n13031 VSS.n2492 0.00101585
R12781 VSS.n2471 VSS.n2465 0.00101585
R12782 VSS.n2366 VSS.n2364 0.00101585
R12783 VSS.n13113 VSS.n13111 0.00101585
R12784 VSS.n1485 VSS.n1482 0.00101585
R12785 VSS.n13658 VSS.n13657 0.00101585
R12786 VSS.n13883 VSS.n13881 0.00101585
R12787 VSS.n13629 VSS.n13233 0.00101585
R12788 VSS.n826 VSS.n822 0.00101585
R12789 VSS.n2222 VSS.n2220 0.00101585
R12790 VSS.n2157 VSS.n2155 0.00101585
R12791 VSS.n1839 VSS.n1835 0.00101585
R12792 VSS.n1823 VSS.n1821 0.00101585
R12793 VSS.n1787 VSS.n1785 0.00101585
R12794 VSS.n1960 VSS.n1954 0.00101585
R12795 VSS.n12962 VSS.n12960 0.00101585
R12796 VSS.n2778 VSS.n2777 0.00101585
R12797 VSS.n12885 VSS.n12883 0.00101585
R12798 VSS.n3042 VSS.n3041 0.00101585
R12799 VSS.n3028 VSS.n3026 0.00101585
R12800 VSS.n2965 VSS.n2963 0.00101585
R12801 VSS.n2512 VSS.n2506 0.00101585
R12802 VSS.n12255 VSS.n12254 0.00101585
R12803 VSS.n12148 VSS.n12147 0.00101585
R12804 VSS.n11980 VSS.n11979 0.00101585
R12805 VSS.n3552 VSS.n3551 0.00101585
R12806 VSS.n12604 VSS.n12603 0.00101585
R12807 VSS.n3145 VSS.n3144 0.00101585
R12808 VSS.n11605 VSS.n11604 0.00101585
R12809 VSS.n4541 VSS.n4536 0.00101562
R12810 VSS.n12323 VSS.n12321 0.00101562
R12811 VSS.n12180 VSS.n12178 0.00101562
R12812 VSS.n12198 VSS.n12196 0.00101562
R12813 VSS.n14494 VSS.n14492 0.00101562
R12814 VSS.n12567 VSS.n12565 0.00101562
R12815 VSS.n3414 VSS.n3412 0.00101562
R12816 VSS.n11899 VSS.n11897 0.00101562
R12817 VSS.n12012 VSS.n12010 0.00101562
R12818 VSS.n13460 VSS.n13457 0.001014
R12819 VSS.n13592 VSS.n13503 0.001014
R12820 VSS.n14005 VSS.n1738 0.001014
R12821 VSS.n12790 VSS.n12786 0.001014
R12822 VSS.n4070 VSS.n4067 0.001014
R12823 VSS.n10885 VSS.n10881 0.001014
R12824 VSS.n10930 VSS.n10929 0.001014
R12825 VSS.n11036 VSS.n11032 0.001014
R12826 VSS.n9034 VSS.n9031 0.001014
R12827 VSS.n9646 VSS.n9643 0.001014
R12828 VSS.n7580 VSS.n7579 0.001014
R12829 VSS.n8472 VSS.n8469 0.001014
R12830 VSS.n8801 VSS.n8800 0.001014
R12831 VSS.n7535 VSS.n7532 0.001014
R12832 VSS.n8658 VSS.n8655 0.001014
R12833 VSS.n8593 VSS.n8590 0.001014
R12834 VSS.n8289 VSS.n8286 0.001014
R12835 VSS.n8228 VSS.n8227 0.001014
R12836 VSS.n8203 VSS.n8199 0.001014
R12837 VSS.n6170 VSS.n6167 0.001014
R12838 VSS.n6229 VSS.n6219 0.001014
R12839 VSS.n6704 VSS.n6699 0.001014
R12840 VSS.n8077 VSS.n8043 0.001014
R12841 VSS.n8135 VSS.n8134 0.001014
R12842 VSS.n8057 VSS.n8056 0.001014
R12843 VSS.n7961 VSS.n7956 0.001014
R12844 VSS.n8171 VSS.n8167 0.001014
R12845 VSS.n9576 VSS.n7562 0.001014
R12846 VSS.n8551 VSS.n8548 0.001014
R12847 VSS.n9393 VSS.n9390 0.001014
R12848 VSS.n7412 VSS.n7409 0.001014
R12849 VSS.n7450 VSS.n7447 0.001014
R12850 VSS.n3948 VSS.n3945 0.001014
R12851 VSS.n9087 VSS.n9084 0.001014
R12852 VSS.n9323 VSS.n9320 0.001014
R12853 VSS.n9009 VSS.n9005 0.001014
R12854 VSS.n9299 VSS.n9297 0.001014
R12855 VSS.n7173 VSS.n7169 0.001014
R12856 VSS.n7245 VSS.n7243 0.001014
R12857 VSS.n7320 VSS.n7268 0.001014
R12858 VSS.n9224 VSS.n9223 0.001014
R12859 VSS.n9248 VSS.n9166 0.001014
R12860 VSS.n7863 VSS.n7862 0.001014
R12861 VSS.n8971 VSS.n7627 0.001014
R12862 VSS.n7761 VSS.n7662 0.001014
R12863 VSS.n7086 VSS.n7076 0.001014
R12864 VSS.n7101 VSS.n7095 0.001014
R12865 VSS.n8907 VSS.n8906 0.001014
R12866 VSS.n7882 VSS.n7878 0.001014
R12867 VSS.n6648 VSS.n6639 0.001014
R12868 VSS.n6617 VSS.n6613 0.001014
R12869 VSS.n6600 VSS.n6591 0.001014
R12870 VSS.n6569 VSS.n6565 0.001014
R12871 VSS.n6552 VSS.n6551 0.001014
R12872 VSS.n6502 VSS.n6493 0.001014
R12873 VSS.n6313 VSS.n6303 0.001014
R12874 VSS.n6374 VSS.n6322 0.001014
R12875 VSS.n6771 VSS.n6685 0.001014
R12876 VSS.n6665 VSS.n6661 0.001014
R12877 VSS.n6020 VSS.n6017 0.001014
R12878 VSS.n5870 VSS.n5867 0.001014
R12879 VSS.n5822 VSS.n5819 0.001014
R12880 VSS.n5689 VSS.n5686 0.001014
R12881 VSS.n5641 VSS.n5638 0.001014
R12882 VSS.n5509 VSS.n5506 0.001014
R12883 VSS.n5461 VSS.n5458 0.001014
R12884 VSS.n5329 VSS.n5326 0.001014
R12885 VSS.n5281 VSS.n5278 0.001014
R12886 VSS.n10063 VSS.n10060 0.001014
R12887 VSS.n4602 VSS.n4599 0.001014
R12888 VSS.n3769 VSS.n3766 0.001014
R12889 VSS.n11094 VSS.n11091 0.001014
R12890 VSS.n3737 VSS.n3734 0.001014
R12891 VSS.n6357 VSS.n6356 0.001014
R12892 VSS.n3872 VSS.n3864 0.001014
R12893 VSS.n7303 VSS.n7302 0.001014
R12894 VSS.n3997 VSS.n3994 0.001014
R12895 VSS.n4143 VSS.n4142 0.001014
R12896 VSS.n4365 VSS.n4184 0.001014
R12897 VSS.n4333 VSS.n4252 0.001014
R12898 VSS.n4313 VSS.n4312 0.001014
R12899 VSS.n4423 VSS.n4118 0.001014
R12900 VSS.n668 VSS.n665 0.001014
R12901 VSS.n1252 VSS.n1249 0.001014
R12902 VSS.n1025 VSS.n1022 0.001014
R12903 VSS.n1200 VSS.n1197 0.001014
R12904 VSS.n901 VSS.n892 0.001014
R12905 VSS.n14322 VSS.n14319 0.001014
R12906 VSS.n2408 VSS.n552 0.001014
R12907 VSS.n523 VSS.n520 0.001014
R12908 VSS.n10658 VSS.n10655 0.001014
R12909 VSS.n922 VSS.n917 0.001014
R12910 VSS.n14185 VSS.n14184 0.001014
R12911 VSS.n12375 VSS.n12372 0.001014
R12912 VSS.n12404 VSS.n12403 0.001014
R12913 VSS.n2539 VSS.n2488 0.001014
R12914 VSS.n2377 VSS.n2359 0.001014
R12915 VSS.n13079 VSS.n13078 0.001014
R12916 VSS.n1927 VSS.n1917 0.001014
R12917 VSS.n2283 VSS.n1936 0.001014
R12918 VSS.n878 VSS.n868 0.001014
R12919 VSS.n1102 VSS.n1099 0.001014
R12920 VSS.n1547 VSS.n1544 0.001014
R12921 VSS.n13735 VSS.n13732 0.001014
R12922 VSS.n13787 VSS.n13784 0.001014
R12923 VSS.n13272 VSS.n13269 0.001014
R12924 VSS.n740 VSS.n737 0.001014
R12925 VSS.n1469 VSS.n1466 0.001014
R12926 VSS.n643 VSS.n639 0.001014
R12927 VSS.n1678 VSS.n1677 0.001014
R12928 VSS.n14065 VSS.n1657 0.001014
R12929 VSS.n13220 VSS.n13210 0.001014
R12930 VSS.n13538 VSS.n13229 0.001014
R12931 VSS.n853 VSS.n852 0.001014
R12932 VSS.n1418 VSS.n819 0.001014
R12933 VSS.n1998 VSS.n1994 0.001014
R12934 VSS.n2073 VSS.n2069 0.001014
R12935 VSS.n1872 VSS.n1863 0.001014
R12936 VSS.n12676 VSS.n12675 0.001014
R12937 VSS.n1798 VSS.n1780 0.001014
R12938 VSS.n2302 VSS.n1968 0.001014
R12939 VSS.n2260 VSS.n2258 0.001014
R12940 VSS.n2577 VSS.n2573 0.001014
R12941 VSS.n2706 VSS.n2705 0.001014
R12942 VSS.n12935 VSS.n2684 0.001014
R12943 VSS.n2796 VSS.n2794 0.001014
R12944 VSS.n2758 VSS.n2754 0.001014
R12945 VSS.n2886 VSS.n2885 0.001014
R12946 VSS.n12858 VSS.n2864 0.001014
R12947 VSS.n3067 VSS.n3066 0.001014
R12948 VSS.n3003 VSS.n2958 0.001014
R12949 VSS.n13007 VSS.n2520 0.001014
R12950 VSS.n2615 VSS.n2613 0.001014
R12951 VSS.n11661 VSS.n11658 0.001014
R12952 VSS.n12231 VSS.n12228 0.001014
R12953 VSS.n11730 VSS.n11727 0.001014
R12954 VSS.n12124 VSS.n12121 0.001014
R12955 VSS.n12076 VSS.n12073 0.001014
R12956 VSS.n11956 VSS.n11953 0.001014
R12957 VSS.n11862 VSS.n11859 0.001014
R12958 VSS.n3528 VSS.n3525 0.001014
R12959 VSS.n3480 VSS.n3477 0.001014
R12960 VSS.n3103 VSS.n3100 0.001014
R12961 VSS.n3136 VSS.n3133 0.001014
R12962 VSS.n3231 VSS.n3228 0.001014
R12963 VSS.n2987 VSS.n2986 0.001014
R12964 VSS.n13978 VSS.n13977 0.001014
R12965 VSS.n13521 VSS.n13520 0.001014
R12966 VSS.n13324 VSS.n13321 0.001014
R12967 VSS.n11478 VSS.n11477 0.00101218
R12968 VSS.n9744 VSS.n9742 0.0010119
R12969 VSS.n14508 VSS.n8 0.00100934
R12970 VSS.n14508 VSS.n14507 0.00100934
R12971 VSS.n3196 VSS.n3194 0.00100934
R12972 VSS.n11512 VSS.n11511 0.00100876
R12973 VSS.n4708 VSS.n4707 0.00100763
R12974 VSS.n4667 VSS.n4666 0.00100763
R12975 VSS.n4674 VSS.n4673 0.00100763
R12976 VSS.n4676 VSS.n4675 0.00100763
R12977 VSS.n4683 VSS.n4682 0.00100763
R12978 VSS.n4685 VSS.n4684 0.00100763
R12979 VSS.n4694 VSS.n4693 0.00100763
R12980 VSS.n4696 VSS.n4695 0.00100763
R12981 VSS.n4705 VSS.n4704 0.00100763
R12982 VSS.n4717 VSS.n4716 0.00100763
R12983 VSS.n5182 VSS.n5181 0.00100763
R12984 VSS.n4565 VSS.n4564 0.00100763
R12985 VSS.n10129 VSS.n10128 0.00100763
R12986 VSS.n3707 VSS.n3706 0.00100763
R12987 VSS.n3705 VSS.n3704 0.00100763
R12988 VSS.n3372 VSS.n3371 0.00100763
R12989 VSS.n6135 VSS.n6134 0.00100763
R12990 VSS.n12295 VSS.n12294 0.00100763
R12991 VSS.n12323 VSS.n12322 0.00100763
R12992 VSS.n11559 VSS.n11558 0.00100763
R12993 VSS.n12180 VSS.n12179 0.00100763
R12994 VSS.n12198 VSS.n12197 0.00100763
R12995 VSS.n14494 VSS.n14493 0.00100763
R12996 VSS.n14484 VSS.n14483 0.00100763
R12997 VSS.n3317 VSS.n3316 0.00100763
R12998 VSS.n12567 VSS.n12566 0.00100763
R12999 VSS.n3414 VSS.n3413 0.00100763
R13000 VSS.n3584 VSS.n3583 0.00100763
R13001 VSS.n11899 VSS.n11898 0.00100763
R13002 VSS.n12012 VSS.n12011 0.00100763
R13003 VSS.n12028 VSS.n12027 0.00100763
R13004 VSS.n10626 VSS.n10622 0.00100763
R13005 VSS.n11501 VSS.n11500 0.00100757
R13006 VSS.n7504 VSS.n7502 0.00100756
R13007 VSS.n7511 VSS.n7509 0.00100756
R13008 VSS.n8327 VSS.n8325 0.00100756
R13009 VSS.n8334 VSS.n8332 0.00100756
R13010 VSS.n3962 VSS.n3960 0.00100756
R13011 VSS.n4542 VSS.n4541 0.00100756
R13012 VSS.n9025 VSS.n9021 0.00100746
R13013 VSS.n8822 VSS.n8821 0.00100746
R13014 VSS.n8784 VSS.n8783 0.00100746
R13015 VSS.n7526 VSS.n7522 0.00100746
R13016 VSS.n8570 VSS.n8569 0.00100746
R13017 VSS.n8779 VSS.n8778 0.00100746
R13018 VSS.n6743 VSS.n6697 0.00100746
R13019 VSS.n8150 VSS.n8149 0.00100746
R13020 VSS.n8039 VSS.n8038 0.00100746
R13021 VSS.n8875 VSS.n7954 0.00100746
R13022 VSS.n8189 VSS.n8188 0.00100746
R13023 VSS.n7570 VSS.n7569 0.00100746
R13024 VSS.n8463 VSS.n8462 0.00100746
R13025 VSS.n9370 VSS.n9369 0.00100746
R13026 VSS.n7427 VSS.n7426 0.00100746
R13027 VSS.n9064 VSS.n9063 0.00100746
R13028 VSS.n9017 VSS.n8999 0.00100746
R13029 VSS.n7181 VSS.n7163 0.00100746
R13030 VSS.n7264 VSS.n7263 0.00100746
R13031 VSS.n9214 VSS.n9213 0.00100746
R13032 VSS.n7853 VSS.n7852 0.00100746
R13033 VSS.n7638 VSS.n7616 0.00100746
R13034 VSS.n7673 VSS.n7651 0.00100746
R13035 VSS.n7091 VSS.n7090 0.00100746
R13036 VSS.n7943 VSS.n7942 0.00100746
R13037 VSS.n6631 VSS.n6630 0.00100746
R13038 VSS.n6583 VSS.n6582 0.00100746
R13039 VSS.n6542 VSS.n6541 0.00100746
R13040 VSS.n6485 VSS.n6484 0.00100746
R13041 VSS.n6318 VSS.n6317 0.00100746
R13042 VSS.n6678 VSS.n6677 0.00100746
R13043 VSS.n5997 VSS.n5996 0.00100746
R13044 VSS.n5799 VSS.n5798 0.00100746
R13045 VSS.n5618 VSS.n5617 0.00100746
R13046 VSS.n5438 VSS.n5437 0.00100746
R13047 VSS.n5258 VSS.n5257 0.00100746
R13048 VSS.n3760 VSS.n3759 0.00100746
R13049 VSS.n6184 VSS.n6183 0.00100746
R13050 VSS.n11074 VSS.n11073 0.00100746
R13051 VSS.n11027 VSS.n3836 0.00100746
R13052 VSS.n10946 VSS.n10945 0.00100746
R13053 VSS.n10876 VSS.n3904 0.00100746
R13054 VSS.n4057 VSS.n4056 0.00100746
R13055 VSS.n4267 VSS.n4249 0.00100746
R13056 VSS.n4378 VSS.n4181 0.00100746
R13057 VSS.n4452 VSS.n4451 0.00100746
R13058 VSS.n659 VSS.n657 0.00100746
R13059 VSS.n1002 VSS.n1001 0.00100746
R13060 VSS.n14200 VSS.n14199 0.00100746
R13061 VSS.n10695 VSS.n10694 0.00100746
R13062 VSS.n514 VSS.n510 0.00100746
R13063 VSS.n1133 VSS.n915 0.00100746
R13064 VSS.n2484 VSS.n2483 0.00100746
R13065 VSS.n2454 VSS.n2453 0.00100746
R13066 VSS.n13093 VSS.n2357 0.00100746
R13067 VSS.n1932 VSS.n1931 0.00100746
R13068 VSS.n2399 VSS.n555 0.00100746
R13069 VSS.n884 VSS.n883 0.00100746
R13070 VSS.n14306 VSS.n14305 0.00100746
R13071 VSS.n1524 VSS.n1523 0.00100746
R13072 VSS.n13764 VSS.n13763 0.00100746
R13073 VSS.n717 VSS.n716 0.00100746
R13074 VSS.n651 VSS.n633 0.00100746
R13075 VSS.n1668 VSS.n1646 0.00100746
R13076 VSS.n13225 VSS.n13224 0.00100746
R13077 VSS.n843 VSS.n842 0.00100746
R13078 VSS.n2006 VSS.n1988 0.00100746
R13079 VSS.n2081 VSS.n2063 0.00100746
R13080 VSS.n1855 VSS.n1854 0.00100746
R13081 VSS.n13927 VSS.n1778 0.00100746
R13082 VSS.n1975 VSS.n1953 0.00100746
R13083 VSS.n2585 VSS.n2567 0.00100746
R13084 VSS.n2695 VSS.n2673 0.00100746
R13085 VSS.n2766 VSS.n2748 0.00100746
R13086 VSS.n2875 VSS.n2853 0.00100746
R13087 VSS.n12722 VSS.n2956 0.00100746
R13088 VSS.n2527 VSS.n2505 0.00100746
R13089 VSS.n11700 VSS.n11699 0.00100746
R13090 VSS.n12053 VSS.n12052 0.00100746
R13091 VSS.n11832 VSS.n11831 0.00100746
R13092 VSS.n3457 VSS.n3456 0.00100746
R13093 VSS.n3222 VSS.n3221 0.00100746
R13094 VSS.n12389 VSS.n12388 0.00100746
R13095 VSS.n12781 VSS.n2941 0.00100746
R13096 VSS.n1764 VSS.n1735 0.00100746
R13097 VSS.n13583 VSS.n13500 0.00100746
R13098 VSS.n13454 VSS.n13453 0.00100746
R13099 VSS.n13343 VSS.n13342 0.001007
R13100 VSS.n13301 VSS.n13300 0.001007
R13101 VSS.n13580 VSS.n13579 0.001007
R13102 VSS.n13556 VSS.n13555 0.001007
R13103 VSS.n13965 VSS.n13964 0.001007
R13104 VSS.n13968 VSS.n13967 0.001007
R13105 VSS.n12757 VSS.n12756 0.001007
R13106 VSS.n2977 VSS.n2945 0.001007
R13107 VSS.n2635 VSS.n2634 0.001007
R13108 VSS.n2028 VSS.n2027 0.001007
R13109 VSS.n836 VSS.n835 0.001007
R13110 VSS.n1612 VSS.n1611 0.001007
R13111 VSS.n4018 VSS.n4017 0.001007
R13112 VSS.n3974 VSS.n3973 0.001007
R13113 VSS.n7338 VSS.n7292 0.001007
R13114 VSS.n7337 VSS.n7336 0.001007
R13115 VSS.n10986 VSS.n10985 0.001007
R13116 VSS.n3860 VSS.n3858 0.001007
R13117 VSS.n6392 VSS.n6346 0.001007
R13118 VSS.n6391 VSS.n6390 0.001007
R13119 VSS.n11133 VSS.n11132 0.001007
R13120 VSS.n3721 VSS.n3720 0.001007
R13121 VSS.n6837 VSS.n6836 0.001007
R13122 VSS.n7938 VSS.n7892 0.001007
R13123 VSS.n9183 VSS.n9182 0.001007
R13124 VSS.n9438 VSS.n9437 0.001007
R13125 VSS.n9666 VSS.n9665 0.001007
R13126 VSS.n9661 VSS.n9660 0.001007
R13127 VSS.n8556 VSS.n8555 0.001007
R13128 VSS.n8347 VSS.n8346 0.001007
R13129 VSS.n8678 VSS.n8677 0.001007
R13130 VSS.n8673 VSS.n8672 0.001007
R13131 VSS.n8741 VSS.n8740 0.001007
R13132 VSS.n8746 VSS.n8743 0.001007
R13133 VSS.n8785 VSS.n8209 0.001007
R13134 VSS.n8068 VSS.n8067 0.001007
R13135 VSS.n9977 VSS.n9976 0.001007
R13136 VSS.n9974 VSS.n9973 0.001007
R13137 VSS.n8120 VSS.n8035 0.001007
R13138 VSS.n8869 VSS.n8868 0.001007
R13139 VSS.n8823 VSS.n8177 0.001007
R13140 VSS.n9561 VSS.n7556 0.001007
R13141 VSS.n7558 VSS.n7557 0.001007
R13142 VSS.n7391 VSS.n7390 0.001007
R13143 VSS.n7396 VSS.n7393 0.001007
R13144 VSS.n3932 VSS.n3931 0.001007
R13145 VSS.n3929 VSS.n3926 0.001007
R13146 VSS.n9443 VSS.n9440 0.001007
R13147 VSS.n9315 VSS.n9314 0.001007
R13148 VSS.n9319 VSS.n9318 0.001007
R13149 VSS.n7221 VSS.n7220 0.001007
R13150 VSS.n7188 VSS.n7187 0.001007
R13151 VSS.n7259 VSS.n7209 0.001007
R13152 VSS.n7375 VSS.n7374 0.001007
R13153 VSS.n9186 VSS.n9184 0.001007
R13154 VSS.n7848 VSS.n7819 0.001007
R13155 VSS.n7830 VSS.n7828 0.001007
R13156 VSS.n7734 VSS.n7733 0.001007
R13157 VSS.n7644 VSS.n7643 0.001007
R13158 VSS.n7699 VSS.n7698 0.001007
R13159 VSS.n7703 VSS.n7702 0.001007
R13160 VSS.n9892 VSS.n9891 0.001007
R13161 VSS.n9889 VSS.n9888 0.001007
R13162 VSS.n8929 VSS.n8928 0.001007
R13163 VSS.n6907 VSS.n6906 0.001007
R13164 VSS.n6860 VSS.n6627 0.001007
R13165 VSS.n6980 VSS.n6979 0.001007
R13166 VSS.n6927 VSS.n6579 0.001007
R13167 VSS.n6537 VSS.n6521 0.001007
R13168 VSS.n6532 VSS.n6530 0.001007
R13169 VSS.n6480 VSS.n6290 0.001007
R13170 VSS.n7061 VSS.n7060 0.001007
R13171 VSS.n6454 VSS.n6453 0.001007
R13172 VSS.n6451 VSS.n6450 0.001007
R13173 VSS.n6840 VSS.n6839 0.001007
R13174 VSS.n5890 VSS.n5889 0.001007
R13175 VSS.n5887 VSS.n5884 0.001007
R13176 VSS.n5709 VSS.n5708 0.001007
R13177 VSS.n5706 VSS.n5703 0.001007
R13178 VSS.n5529 VSS.n5528 0.001007
R13179 VSS.n5526 VSS.n5523 0.001007
R13180 VSS.n5349 VSS.n5348 0.001007
R13181 VSS.n5346 VSS.n5343 0.001007
R13182 VSS.n10083 VSS.n10082 0.001007
R13183 VSS.n10080 VSS.n10077 0.001007
R13184 VSS.n4580 VSS.n4579 0.001007
R13185 VSS.n4607 VSS.n4604 0.001007
R13186 VSS.n6075 VSS.n6074 0.001007
R13187 VSS.n10775 VSS.n10774 0.001007
R13188 VSS.n4415 VSS.n4113 0.001007
R13189 VSS.n4403 VSS.n4402 0.001007
R13190 VSS.n4200 VSS.n4188 0.001007
R13191 VSS.n4300 VSS.n4299 0.001007
R13192 VSS.n4303 VSS.n4302 0.001007
R13193 VSS.n1272 VSS.n1271 0.001007
R13194 VSS.n1269 VSS.n1266 0.001007
R13195 VSS.n1341 VSS.n1340 0.001007
R13196 VSS.n1344 VSS.n1343 0.001007
R13197 VSS.n1105 VSS.n1104 0.001007
R13198 VSS.n960 VSS.n959 0.001007
R13199 VSS.n14227 VSS.n14226 0.001007
R13200 VSS.n14156 VSS.n570 0.001007
R13201 VSS.n10673 VSS.n10672 0.001007
R13202 VSS.n606 VSS.n603 0.001007
R13203 VSS.n13133 VSS.n13132 0.001007
R13204 VSS.n12414 VSS.n2479 0.001007
R13205 VSS.n13053 VSS.n13052 0.001007
R13206 VSS.n2457 VSS.n2456 0.001007
R13207 VSS.n13130 VSS.n13129 0.001007
R13208 VSS.n1395 VSS.n1394 0.001007
R13209 VSS.n1171 VSS.n880 0.001007
R13210 VSS.n13716 VSS.n13713 0.001007
R13211 VSS.n13719 VSS.n13718 0.001007
R13212 VSS.n13256 VSS.n13253 0.001007
R13213 VSS.n13251 VSS.n13250 0.001007
R13214 VSS.n1615 VSS.n1614 0.001007
R13215 VSS.n1686 VSS.n1685 0.001007
R13216 VSS.n1465 VSS.n1464 0.001007
R13217 VSS.n13693 VSS.n13670 0.001007
R13218 VSS.n13698 VSS.n13697 0.001007
R13219 VSS.n13903 VSS.n13902 0.001007
R13220 VSS.n13900 VSS.n13899 0.001007
R13221 VSS.n839 VSS.n837 0.001007
R13222 VSS.n2211 VSS.n2210 0.001007
R13223 VSS.n2215 VSS.n2214 0.001007
R13224 VSS.n2127 VSS.n2126 0.001007
R13225 VSS.n2131 VSS.n2130 0.001007
R13226 VSS.n12649 VSS.n1850 0.001007
R13227 VSS.n13196 VSS.n13195 0.001007
R13228 VSS.n12687 VSS.n12686 0.001007
R13229 VSS.n13924 VSS.n13923 0.001007
R13230 VSS.n1980 VSS.n1979 0.001007
R13231 VSS.n2717 VSS.n2716 0.001007
R13232 VSS.n2665 VSS.n2664 0.001007
R13233 VSS.n2810 VSS.n2787 0.001007
R13234 VSS.n2815 VSS.n2814 0.001007
R13235 VSS.n2897 VSS.n2896 0.001007
R13236 VSS.n2846 VSS.n2845 0.001007
R13237 VSS.n12634 VSS.n3054 0.001007
R13238 VSS.n12639 VSS.n12638 0.001007
R13239 VSS.n3078 VSS.n3077 0.001007
R13240 VSS.n12719 VSS.n12718 0.001007
R13241 VSS.n2608 VSS.n2607 0.001007
R13242 VSS.n12251 VSS.n12250 0.001007
R13243 VSS.n12248 VSS.n12245 0.001007
R13244 VSS.n12144 VSS.n12143 0.001007
R13245 VSS.n12141 VSS.n12138 0.001007
R13246 VSS.n11976 VSS.n11975 0.001007
R13247 VSS.n11973 VSS.n11970 0.001007
R13248 VSS.n3548 VSS.n3547 0.001007
R13249 VSS.n3545 VSS.n3542 0.001007
R13250 VSS.n12600 VSS.n12599 0.001007
R13251 VSS.n12597 VSS.n12594 0.001007
R13252 VSS.n3120 VSS.n3119 0.001007
R13253 VSS.n3141 VSS.n3138 0.001007
R13254 VSS.n11625 VSS.n11624 0.001007
R13255 VSS.n13334 VSS.n13333 0.001007
R13256 VSS.n13340 VSS.n13339 0.001007
R13257 VSS.n13346 VSS.n13345 0.001007
R13258 VSS.n13446 VSS.n13443 0.001007
R13259 VSS.n13436 VSS.n13433 0.001007
R13260 VSS.n13409 VSS.n13406 0.001007
R13261 VSS.n13475 VSS.n13474 0.001007
R13262 VSS.n13472 VSS.n13469 0.001007
R13263 VSS.n13466 VSS.n13463 0.001007
R13264 VSS.n13568 VSS.n13567 0.001007
R13265 VSS.n13561 VSS.n13560 0.001007
R13266 VSS.n13577 VSS.n13576 0.001007
R13267 VSS.n13495 VSS.n13488 0.001007
R13268 VSS.n13486 VSS.n13483 0.001007
R13269 VSS.n13604 VSS.n13484 0.001007
R13270 VSS.n13506 VSS.n13501 0.001007
R13271 VSS.n13602 VSS.n13505 0.001007
R13272 VSS.n13593 VSS.n13504 0.001007
R13273 VSS.n13951 VSS.n13950 0.001007
R13274 VSS.n13957 VSS.n13956 0.001007
R13275 VSS.n13960 VSS.n13959 0.001007
R13276 VSS.n1730 VSS.n1723 0.001007
R13277 VSS.n1721 VSS.n1718 0.001007
R13278 VSS.n14017 VSS.n1719 0.001007
R13279 VSS.n1741 VSS.n1736 0.001007
R13280 VSS.n14015 VSS.n1740 0.001007
R13281 VSS.n14006 VSS.n1739 0.001007
R13282 VSS.n12744 VSS.n12743 0.001007
R13283 VSS.n12747 VSS.n12746 0.001007
R13284 VSS.n12754 VSS.n12753 0.001007
R13285 VSS.n12768 VSS.n2939 0.001007
R13286 VSS.n12776 VSS.n2937 0.001007
R13287 VSS.n12780 VSS.n2936 0.001007
R13288 VSS.n2942 VSS.n2932 0.001007
R13289 VSS.n12797 VSS.n2934 0.001007
R13290 VSS.n12795 VSS.n12787 0.001007
R13291 VSS.n2605 VSS.n2604 0.001007
R13292 VSS.n2025 VSS.n2024 0.001007
R13293 VSS.n829 VSS.n823 0.001007
R13294 VSS.n834 VSS.n833 0.001007
R13295 VSS.n1437 VSS.n1436 0.001007
R13296 VSS.n1491 VSS.n1490 0.001007
R13297 VSS.n1497 VSS.n1496 0.001007
R13298 VSS.n1607 VSS.n1606 0.001007
R13299 VSS.n4007 VSS.n4006 0.001007
R13300 VSS.n4013 VSS.n4012 0.001007
R13301 VSS.n4021 VSS.n4020 0.001007
R13302 VSS.n4049 VSS.n4046 0.001007
R13303 VSS.n4085 VSS.n4084 0.001007
R13304 VSS.n4039 VSS.n4036 0.001007
R13305 VSS.n4064 VSS.n4061 0.001007
R13306 VSS.n4082 VSS.n4079 0.001007
R13307 VSS.n4076 VSS.n4073 0.001007
R13308 VSS.n7288 VSS.n7287 0.001007
R13309 VSS.n7346 VSS.n7290 0.001007
R13310 VSS.n7345 VSS.n7344 0.001007
R13311 VSS.n10863 VSS.n3902 0.001007
R13312 VSS.n10871 VSS.n3900 0.001007
R13313 VSS.n10875 VSS.n3899 0.001007
R13314 VSS.n3905 VSS.n3895 0.001007
R13315 VSS.n10892 VSS.n3897 0.001007
R13316 VSS.n10890 VSS.n10882 0.001007
R13317 VSS.n10974 VSS.n3874 0.001007
R13318 VSS.n10970 VSS.n3875 0.001007
R13319 VSS.n10981 VSS.n3876 0.001007
R13320 VSS.n10909 VSS.n10908 0.001007
R13321 VSS.n10916 VSS.n10915 0.001007
R13322 VSS.n10948 VSS.n10947 0.001007
R13323 VSS.n10923 VSS.n10922 0.001007
R13324 VSS.n10937 VSS.n10936 0.001007
R13325 VSS.n10934 VSS.n10933 0.001007
R13326 VSS.n6342 VSS.n6341 0.001007
R13327 VSS.n6400 VSS.n6344 0.001007
R13328 VSS.n6399 VSS.n6398 0.001007
R13329 VSS.n11014 VSS.n3834 0.001007
R13330 VSS.n11022 VSS.n3832 0.001007
R13331 VSS.n11026 VSS.n3831 0.001007
R13332 VSS.n3837 VSS.n3827 0.001007
R13333 VSS.n11043 VSS.n3829 0.001007
R13334 VSS.n11041 VSS.n11033 0.001007
R13335 VSS.n3747 VSS.n3746 0.001007
R13336 VSS.n3753 VSS.n3752 0.001007
R13337 VSS.n11130 VSS.n11129 0.001007
R13338 VSS.n6829 VSS.n6828 0.001007
R13339 VSS.n7925 VSS.n7889 0.001007
R13340 VSS.n7930 VSS.n7890 0.001007
R13341 VSS.n7934 VSS.n7891 0.001007
R13342 VSS.n9176 VSS.n9170 0.001007
R13343 VSS.n9181 VSS.n9180 0.001007
R13344 VSS.n9267 VSS.n9266 0.001007
R13345 VSS.n9345 VSS.n9344 0.001007
R13346 VSS.n9351 VSS.n9350 0.001007
R13347 VSS.n9435 VSS.n9434 0.001007
R13348 VSS.n9678 VSS.n9677 0.001007
R13349 VSS.n9672 VSS.n9671 0.001007
R13350 VSS.n9692 VSS.n9691 0.001007
R13351 VSS.n9133 VSS.n9130 0.001007
R13352 VSS.n9127 VSS.n9124 0.001007
R13353 VSS.n9030 VSS.n9027 0.001007
R13354 VSS.n9139 VSS.n9138 0.001007
R13355 VSS.n9046 VSS.n9043 0.001007
R13356 VSS.n9040 VSS.n9037 0.001007
R13357 VSS.n9658 VSS.n9655 0.001007
R13358 VSS.n9652 VSS.n9649 0.001007
R13359 VSS.n9689 VSS.n9686 0.001007
R13360 VSS.n8272 VSS.n8271 0.001007
R13361 VSS.n8276 VSS.n8264 0.001007
R13362 VSS.n8282 VSS.n8278 0.001007
R13363 VSS.n8280 VSS.n8279 0.001007
R13364 VSS.n9552 VSS.n9551 0.001007
R13365 VSS.n7576 VSS.n7575 0.001007
R13366 VSS.n7583 VSS.n7582 0.001007
R13367 VSS.n8497 VSS.n8179 0.001007
R13368 VSS.n8501 VSS.n8180 0.001007
R13369 VSS.n8506 VSS.n8181 0.001007
R13370 VSS.n8184 VSS.n8182 0.001007
R13371 VSS.n8357 VSS.n8356 0.001007
R13372 VSS.n8363 VSS.n8362 0.001007
R13373 VSS.n8559 VSS.n8558 0.001007
R13374 VSS.n8455 VSS.n8452 0.001007
R13375 VSS.n8440 VSS.n8437 0.001007
R13376 VSS.n8445 VSS.n8442 0.001007
R13377 VSS.n8468 VSS.n8465 0.001007
R13378 VSS.n8484 VSS.n8483 0.001007
R13379 VSS.n8478 VSS.n8475 0.001007
R13380 VSS.n8376 VSS.n8375 0.001007
R13381 VSS.n8380 VSS.n8368 0.001007
R13382 VSS.n8386 VSS.n8382 0.001007
R13383 VSS.n8384 VSS.n8383 0.001007
R13384 VSS.n8814 VSS.n8813 0.001007
R13385 VSS.n8807 VSS.n8798 0.001007
R13386 VSS.n8805 VSS.n8804 0.001007
R13387 VSS.n8396 VSS.n8211 0.001007
R13388 VSS.n8400 VSS.n8212 0.001007
R13389 VSS.n8405 VSS.n8213 0.001007
R13390 VSS.n8216 VSS.n8214 0.001007
R13391 VSS.n8690 VSS.n8689 0.001007
R13392 VSS.n8684 VSS.n8683 0.001007
R13393 VSS.n8704 VSS.n8703 0.001007
R13394 VSS.n9630 VSS.n9627 0.001007
R13395 VSS.n9636 VSS.n9635 0.001007
R13396 VSS.n7531 VSS.n7528 0.001007
R13397 VSS.n9618 VSS.n9615 0.001007
R13398 VSS.n7547 VSS.n7544 0.001007
R13399 VSS.n7541 VSS.n7538 0.001007
R13400 VSS.n8670 VSS.n8667 0.001007
R13401 VSS.n8664 VSS.n8661 0.001007
R13402 VSS.n8701 VSS.n8698 0.001007
R13403 VSS.n8311 VSS.n8310 0.001007
R13404 VSS.n8317 VSS.n8316 0.001007
R13405 VSS.n8738 VSS.n8737 0.001007
R13406 VSS.n8587 VSS.n8584 0.001007
R13407 VSS.n8581 VSS.n8578 0.001007
R13408 VSS.n8617 VSS.n8616 0.001007
R13409 VSS.n8575 VSS.n8572 0.001007
R13410 VSS.n8612 VSS.n8609 0.001007
R13411 VSS.n8605 VSS.n8602 0.001007
R13412 VSS.n8599 VSS.n8596 0.001007
R13413 VSS.n8301 VSS.n8298 0.001007
R13414 VSS.n8295 VSS.n8292 0.001007
R13415 VSS.n8751 VSS.n8750 0.001007
R13416 VSS.n8258 VSS.n8255 0.001007
R13417 VSS.n8256 VSS.n8244 0.001007
R13418 VSS.n8777 VSS.n8776 0.001007
R13419 VSS.n8240 VSS.n8239 0.001007
R13420 VSS.n8234 VSS.n8224 0.001007
R13421 VSS.n8232 VSS.n8231 0.001007
R13422 VSS.n8789 VSS.n8198 0.001007
R13423 VSS.n8208 VSS.n8200 0.001007
R13424 VSS.n8787 VSS.n8196 0.001007
R13425 VSS.n6199 VSS.n6196 0.001007
R13426 VSS.n6205 VSS.n6204 0.001007
R13427 VSS.n6189 VSS.n6186 0.001007
R13428 VSS.n6166 VSS.n6163 0.001007
R13429 VSS.n6161 VSS.n6158 0.001007
R13430 VSS.n6176 VSS.n6173 0.001007
R13431 VSS.n9980 VSS.n9979 0.001007
R13432 VSS.n6222 VSS.n6217 0.001007
R13433 VSS.n6220 VSS.n6218 0.001007
R13434 VSS.n6756 VSS.n6714 0.001007
R13435 VSS.n6752 VSS.n6713 0.001007
R13436 VSS.n6748 VSS.n6712 0.001007
R13437 VSS.n6744 VSS.n6698 0.001007
R13438 VSS.n6764 VSS.n6695 0.001007
R13439 VSS.n6762 VSS.n6696 0.001007
R13440 VSS.n6709 VSS.n6700 0.001007
R13441 VSS.n9966 VSS.n9965 0.001007
R13442 VSS.n9960 VSS.n9959 0.001007
R13443 VSS.n9969 VSS.n9968 0.001007
R13444 VSS.n8028 VSS.n8021 0.001007
R13445 VSS.n8033 VSS.n8032 0.001007
R13446 VSS.n8154 VSS.n8019 0.001007
R13447 VSS.n8152 VSS.n8151 0.001007
R13448 VSS.n8109 VSS.n8094 0.001007
R13449 VSS.n8105 VSS.n8093 0.001007
R13450 VSS.n8101 VSS.n8092 0.001007
R13451 VSS.n8042 VSS.n8041 0.001007
R13452 VSS.n8091 VSS.n8090 0.001007
R13453 VSS.n8084 VSS.n8045 0.001007
R13454 VSS.n8080 VSS.n8044 0.001007
R13455 VSS.n8142 VSS.n8141 0.001007
R13456 VSS.n8137 VSS.n8130 0.001007
R13457 VSS.n8128 VSS.n8127 0.001007
R13458 VSS.n8071 VSS.n8070 0.001007
R13459 VSS.n8065 VSS.n8064 0.001007
R13460 VSS.n8060 VSS.n8059 0.001007
R13461 VSS.n8888 VSS.n7971 0.001007
R13462 VSS.n8884 VSS.n7970 0.001007
R13463 VSS.n8880 VSS.n7969 0.001007
R13464 VSS.n8876 VSS.n7955 0.001007
R13465 VSS.n8896 VSS.n7951 0.001007
R13466 VSS.n8894 VSS.n7952 0.001007
R13467 VSS.n7966 VSS.n7957 0.001007
R13468 VSS.n8861 VSS.n8860 0.001007
R13469 VSS.n8858 VSS.n8857 0.001007
R13470 VSS.n8866 VSS.n8865 0.001007
R13471 VSS.n8827 VSS.n8166 0.001007
R13472 VSS.n8176 VSS.n8168 0.001007
R13473 VSS.n8825 VSS.n8164 0.001007
R13474 VSS.n9581 VSS.n9579 0.001007
R13475 VSS.n9565 VSS.n7559 0.001007
R13476 VSS.n9569 VSS.n7560 0.001007
R13477 VSS.n7563 VSS.n7561 0.001007
R13478 VSS.n9590 VSS.n9589 0.001007
R13479 VSS.n9593 VSS.n9592 0.001007
R13480 VSS.n8535 VSS.n8532 0.001007
R13481 VSS.n8541 VSS.n8538 0.001007
R13482 VSS.n8547 VSS.n8544 0.001007
R13483 VSS.n9387 VSS.n9384 0.001007
R13484 VSS.n9381 VSS.n9378 0.001007
R13485 VSS.n9417 VSS.n9416 0.001007
R13486 VSS.n9375 VSS.n9372 0.001007
R13487 VSS.n9412 VSS.n9409 0.001007
R13488 VSS.n9405 VSS.n9402 0.001007
R13489 VSS.n9399 VSS.n9396 0.001007
R13490 VSS.n7388 VSS.n7387 0.001007
R13491 VSS.n9789 VSS.n9788 0.001007
R13492 VSS.n7402 VSS.n7399 0.001007
R13493 VSS.n7408 VSS.n7405 0.001007
R13494 VSS.n7418 VSS.n7415 0.001007
R13495 VSS.n9782 VSS.n9779 0.001007
R13496 VSS.n7444 VSS.n7441 0.001007
R13497 VSS.n7438 VSS.n7435 0.001007
R13498 VSS.n7474 VSS.n7473 0.001007
R13499 VSS.n7432 VSS.n7429 0.001007
R13500 VSS.n7469 VSS.n7466 0.001007
R13501 VSS.n7462 VSS.n7459 0.001007
R13502 VSS.n7456 VSS.n7453 0.001007
R13503 VSS.n3924 VSS.n3923 0.001007
R13504 VSS.n10836 VSS.n10835 0.001007
R13505 VSS.n3938 VSS.n3935 0.001007
R13506 VSS.n3944 VSS.n3941 0.001007
R13507 VSS.n3954 VSS.n3951 0.001007
R13508 VSS.n10829 VSS.n10826 0.001007
R13509 VSS.n9081 VSS.n9078 0.001007
R13510 VSS.n9075 VSS.n9072 0.001007
R13511 VSS.n9111 VSS.n9110 0.001007
R13512 VSS.n9069 VSS.n9066 0.001007
R13513 VSS.n9106 VSS.n9103 0.001007
R13514 VSS.n9099 VSS.n9096 0.001007
R13515 VSS.n9093 VSS.n9090 0.001007
R13516 VSS.n9335 VSS.n9332 0.001007
R13517 VSS.n9329 VSS.n9326 0.001007
R13518 VSS.n9448 VSS.n9447 0.001007
R13519 VSS.n9277 VSS.n9003 0.001007
R13520 VSS.n9282 VSS.n9002 0.001007
R13521 VSS.n9286 VSS.n9001 0.001007
R13522 VSS.n9289 VSS.n9000 0.001007
R13523 VSS.n9015 VSS.n8996 0.001007
R13524 VSS.n9517 VSS.n8998 0.001007
R13525 VSS.n9014 VSS.n9006 0.001007
R13526 VSS.n9493 VSS.n9491 0.001007
R13527 VSS.n9310 VSS.n9292 0.001007
R13528 VSS.n9308 VSS.n9307 0.001007
R13529 VSS.n9302 VSS.n9301 0.001007
R13530 VSS.n9503 VSS.n9502 0.001007
R13531 VSS.n9506 VSS.n9505 0.001007
R13532 VSS.n7237 VSS.n7236 0.001007
R13533 VSS.n7226 VSS.n7225 0.001007
R13534 VSS.n7234 VSS.n7233 0.001007
R13535 VSS.n9474 VSS.n7167 0.001007
R13536 VSS.n9477 VSS.n7166 0.001007
R13537 VSS.n9478 VSS.n7165 0.001007
R13538 VSS.n7182 VSS.n7164 0.001007
R13539 VSS.n7179 VSS.n7160 0.001007
R13540 VSS.n9839 VSS.n7162 0.001007
R13541 VSS.n7178 VSS.n7170 0.001007
R13542 VSS.n9824 VSS.n9823 0.001007
R13543 VSS.n9818 VSS.n9817 0.001007
R13544 VSS.n9828 VSS.n9827 0.001007
R13545 VSS.n7200 VSS.n7195 0.001007
R13546 VSS.n7207 VSS.n7206 0.001007
R13547 VSS.n7257 VSS.n7256 0.001007
R13548 VSS.n7214 VSS.n7213 0.001007
R13549 VSS.n7249 VSS.n7248 0.001007
R13550 VSS.n7356 VSS.n7273 0.001007
R13551 VSS.n7360 VSS.n7274 0.001007
R13552 VSS.n7267 VSS.n7266 0.001007
R13553 VSS.n7316 VSS.n7271 0.001007
R13554 VSS.n7326 VSS.n7270 0.001007
R13555 VSS.n7319 VSS.n7269 0.001007
R13556 VSS.n7193 VSS.n7192 0.001007
R13557 VSS.n9193 VSS.n9191 0.001007
R13558 VSS.n9203 VSS.n9202 0.001007
R13559 VSS.n9204 VSS.n9189 0.001007
R13560 VSS.n9212 VSS.n9211 0.001007
R13561 VSS.n9238 VSS.n9237 0.001007
R13562 VSS.n9220 VSS.n9219 0.001007
R13563 VSS.n9227 VSS.n9226 0.001007
R13564 VSS.n9256 VSS.n9168 0.001007
R13565 VSS.n9251 VSS.n9167 0.001007
R13566 VSS.n9264 VSS.n9185 0.001007
R13567 VSS.n8960 VSS.n8959 0.001007
R13568 VSS.n7845 VSS.n7826 0.001007
R13569 VSS.n7825 VSS.n7820 0.001007
R13570 VSS.n7903 VSS.n7897 0.001007
R13571 VSS.n7906 VSS.n7905 0.001007
R13572 VSS.n7913 VSS.n7912 0.001007
R13573 VSS.n7910 VSS.n7909 0.001007
R13574 VSS.n8945 VSS.n8944 0.001007
R13575 VSS.n7859 VSS.n7858 0.001007
R13576 VSS.n7866 VSS.n7865 0.001007
R13577 VSS.n7840 VSS.n7817 0.001007
R13578 VSS.n7835 VSS.n7816 0.001007
R13579 VSS.n8957 VSS.n7829 0.001007
R13580 VSS.n7750 VSS.n7749 0.001007
R13581 VSS.n7739 VSS.n7738 0.001007
R13582 VSS.n7747 VSS.n7746 0.001007
R13583 VSS.n7622 VSS.n7619 0.001007
R13584 VSS.n7618 VSS.n7613 0.001007
R13585 VSS.n8986 VSS.n7615 0.001007
R13586 VSS.n7637 VSS.n7617 0.001007
R13587 VSS.n8967 VSS.n7630 0.001007
R13588 VSS.n8968 VSS.n7629 0.001007
R13589 VSS.n8972 VSS.n7628 0.001007
R13590 VSS.n7797 VSS.n7796 0.001007
R13591 VSS.n7791 VSS.n7790 0.001007
R13592 VSS.n7801 VSS.n7800 0.001007
R13593 VSS.n7691 VSS.n7690 0.001007
R13594 VSS.n7678 VSS.n7676 0.001007
R13595 VSS.n7682 VSS.n7679 0.001007
R13596 VSS.n7657 VSS.n7654 0.001007
R13597 VSS.n7653 VSS.n7648 0.001007
R13598 VSS.n7776 VSS.n7650 0.001007
R13599 VSS.n7672 VSS.n7652 0.001007
R13600 VSS.n7757 VSS.n7665 0.001007
R13601 VSS.n7758 VSS.n7664 0.001007
R13602 VSS.n7762 VSS.n7663 0.001007
R13603 VSS.n7718 VSS.n7717 0.001007
R13604 VSS.n7712 VSS.n7711 0.001007
R13605 VSS.n7722 VSS.n7721 0.001007
R13606 VSS.n9875 VSS.n9874 0.001007
R13607 VSS.n9881 VSS.n9880 0.001007
R13608 VSS.n9895 VSS.n9894 0.001007
R13609 VSS.n7079 VSS.n7074 0.001007
R13610 VSS.n7077 VSS.n7075 0.001007
R13611 VSS.n7125 VSS.n7117 0.001007
R13612 VSS.n7130 VSS.n7118 0.001007
R13613 VSS.n7094 VSS.n7093 0.001007
R13614 VSS.n7115 VSS.n7114 0.001007
R13615 VSS.n7109 VSS.n7097 0.001007
R13616 VSS.n7102 VSS.n7096 0.001007
R13617 VSS.n9884 VSS.n9883 0.001007
R13618 VSS.n7982 VSS.n7981 0.001007
R13619 VSS.n7991 VSS.n7990 0.001007
R13620 VSS.n7996 VSS.n7995 0.001007
R13621 VSS.n8920 VSS.n8919 0.001007
R13622 VSS.n8913 VSS.n8904 0.001007
R13623 VSS.n8911 VSS.n8910 0.001007
R13624 VSS.n8933 VSS.n7876 0.001007
R13625 VSS.n7887 VSS.n7879 0.001007
R13626 VSS.n8931 VSS.n7874 0.001007
R13627 VSS.n6800 VSS.n6637 0.001007
R13628 VSS.n6803 VSS.n6636 0.001007
R13629 VSS.n6804 VSS.n6635 0.001007
R13630 VSS.n6634 VSS.n6633 0.001007
R13631 VSS.n6853 VSS.n6852 0.001007
R13632 VSS.n6646 VSS.n6641 0.001007
R13633 VSS.n6647 VSS.n6640 0.001007
R13634 VSS.n6896 VSS.n6895 0.001007
R13635 VSS.n6900 VSS.n6899 0.001007
R13636 VSS.n6910 VSS.n6909 0.001007
R13637 VSS.n6625 VSS.n6624 0.001007
R13638 VSS.n6620 VSS.n6614 0.001007
R13639 VSS.n6890 VSS.n6889 0.001007
R13640 VSS.n6868 VSS.n6589 0.001007
R13641 VSS.n6871 VSS.n6588 0.001007
R13642 VSS.n6872 VSS.n6587 0.001007
R13643 VSS.n6586 VSS.n6585 0.001007
R13644 VSS.n6920 VSS.n6919 0.001007
R13645 VSS.n6598 VSS.n6593 0.001007
R13646 VSS.n6599 VSS.n6592 0.001007
R13647 VSS.n6969 VSS.n6968 0.001007
R13648 VSS.n6973 VSS.n6972 0.001007
R13649 VSS.n6983 VSS.n6982 0.001007
R13650 VSS.n6577 VSS.n6576 0.001007
R13651 VSS.n6572 VSS.n6566 0.001007
R13652 VSS.n6963 VSS.n6962 0.001007
R13653 VSS.n7042 VSS.n7041 0.001007
R13654 VSS.n6534 VSS.n6528 0.001007
R13655 VSS.n6527 VSS.n6522 0.001007
R13656 VSS.n6938 VSS.n6932 0.001007
R13657 VSS.n6941 VSS.n6940 0.001007
R13658 VSS.n6948 VSS.n6947 0.001007
R13659 VSS.n6945 VSS.n6944 0.001007
R13660 VSS.n6993 VSS.n6992 0.001007
R13661 VSS.n6548 VSS.n6547 0.001007
R13662 VSS.n6555 VSS.n6554 0.001007
R13663 VSS.n7011 VSS.n6519 0.001007
R13664 VSS.n7005 VSS.n6518 0.001007
R13665 VSS.n7039 VSS.n6531 0.001007
R13666 VSS.n6465 VSS.n6294 0.001007
R13667 VSS.n6478 VSS.n6477 0.001007
R13668 VSS.n6470 VSS.n6469 0.001007
R13669 VSS.n7021 VSS.n6491 0.001007
R13670 VSS.n7024 VSS.n6490 0.001007
R13671 VSS.n7025 VSS.n6489 0.001007
R13672 VSS.n6488 VSS.n6487 0.001007
R13673 VSS.n7052 VSS.n7051 0.001007
R13674 VSS.n6500 VSS.n6495 0.001007
R13675 VSS.n6501 VSS.n6494 0.001007
R13676 VSS.n6288 VSS.n6286 0.001007
R13677 VSS.n6282 VSS.n6276 0.001007
R13678 VSS.n6274 VSS.n6273 0.001007
R13679 VSS.n6437 VSS.n6436 0.001007
R13680 VSS.n6443 VSS.n6442 0.001007
R13681 VSS.n6457 VSS.n6456 0.001007
R13682 VSS.n6306 VSS.n6301 0.001007
R13683 VSS.n6304 VSS.n6302 0.001007
R13684 VSS.n6410 VSS.n6327 0.001007
R13685 VSS.n6414 VSS.n6328 0.001007
R13686 VSS.n6321 VSS.n6320 0.001007
R13687 VSS.n6370 VSS.n6325 0.001007
R13688 VSS.n6380 VSS.n6324 0.001007
R13689 VSS.n6373 VSS.n6323 0.001007
R13690 VSS.n6446 VSS.n6445 0.001007
R13691 VSS.n6823 VSS.n6822 0.001007
R13692 VSS.n6832 VSS.n6831 0.001007
R13693 VSS.n6722 VSS.n6681 0.001007
R13694 VSS.n6728 VSS.n6682 0.001007
R13695 VSS.n6734 VSS.n6683 0.001007
R13696 VSS.n6785 VSS.n6784 0.001007
R13697 VSS.n6778 VSS.n6687 0.001007
R13698 VSS.n6774 VSS.n6686 0.001007
R13699 VSS.n6673 VSS.n6672 0.001007
R13700 VSS.n6668 VSS.n6662 0.001007
R13701 VSS.n6843 VSS.n6842 0.001007
R13702 VSS.n6014 VSS.n6011 0.001007
R13703 VSS.n6008 VSS.n6005 0.001007
R13704 VSS.n6044 VSS.n6043 0.001007
R13705 VSS.n6002 VSS.n5999 0.001007
R13706 VSS.n6039 VSS.n6036 0.001007
R13707 VSS.n6032 VSS.n6029 0.001007
R13708 VSS.n6026 VSS.n6023 0.001007
R13709 VSS.n5860 VSS.n5859 0.001007
R13710 VSS.n5854 VSS.n5853 0.001007
R13711 VSS.n5899 VSS.n5898 0.001007
R13712 VSS.n5882 VSS.n5879 0.001007
R13713 VSS.n5876 VSS.n5873 0.001007
R13714 VSS.n5866 VSS.n5863 0.001007
R13715 VSS.n5816 VSS.n5813 0.001007
R13716 VSS.n5810 VSS.n5807 0.001007
R13717 VSS.n5846 VSS.n5845 0.001007
R13718 VSS.n5804 VSS.n5801 0.001007
R13719 VSS.n5841 VSS.n5838 0.001007
R13720 VSS.n5834 VSS.n5831 0.001007
R13721 VSS.n5828 VSS.n5825 0.001007
R13722 VSS.n5679 VSS.n5678 0.001007
R13723 VSS.n5673 VSS.n5672 0.001007
R13724 VSS.n5718 VSS.n5717 0.001007
R13725 VSS.n5701 VSS.n5698 0.001007
R13726 VSS.n5695 VSS.n5692 0.001007
R13727 VSS.n5685 VSS.n5682 0.001007
R13728 VSS.n5635 VSS.n5632 0.001007
R13729 VSS.n5629 VSS.n5626 0.001007
R13730 VSS.n5665 VSS.n5664 0.001007
R13731 VSS.n5623 VSS.n5620 0.001007
R13732 VSS.n5660 VSS.n5657 0.001007
R13733 VSS.n5653 VSS.n5650 0.001007
R13734 VSS.n5647 VSS.n5644 0.001007
R13735 VSS.n5499 VSS.n5498 0.001007
R13736 VSS.n5493 VSS.n5492 0.001007
R13737 VSS.n5538 VSS.n5537 0.001007
R13738 VSS.n5521 VSS.n5518 0.001007
R13739 VSS.n5515 VSS.n5512 0.001007
R13740 VSS.n5505 VSS.n5502 0.001007
R13741 VSS.n5455 VSS.n5452 0.001007
R13742 VSS.n5449 VSS.n5446 0.001007
R13743 VSS.n5485 VSS.n5484 0.001007
R13744 VSS.n5443 VSS.n5440 0.001007
R13745 VSS.n5480 VSS.n5477 0.001007
R13746 VSS.n5473 VSS.n5470 0.001007
R13747 VSS.n5467 VSS.n5464 0.001007
R13748 VSS.n5319 VSS.n5318 0.001007
R13749 VSS.n5313 VSS.n5312 0.001007
R13750 VSS.n5358 VSS.n5357 0.001007
R13751 VSS.n5341 VSS.n5338 0.001007
R13752 VSS.n5335 VSS.n5332 0.001007
R13753 VSS.n5325 VSS.n5322 0.001007
R13754 VSS.n5275 VSS.n5272 0.001007
R13755 VSS.n5269 VSS.n5266 0.001007
R13756 VSS.n5305 VSS.n5304 0.001007
R13757 VSS.n5263 VSS.n5260 0.001007
R13758 VSS.n5300 VSS.n5297 0.001007
R13759 VSS.n5293 VSS.n5290 0.001007
R13760 VSS.n5287 VSS.n5284 0.001007
R13761 VSS.n10053 VSS.n10052 0.001007
R13762 VSS.n10047 VSS.n10046 0.001007
R13763 VSS.n10092 VSS.n10091 0.001007
R13764 VSS.n10075 VSS.n10072 0.001007
R13765 VSS.n10069 VSS.n10066 0.001007
R13766 VSS.n10059 VSS.n10056 0.001007
R13767 VSS.n4617 VSS.n4616 0.001007
R13768 VSS.n4623 VSS.n4622 0.001007
R13769 VSS.n4586 VSS.n4583 0.001007
R13770 VSS.n4592 VSS.n4589 0.001007
R13771 VSS.n4598 VSS.n4595 0.001007
R13772 VSS.n3802 VSS.n3799 0.001007
R13773 VSS.n3808 VSS.n3805 0.001007
R13774 VSS.n3765 VSS.n3762 0.001007
R13775 VSS.n3790 VSS.n3787 0.001007
R13776 VSS.n3781 VSS.n3778 0.001007
R13777 VSS.n3775 VSS.n3772 0.001007
R13778 VSS.n4628 VSS.n4627 0.001007
R13779 VSS.n6067 VSS.n6066 0.001007
R13780 VSS.n6081 VSS.n6080 0.001007
R13781 VSS.n5986 VSS.n5985 0.001007
R13782 VSS.n5980 VSS.n5979 0.001007
R13783 VSS.n6061 VSS.n6058 0.001007
R13784 VSS.n6055 VSS.n6052 0.001007
R13785 VSS.n6072 VSS.n6069 0.001007
R13786 VSS.n11066 VSS.n11063 0.001007
R13787 VSS.n11109 VSS.n11108 0.001007
R13788 VSS.n11056 VSS.n11053 0.001007
R13789 VSS.n11088 VSS.n11085 0.001007
R13790 VSS.n11106 VSS.n11103 0.001007
R13791 VSS.n11100 VSS.n11097 0.001007
R13792 VSS.n11138 VSS.n11137 0.001007
R13793 VSS.n3727 VSS.n3724 0.001007
R13794 VSS.n3733 VSS.n3730 0.001007
R13795 VSS.n6349 VSS.n6348 0.001007
R13796 VSS.n6354 VSS.n6353 0.001007
R13797 VSS.n6361 VSS.n6360 0.001007
R13798 VSS.n3862 VSS.n3855 0.001007
R13799 VSS.n10988 VSS.n3857 0.001007
R13800 VSS.n3865 VSS.n3863 0.001007
R13801 VSS.n7295 VSS.n7294 0.001007
R13802 VSS.n7300 VSS.n7299 0.001007
R13803 VSS.n7307 VSS.n7306 0.001007
R13804 VSS.n3981 VSS.n3978 0.001007
R13805 VSS.n3987 VSS.n3984 0.001007
R13806 VSS.n3993 VSS.n3990 0.001007
R13807 VSS.n4126 VSS.n4125 0.001007
R13808 VSS.n10777 VSS.n4110 0.001007
R13809 VSS.n4127 VSS.n4112 0.001007
R13810 VSS.n4222 VSS.n4196 0.001007
R13811 VSS.n10757 VSS.n10756 0.001007
R13812 VSS.n10767 VSS.n10764 0.001007
R13813 VSS.n10765 VSS.n4453 0.001007
R13814 VSS.n4447 VSS.n4446 0.001007
R13815 VSS.n4149 VSS.n4140 0.001007
R13816 VSS.n4147 VSS.n4146 0.001007
R13817 VSS.n4398 VSS.n4193 0.001007
R13818 VSS.n4394 VSS.n4192 0.001007
R13819 VSS.n4389 VSS.n4191 0.001007
R13820 VSS.n4171 VSS.n4168 0.001007
R13821 VSS.n4173 VSS.n4167 0.001007
R13822 VSS.n4166 VSS.n4164 0.001007
R13823 VSS.n4406 VSS.n4165 0.001007
R13824 VSS.n4379 VSS.n4183 0.001007
R13825 VSS.n4362 VSS.n4182 0.001007
R13826 VSS.n4366 VSS.n4185 0.001007
R13827 VSS.n4286 VSS.n4285 0.001007
R13828 VSS.n4292 VSS.n4291 0.001007
R13829 VSS.n4295 VSS.n4294 0.001007
R13830 VSS.n4244 VSS.n4237 0.001007
R13831 VSS.n4235 VSS.n4232 0.001007
R13832 VSS.n4345 VSS.n4233 0.001007
R13833 VSS.n4255 VSS.n4250 0.001007
R13834 VSS.n4343 VSS.n4254 0.001007
R13835 VSS.n4334 VSS.n4253 0.001007
R13836 VSS.n4306 VSS.n4305 0.001007
R13837 VSS.n4319 VSS.n4318 0.001007
R13838 VSS.n4309 VSS.n4308 0.001007
R13839 VSS.n4211 VSS.n4194 0.001007
R13840 VSS.n4218 VSS.n4189 0.001007
R13841 VSS.n4418 VSS.n4115 0.001007
R13842 VSS.n4419 VSS.n4116 0.001007
R13843 VSS.n4420 VSS.n4117 0.001007
R13844 VSS.n1284 VSS.n1283 0.001007
R13845 VSS.n1278 VSS.n1277 0.001007
R13846 VSS.n1298 VSS.n1297 0.001007
R13847 VSS.n786 VSS.n783 0.001007
R13848 VSS.n780 VSS.n777 0.001007
R13849 VSS.n664 VSS.n661 0.001007
R13850 VSS.n792 VSS.n791 0.001007
R13851 VSS.n680 VSS.n677 0.001007
R13852 VSS.n674 VSS.n671 0.001007
R13853 VSS.n1264 VSS.n1261 0.001007
R13854 VSS.n1258 VSS.n1255 0.001007
R13855 VSS.n1295 VSS.n1292 0.001007
R13856 VSS.n1222 VSS.n1221 0.001007
R13857 VSS.n1228 VSS.n1227 0.001007
R13858 VSS.n1336 VSS.n1335 0.001007
R13859 VSS.n1019 VSS.n1016 0.001007
R13860 VSS.n1013 VSS.n1010 0.001007
R13861 VSS.n1049 VSS.n1048 0.001007
R13862 VSS.n1007 VSS.n1004 0.001007
R13863 VSS.n1044 VSS.n1041 0.001007
R13864 VSS.n1037 VSS.n1034 0.001007
R13865 VSS.n1031 VSS.n1028 0.001007
R13866 VSS.n1212 VSS.n1209 0.001007
R13867 VSS.n1206 VSS.n1203 0.001007
R13868 VSS.n1349 VSS.n1348 0.001007
R13869 VSS.n943 VSS.n890 0.001007
R13870 VSS.n947 VSS.n889 0.001007
R13871 VSS.n952 VSS.n888 0.001007
R13872 VSS.n887 VSS.n886 0.001007
R13873 VSS.n1164 VSS.n1163 0.001007
R13874 VSS.n899 VSS.n894 0.001007
R13875 VSS.n900 VSS.n893 0.001007
R13876 VSS.n596 VSS.n589 0.001007
R13877 VSS.n601 VSS.n600 0.001007
R13878 VSS.n14204 VSS.n587 0.001007
R13879 VSS.n14202 VSS.n14201 0.001007
R13880 VSS.n970 VSS.n969 0.001007
R13881 VSS.n976 VSS.n975 0.001007
R13882 VSS.n1086 VSS.n1085 0.001007
R13883 VSS.n14299 VSS.n14296 0.001007
R13884 VSS.n14293 VSS.n14290 0.001007
R13885 VSS.n14334 VSS.n14333 0.001007
R13886 VSS.n14287 VSS.n14284 0.001007
R13887 VSS.n14318 VSS.n14315 0.001007
R13888 VSS.n14313 VSS.n14310 0.001007
R13889 VSS.n14328 VSS.n14325 0.001007
R13890 VSS.n14170 VSS.n578 0.001007
R13891 VSS.n14222 VSS.n575 0.001007
R13892 VSS.n14218 VSS.n574 0.001007
R13893 VSS.n14213 VSS.n573 0.001007
R13894 VSS.n562 VSS.n557 0.001007
R13895 VSS.n14232 VSS.n548 0.001007
R13896 VSS.n14230 VSS.n549 0.001007
R13897 VSS.n2402 VSS.n551 0.001007
R13898 VSS.n2406 VSS.n550 0.001007
R13899 VSS.n2411 VSS.n553 0.001007
R13900 VSS.n10681 VSS.n10680 0.001007
R13901 VSS.n10687 VSS.n10686 0.001007
R13902 VSS.n10706 VSS.n10705 0.001007
R13903 VSS.n10692 VSS.n10691 0.001007
R13904 VSS.n14271 VSS.n14268 0.001007
R13905 VSS.n14277 VSS.n14276 0.001007
R13906 VSS.n519 VSS.n516 0.001007
R13907 VSS.n14259 VSS.n14256 0.001007
R13908 VSS.n535 VSS.n532 0.001007
R13909 VSS.n529 VSS.n526 0.001007
R13910 VSS.n10670 VSS.n10667 0.001007
R13911 VSS.n10664 VSS.n10661 0.001007
R13912 VSS.n10703 VSS.n10700 0.001007
R13913 VSS.n1146 VSS.n932 0.001007
R13914 VSS.n1142 VSS.n931 0.001007
R13915 VSS.n1138 VSS.n930 0.001007
R13916 VSS.n1134 VSS.n916 0.001007
R13917 VSS.n1154 VSS.n913 0.001007
R13918 VSS.n1152 VSS.n914 0.001007
R13919 VSS.n927 VSS.n918 0.001007
R13920 VSS.n14192 VSS.n14191 0.001007
R13921 VSS.n14187 VSS.n14180 0.001007
R13922 VSS.n14178 VSS.n14177 0.001007
R13923 VSS.n12450 VSS.n12447 0.001007
R13924 VSS.n12444 VSS.n12441 0.001007
R13925 VSS.n12438 VSS.n12435 0.001007
R13926 VSS.n12394 VSS.n12391 0.001007
R13927 VSS.n12371 VSS.n12368 0.001007
R13928 VSS.n12455 VSS.n12454 0.001007
R13929 VSS.n12381 VSS.n12378 0.001007
R13930 VSS.n12417 VSS.n12416 0.001007
R13931 VSS.n12412 VSS.n12411 0.001007
R13932 VSS.n12407 VSS.n12406 0.001007
R13933 VSS.n13034 VSS.n2493 0.001007
R13934 VSS.n13038 VSS.n2494 0.001007
R13935 VSS.n2487 VSS.n2486 0.001007
R13936 VSS.n2535 VSS.n2491 0.001007
R13937 VSS.n2545 VSS.n2490 0.001007
R13938 VSS.n2538 VSS.n2489 0.001007
R13939 VSS.n2477 VSS.n2476 0.001007
R13940 VSS.n2470 VSS.n2466 0.001007
R13941 VSS.n13056 VSS.n13055 0.001007
R13942 VSS.n2438 VSS.n2432 0.001007
R13943 VSS.n2443 VSS.n2440 0.001007
R13944 VSS.n2441 VSS.n2393 0.001007
R13945 VSS.n2452 VSS.n2451 0.001007
R13946 VSS.n2370 VSS.n2369 0.001007
R13947 VSS.n13103 VSS.n13102 0.001007
R13948 VSS.n2372 VSS.n2358 0.001007
R13949 VSS.n2375 VSS.n2362 0.001007
R13950 VSS.n2385 VSS.n2361 0.001007
R13951 VSS.n2378 VSS.n2360 0.001007
R13952 VSS.n13086 VSS.n13085 0.001007
R13953 VSS.n13081 VSS.n13074 0.001007
R13954 VSS.n13072 VSS.n13071 0.001007
R13955 VSS.n13136 VSS.n13135 0.001007
R13956 VSS.n1920 VSS.n1915 0.001007
R13957 VSS.n1918 VSS.n1916 0.001007
R13958 VSS.n2337 VSS.n1942 0.001007
R13959 VSS.n2333 VSS.n1941 0.001007
R13960 VSS.n2329 VSS.n1940 0.001007
R13961 VSS.n1935 VSS.n1934 0.001007
R13962 VSS.n2294 VSS.n1939 0.001007
R13963 VSS.n2290 VSS.n1938 0.001007
R13964 VSS.n2286 VSS.n1937 0.001007
R13965 VSS.n13122 VSS.n13121 0.001007
R13966 VSS.n13116 VSS.n13115 0.001007
R13967 VSS.n13125 VSS.n13124 0.001007
R13968 VSS.n14159 VSS.n576 0.001007
R13969 VSS.n14166 VSS.n571 0.001007
R13970 VSS.n1375 VSS.n1373 0.001007
R13971 VSS.n1398 VSS.n1397 0.001007
R13972 VSS.n871 VSS.n866 0.001007
R13973 VSS.n869 VSS.n867 0.001007
R13974 VSS.n1385 VSS.n1384 0.001007
R13975 VSS.n1388 VSS.n1387 0.001007
R13976 VSS.n1110 VSS.n1109 0.001007
R13977 VSS.n1092 VSS.n1089 0.001007
R13978 VSS.n1098 VSS.n1095 0.001007
R13979 VSS.n1541 VSS.n1538 0.001007
R13980 VSS.n1535 VSS.n1532 0.001007
R13981 VSS.n1571 VSS.n1570 0.001007
R13982 VSS.n1529 VSS.n1526 0.001007
R13983 VSS.n1566 VSS.n1563 0.001007
R13984 VSS.n1559 VSS.n1556 0.001007
R13985 VSS.n1553 VSS.n1550 0.001007
R13986 VSS.n13711 VSS.n13710 0.001007
R13987 VSS.n13857 VSS.n13856 0.001007
R13988 VSS.n13725 VSS.n13722 0.001007
R13989 VSS.n13731 VSS.n13728 0.001007
R13990 VSS.n13741 VSS.n13738 0.001007
R13991 VSS.n13850 VSS.n13847 0.001007
R13992 VSS.n13781 VSS.n13778 0.001007
R13993 VSS.n13775 VSS.n13772 0.001007
R13994 VSS.n13811 VSS.n13810 0.001007
R13995 VSS.n13769 VSS.n13766 0.001007
R13996 VSS.n13806 VSS.n13803 0.001007
R13997 VSS.n13799 VSS.n13796 0.001007
R13998 VSS.n13793 VSS.n13790 0.001007
R13999 VSS.n13248 VSS.n13247 0.001007
R14000 VSS.n13392 VSS.n13391 0.001007
R14001 VSS.n13262 VSS.n13259 0.001007
R14002 VSS.n13268 VSS.n13265 0.001007
R14003 VSS.n13278 VSS.n13275 0.001007
R14004 VSS.n13385 VSS.n13382 0.001007
R14005 VSS.n734 VSS.n731 0.001007
R14006 VSS.n728 VSS.n725 0.001007
R14007 VSS.n764 VSS.n763 0.001007
R14008 VSS.n722 VSS.n719 0.001007
R14009 VSS.n759 VSS.n756 0.001007
R14010 VSS.n752 VSS.n749 0.001007
R14011 VSS.n746 VSS.n743 0.001007
R14012 VSS.n1481 VSS.n1478 0.001007
R14013 VSS.n1475 VSS.n1472 0.001007
R14014 VSS.n1620 VSS.n1619 0.001007
R14015 VSS.n1447 VSS.n637 0.001007
R14016 VSS.n1452 VSS.n636 0.001007
R14017 VSS.n1456 VSS.n635 0.001007
R14018 VSS.n1459 VSS.n634 0.001007
R14019 VSS.n649 VSS.n630 0.001007
R14020 VSS.n14116 VSS.n632 0.001007
R14021 VSS.n648 VSS.n640 0.001007
R14022 VSS.n14092 VSS.n14090 0.001007
R14023 VSS.n1690 VSS.n1689 0.001007
R14024 VSS.n1693 VSS.n1692 0.001007
R14025 VSS.n1682 VSS.n1681 0.001007
R14026 VSS.n14102 VSS.n14101 0.001007
R14027 VSS.n14105 VSS.n14104 0.001007
R14028 VSS.n13678 VSS.n13674 0.001007
R14029 VSS.n13691 VSS.n13690 0.001007
R14030 VSS.n13683 VSS.n13682 0.001007
R14031 VSS.n1652 VSS.n1649 0.001007
R14032 VSS.n1648 VSS.n1643 0.001007
R14033 VSS.n14080 VSS.n1645 0.001007
R14034 VSS.n1667 VSS.n1647 0.001007
R14035 VSS.n14061 VSS.n1660 0.001007
R14036 VSS.n14062 VSS.n1659 0.001007
R14037 VSS.n14066 VSS.n1658 0.001007
R14038 VSS.n13666 VSS.n13665 0.001007
R14039 VSS.n13661 VSS.n13660 0.001007
R14040 VSS.n13669 VSS.n13668 0.001007
R14041 VSS.n13886 VSS.n13885 0.001007
R14042 VSS.n13892 VSS.n13891 0.001007
R14043 VSS.n13906 VSS.n13905 0.001007
R14044 VSS.n13213 VSS.n13208 0.001007
R14045 VSS.n13211 VSS.n13209 0.001007
R14046 VSS.n13632 VSS.n13234 0.001007
R14047 VSS.n13636 VSS.n13235 0.001007
R14048 VSS.n13228 VSS.n13227 0.001007
R14049 VSS.n13534 VSS.n13232 0.001007
R14050 VSS.n13544 VSS.n13231 0.001007
R14051 VSS.n13537 VSS.n13230 0.001007
R14052 VSS.n13895 VSS.n13894 0.001007
R14053 VSS.n1183 VSS.n1182 0.001007
R14054 VSS.n1187 VSS.n1175 0.001007
R14055 VSS.n1193 VSS.n1189 0.001007
R14056 VSS.n1191 VSS.n1190 0.001007
R14057 VSS.n1408 VSS.n1407 0.001007
R14058 VSS.n849 VSS.n848 0.001007
R14059 VSS.n856 VSS.n855 0.001007
R14060 VSS.n1426 VSS.n821 0.001007
R14061 VSS.n1421 VSS.n820 0.001007
R14062 VSS.n1434 VSS.n838 0.001007
R14063 VSS.n2202 VSS.n2201 0.001007
R14064 VSS.n2191 VSS.n2055 0.001007
R14065 VSS.n2199 VSS.n2198 0.001007
R14066 VSS.n2041 VSS.n1992 0.001007
R14067 VSS.n2046 VSS.n1991 0.001007
R14068 VSS.n2050 VSS.n1990 0.001007
R14069 VSS.n2008 VSS.n1989 0.001007
R14070 VSS.n2004 VSS.n1985 0.001007
R14071 VSS.n2246 VSS.n1987 0.001007
R14072 VSS.n2003 VSS.n1995 0.001007
R14073 VSS.n2231 VSS.n2230 0.001007
R14074 VSS.n2225 VSS.n2224 0.001007
R14075 VSS.n2235 VSS.n2234 0.001007
R14076 VSS.n2119 VSS.n2118 0.001007
R14077 VSS.n2106 VSS.n2104 0.001007
R14078 VSS.n2110 VSS.n2107 0.001007
R14079 VSS.n2090 VSS.n2067 0.001007
R14080 VSS.n2095 VSS.n2066 0.001007
R14081 VSS.n2099 VSS.n2065 0.001007
R14082 VSS.n2083 VSS.n2064 0.001007
R14083 VSS.n2079 VSS.n2060 0.001007
R14084 VSS.n2181 VSS.n2062 0.001007
R14085 VSS.n2078 VSS.n2070 0.001007
R14086 VSS.n2166 VSS.n2165 0.001007
R14087 VSS.n2160 VSS.n2159 0.001007
R14088 VSS.n2170 VSS.n2169 0.001007
R14089 VSS.n12665 VSS.n12664 0.001007
R14090 VSS.n12654 VSS.n12653 0.001007
R14091 VSS.n12662 VSS.n12661 0.001007
R14092 VSS.n2138 VSS.n1861 0.001007
R14093 VSS.n2141 VSS.n1860 0.001007
R14094 VSS.n2142 VSS.n1859 0.001007
R14095 VSS.n1858 VSS.n1857 0.001007
R14096 VSS.n13187 VSS.n13186 0.001007
R14097 VSS.n1870 VSS.n1865 0.001007
R14098 VSS.n1871 VSS.n1864 0.001007
R14099 VSS.n1848 VSS.n1846 0.001007
R14100 VSS.n1842 VSS.n1836 0.001007
R14101 VSS.n1834 VSS.n1833 0.001007
R14102 VSS.n1827 VSS.n1826 0.001007
R14103 VSS.n1820 VSS.n1819 0.001007
R14104 VSS.n12690 VSS.n12689 0.001007
R14105 VSS.n12684 VSS.n12683 0.001007
R14106 VSS.n12679 VSS.n12678 0.001007
R14107 VSS.n1791 VSS.n1790 0.001007
R14108 VSS.n13937 VSS.n13936 0.001007
R14109 VSS.n1793 VSS.n1779 0.001007
R14110 VSS.n1796 VSS.n1783 0.001007
R14111 VSS.n1806 VSS.n1782 0.001007
R14112 VSS.n1799 VSS.n1781 0.001007
R14113 VSS.n13921 VSS.n13920 0.001007
R14114 VSS.n2020 VSS.n2019 0.001007
R14115 VSS.n2031 VSS.n2030 0.001007
R14116 VSS.n1959 VSS.n1955 0.001007
R14117 VSS.n1966 VSS.n1965 0.001007
R14118 VSS.n2321 VSS.n2320 0.001007
R14119 VSS.n2314 VSS.n1971 0.001007
R14120 VSS.n2310 VSS.n1970 0.001007
R14121 VSS.n2305 VSS.n1969 0.001007
R14122 VSS.n2269 VSS.n2268 0.001007
R14123 VSS.n2263 VSS.n2262 0.001007
R14124 VSS.n2273 VSS.n2272 0.001007
R14125 VSS.n2648 VSS.n2571 0.001007
R14126 VSS.n2653 VSS.n2570 0.001007
R14127 VSS.n2657 VSS.n2569 0.001007
R14128 VSS.n2587 VSS.n2568 0.001007
R14129 VSS.n2583 VSS.n2564 0.001007
R14130 VSS.n12986 VSS.n2566 0.001007
R14131 VSS.n2582 VSS.n2574 0.001007
R14132 VSS.n12971 VSS.n12970 0.001007
R14133 VSS.n12975 VSS.n12974 0.001007
R14134 VSS.n2720 VSS.n2719 0.001007
R14135 VSS.n2714 VSS.n2713 0.001007
R14136 VSS.n2709 VSS.n2708 0.001007
R14137 VSS.n12965 VSS.n12964 0.001007
R14138 VSS.n2679 VSS.n2676 0.001007
R14139 VSS.n2675 VSS.n2670 0.001007
R14140 VSS.n12950 VSS.n2672 0.001007
R14141 VSS.n2694 VSS.n2674 0.001007
R14142 VSS.n12931 VSS.n2687 0.001007
R14143 VSS.n12932 VSS.n2686 0.001007
R14144 VSS.n12936 VSS.n2685 0.001007
R14145 VSS.n2784 VSS.n2783 0.001007
R14146 VSS.n2816 VSS.n2786 0.001007
R14147 VSS.n2808 VSS.n2807 0.001007
R14148 VSS.n2792 VSS.n2791 0.001007
R14149 VSS.n2800 VSS.n2799 0.001007
R14150 VSS.n2775 VSS.n2774 0.001007
R14151 VSS.n2829 VSS.n2752 0.001007
R14152 VSS.n2834 VSS.n2751 0.001007
R14153 VSS.n2838 VSS.n2750 0.001007
R14154 VSS.n2768 VSS.n2749 0.001007
R14155 VSS.n2764 VSS.n2745 0.001007
R14156 VSS.n12909 VSS.n2747 0.001007
R14157 VSS.n2763 VSS.n2755 0.001007
R14158 VSS.n12894 VSS.n12893 0.001007
R14159 VSS.n12898 VSS.n12897 0.001007
R14160 VSS.n2900 VSS.n2899 0.001007
R14161 VSS.n2894 VSS.n2893 0.001007
R14162 VSS.n2889 VSS.n2888 0.001007
R14163 VSS.n12888 VSS.n12887 0.001007
R14164 VSS.n12619 VSS.n3058 0.001007
R14165 VSS.n12632 VSS.n12631 0.001007
R14166 VSS.n12624 VSS.n12623 0.001007
R14167 VSS.n2859 VSS.n2856 0.001007
R14168 VSS.n2855 VSS.n2850 0.001007
R14169 VSS.n12873 VSS.n2852 0.001007
R14170 VSS.n2874 VSS.n2854 0.001007
R14171 VSS.n12854 VSS.n2867 0.001007
R14172 VSS.n12855 VSS.n2866 0.001007
R14173 VSS.n12859 VSS.n2865 0.001007
R14174 VSS.n3050 VSS.n3049 0.001007
R14175 VSS.n3045 VSS.n3044 0.001007
R14176 VSS.n3053 VSS.n3052 0.001007
R14177 VSS.n3032 VSS.n3031 0.001007
R14178 VSS.n3025 VSS.n3024 0.001007
R14179 VSS.n3081 VSS.n3080 0.001007
R14180 VSS.n3075 VSS.n3074 0.001007
R14181 VSS.n3070 VSS.n3069 0.001007
R14182 VSS.n2969 VSS.n2968 0.001007
R14183 VSS.n12732 VSS.n12731 0.001007
R14184 VSS.n2971 VSS.n2957 0.001007
R14185 VSS.n3001 VSS.n2961 0.001007
R14186 VSS.n3011 VSS.n2960 0.001007
R14187 VSS.n3004 VSS.n2959 0.001007
R14188 VSS.n12716 VSS.n12715 0.001007
R14189 VSS.n2600 VSS.n2599 0.001007
R14190 VSS.n2638 VSS.n2637 0.001007
R14191 VSS.n2511 VSS.n2507 0.001007
R14192 VSS.n2518 VSS.n2517 0.001007
R14193 VSS.n13026 VSS.n13025 0.001007
R14194 VSS.n13019 VSS.n2523 0.001007
R14195 VSS.n13015 VSS.n2522 0.001007
R14196 VSS.n13010 VSS.n2521 0.001007
R14197 VSS.n2624 VSS.n2623 0.001007
R14198 VSS.n2618 VSS.n2617 0.001007
R14199 VSS.n2628 VSS.n2627 0.001007
R14200 VSS.n11655 VSS.n11652 0.001007
R14201 VSS.n11649 VSS.n11646 0.001007
R14202 VSS.n11643 VSS.n11640 0.001007
R14203 VSS.n11581 VSS.n11578 0.001007
R14204 VSS.n11678 VSS.n11677 0.001007
R14205 VSS.n11673 VSS.n11670 0.001007
R14206 VSS.n11667 VSS.n11664 0.001007
R14207 VSS.n12221 VSS.n12220 0.001007
R14208 VSS.n12215 VSS.n12214 0.001007
R14209 VSS.n12260 VSS.n12259 0.001007
R14210 VSS.n12243 VSS.n12240 0.001007
R14211 VSS.n12237 VSS.n12234 0.001007
R14212 VSS.n12227 VSS.n12224 0.001007
R14213 VSS.n11724 VSS.n11721 0.001007
R14214 VSS.n11718 VSS.n11715 0.001007
R14215 VSS.n11712 VSS.n11709 0.001007
R14216 VSS.n11705 VSS.n11702 0.001007
R14217 VSS.n11747 VSS.n11746 0.001007
R14218 VSS.n11742 VSS.n11739 0.001007
R14219 VSS.n11736 VSS.n11733 0.001007
R14220 VSS.n12114 VSS.n12113 0.001007
R14221 VSS.n12108 VSS.n12107 0.001007
R14222 VSS.n12153 VSS.n12152 0.001007
R14223 VSS.n12136 VSS.n12133 0.001007
R14224 VSS.n12130 VSS.n12127 0.001007
R14225 VSS.n12120 VSS.n12117 0.001007
R14226 VSS.n12070 VSS.n12067 0.001007
R14227 VSS.n12064 VSS.n12061 0.001007
R14228 VSS.n12100 VSS.n12099 0.001007
R14229 VSS.n12058 VSS.n12055 0.001007
R14230 VSS.n12095 VSS.n12092 0.001007
R14231 VSS.n12088 VSS.n12085 0.001007
R14232 VSS.n12082 VSS.n12079 0.001007
R14233 VSS.n11946 VSS.n11945 0.001007
R14234 VSS.n11940 VSS.n11939 0.001007
R14235 VSS.n11985 VSS.n11984 0.001007
R14236 VSS.n11968 VSS.n11965 0.001007
R14237 VSS.n11962 VSS.n11959 0.001007
R14238 VSS.n11952 VSS.n11949 0.001007
R14239 VSS.n11856 VSS.n11853 0.001007
R14240 VSS.n11850 VSS.n11847 0.001007
R14241 VSS.n11844 VSS.n11841 0.001007
R14242 VSS.n11837 VSS.n11834 0.001007
R14243 VSS.n11879 VSS.n11878 0.001007
R14244 VSS.n11874 VSS.n11871 0.001007
R14245 VSS.n11868 VSS.n11865 0.001007
R14246 VSS.n3518 VSS.n3517 0.001007
R14247 VSS.n3512 VSS.n3511 0.001007
R14248 VSS.n3557 VSS.n3556 0.001007
R14249 VSS.n3540 VSS.n3537 0.001007
R14250 VSS.n3534 VSS.n3531 0.001007
R14251 VSS.n3524 VSS.n3521 0.001007
R14252 VSS.n3474 VSS.n3471 0.001007
R14253 VSS.n3468 VSS.n3465 0.001007
R14254 VSS.n3504 VSS.n3503 0.001007
R14255 VSS.n3462 VSS.n3459 0.001007
R14256 VSS.n3499 VSS.n3496 0.001007
R14257 VSS.n3492 VSS.n3489 0.001007
R14258 VSS.n3486 VSS.n3483 0.001007
R14259 VSS.n3093 VSS.n3092 0.001007
R14260 VSS.n12607 VSS.n12606 0.001007
R14261 VSS.n12592 VSS.n12589 0.001007
R14262 VSS.n3115 VSS.n3112 0.001007
R14263 VSS.n3109 VSS.n3106 0.001007
R14264 VSS.n3099 VSS.n3096 0.001007
R14265 VSS.n3151 VSS.n3150 0.001007
R14266 VSS.n3157 VSS.n3156 0.001007
R14267 VSS.n3168 VSS.n3167 0.001007
R14268 VSS.n3126 VSS.n3123 0.001007
R14269 VSS.n3132 VSS.n3129 0.001007
R14270 VSS.n3264 VSS.n3261 0.001007
R14271 VSS.n3258 VSS.n3255 0.001007
R14272 VSS.n3269 VSS.n3268 0.001007
R14273 VSS.n3227 VSS.n3224 0.001007
R14274 VSS.n3250 VSS.n3247 0.001007
R14275 VSS.n3243 VSS.n3240 0.001007
R14276 VSS.n3237 VSS.n3234 0.001007
R14277 VSS.n3163 VSS.n3160 0.001007
R14278 VSS.n11617 VSS.n11616 0.001007
R14279 VSS.n11601 VSS.n11600 0.001007
R14280 VSS.n11595 VSS.n11594 0.001007
R14281 VSS.n11589 VSS.n11588 0.001007
R14282 VSS.n11611 VSS.n11608 0.001007
R14283 VSS.n11633 VSS.n11632 0.001007
R14284 VSS.n11622 VSS.n11619 0.001007
R14285 VSS.n2980 VSS.n2979 0.001007
R14286 VSS.n2993 VSS.n2992 0.001007
R14287 VSS.n2983 VSS.n2982 0.001007
R14288 VSS.n13971 VSS.n13970 0.001007
R14289 VSS.n13984 VSS.n13983 0.001007
R14290 VSS.n13974 VSS.n13973 0.001007
R14291 VSS.n13513 VSS.n13512 0.001007
R14292 VSS.n13518 VSS.n13517 0.001007
R14293 VSS.n13525 VSS.n13524 0.001007
R14294 VSS.n13308 VSS.n13305 0.001007
R14295 VSS.n13314 VSS.n13311 0.001007
R14296 VSS.n13320 VSS.n13317 0.001007
R14297 VSS.n3284 VSS.n3283 0.001007
R14298 VSS.n3278 VSS.n3277 0.001007
R14299 VSS.n12809 VSS.n12808 0.001007
R14300 VSS.n12821 VSS.n12820 0.001007
R14301 VSS.n12807 VSS.n12805 0.00100685
R14302 VSS.n6095 VSS.n6094 0.00100593
R14303 VSS.n5913 VSS.n5912 0.00100593
R14304 VSS.n5732 VSS.n5731 0.00100593
R14305 VSS.n5552 VSS.n5551 0.00100593
R14306 VSS.n5372 VSS.n5371 0.00100593
R14307 VSS.n5192 VSS.n5191 0.00100593
R14308 VSS.n10140 VSS.n10139 0.00100593
R14309 VSS.n3701 VSS.n3700 0.00100593
R14310 VSS.n12353 VSS.n12352 0.00100593
R14311 VSS.n12270 VSS.n12269 0.00100593
R14312 VSS.n11803 VSS.n11802 0.00100593
R14313 VSS.n11820 VSS.n11819 0.00100593
R14314 VSS.n3391 VSS.n3390 0.00100593
R14315 VSS.n3337 VSS.n3336 0.00100593
R14316 VSS.n3295 VSS.n3294 0.00100593
R14317 VSS.n14507 VSS.n11 0.00100593
R14318 VSS.n4096 VSS.n4095 0.00100588
R14319 VSS.n10634 VSS.n10632 0.00100509
R14320 VSS.n10634 VSS.n10633 0.00100509
R14321 VSS.n3367 VSS.n3328 0.00100509
R14322 VSS.n3373 VSS.n3367 0.00100509
R14323 VSS.n5388 VSS.n4708 0.00100509
R14324 VSS.n5394 VSS.n5388 0.00100509
R14325 VSS.n6127 VSS.n4665 0.00100509
R14326 VSS.n6133 VSS.n6127 0.00100509
R14327 VSS.n6111 VSS.n4667 0.00100509
R14328 VSS.n6117 VSS.n6111 0.00100509
R14329 VSS.n5945 VSS.n4674 0.00100509
R14330 VSS.n5951 VSS.n5945 0.00100509
R14331 VSS.n5929 VSS.n4676 0.00100509
R14332 VSS.n5935 VSS.n5929 0.00100509
R14333 VSS.n5764 VSS.n4683 0.00100509
R14334 VSS.n5770 VSS.n5764 0.00100509
R14335 VSS.n5748 VSS.n4685 0.00100509
R14336 VSS.n5754 VSS.n5748 0.00100509
R14337 VSS.n5584 VSS.n4694 0.00100509
R14338 VSS.n5590 VSS.n5584 0.00100509
R14339 VSS.n5568 VSS.n4696 0.00100509
R14340 VSS.n5574 VSS.n5568 0.00100509
R14341 VSS.n5404 VSS.n4705 0.00100509
R14342 VSS.n5410 VSS.n5404 0.00100509
R14343 VSS.n5224 VSS.n4717 0.00100509
R14344 VSS.n5230 VSS.n5224 0.00100509
R14345 VSS.n5208 VSS.n5182 0.00100509
R14346 VSS.n5214 VSS.n5208 0.00100509
R14347 VSS.n10118 VSS.n4565 0.00100509
R14348 VSS.n10118 VSS.n10117 0.00100509
R14349 VSS.n10156 VSS.n10129 0.00100509
R14350 VSS.n10162 VSS.n10156 0.00100509
R14351 VSS.n11161 VSS.n3707 0.00100509
R14352 VSS.n11161 VSS.n11160 0.00100509
R14353 VSS.n11177 VSS.n3705 0.00100509
R14354 VSS.n11177 VSS.n11176 0.00100509
R14355 VSS.n12285 VSS.n11686 0.00100509
R14356 VSS.n12296 VSS.n12285 0.00100509
R14357 VSS.n12319 VSS.n12313 0.00100509
R14358 VSS.n11561 VSS.n11554 0.00100509
R14359 VSS.n11561 VSS.n11560 0.00100509
R14360 VSS.n3612 VSS.n3606 0.00100509
R14361 VSS.n3612 VSS.n3611 0.00100509
R14362 VSS.n12176 VSS.n12170 0.00100509
R14363 VSS.n12194 VSS.n12188 0.00100509
R14364 VSS.n14466 VSS.n14465 0.00100509
R14365 VSS.n3312 VSS.n3183 0.00100509
R14366 VSS.n3318 VSS.n3312 0.00100509
R14367 VSS.n12558 VSS.n12553 0.00100509
R14368 VSS.n12559 VSS.n12558 0.00100509
R14369 VSS.n3410 VSS.n3404 0.00100509
R14370 VSS.n3574 VSS.n3382 0.00100509
R14371 VSS.n3585 VSS.n3574 0.00100509
R14372 VSS.n11895 VSS.n11889 0.00100509
R14373 VSS.n12003 VSS.n11811 0.00100509
R14374 VSS.n12009 VSS.n12003 0.00100509
R14375 VSS.n12020 VSS.n11810 0.00100509
R14376 VSS.n12026 VSS.n12020 0.00100509
R14377 VSS.n10627 VSS.n10621 0.00100509
R14378 VSS.n10627 VSS.n10626 0.00100509
R14379 VSS.n10635 VSS.n4542 0.00100509
R14380 VSS.n3327 VSS.n3326 0.00100509
R14381 VSS.n12565 VSS.n12564 0.00100509
R14382 VSS.n3182 VSS.n3181 0.00100509
R14383 VSS.n14492 VSS.n14491 0.00100509
R14384 VSS.n11553 VSS.n11552 0.00100509
R14385 VSS.n11190 VSS.n11184 0.00100462
R14386 VSS.n705 VSS.n704 0.00100462
R14387 VSS.n693 VSS.n692 0.00100462
R14388 VSS.n13454 VSS.n13452 0.00100384
R14389 VSS.n13584 VSS.n13500 0.00100384
R14390 VSS.n1765 VSS.n1735 0.00100384
R14391 VSS.n12783 VSS.n2941 0.00100384
R14392 VSS.n4057 VSS.n4055 0.00100384
R14393 VSS.n10878 VSS.n3904 0.00100384
R14394 VSS.n10945 VSS.n10944 0.00100384
R14395 VSS.n11029 VSS.n3836 0.00100384
R14396 VSS.n9025 VSS.n9024 0.00100384
R14397 VSS.n9555 VSS.n7570 0.00100384
R14398 VSS.n8463 VSS.n8461 0.00100384
R14399 VSS.n8817 VSS.n8189 0.00100384
R14400 VSS.n7526 VSS.n7525 0.00100384
R14401 VSS.n8570 VSS.n8566 0.00100384
R14402 VSS.n8778 VSS.n8243 0.00100384
R14403 VSS.n6184 VSS.n6182 0.00100384
R14404 VSS.n6741 VSS.n6697 0.00100384
R14405 VSS.n8116 VSS.n8039 0.00100384
R14406 VSS.n8873 VSS.n7954 0.00100384
R14407 VSS.n9370 VSS.n9366 0.00100384
R14408 VSS.n7427 VSS.n7425 0.00100384
R14409 VSS.n9064 VSS.n9062 0.00100384
R14410 VSS.n9513 VSS.n8999 0.00100384
R14411 VSS.n9835 VSS.n7163 0.00100384
R14412 VSS.n7369 VSS.n7264 0.00100384
R14413 VSS.n9241 VSS.n9214 0.00100384
R14414 VSS.n8948 VSS.n7853 0.00100384
R14415 VSS.n7632 VSS.n7616 0.00100384
R14416 VSS.n7667 VSS.n7651 0.00100384
R14417 VSS.n7139 VSS.n7091 0.00100384
R14418 VSS.n8923 VSS.n7943 0.00100384
R14419 VSS.n6856 VSS.n6631 0.00100384
R14420 VSS.n6923 VSS.n6583 0.00100384
R14421 VSS.n6996 VSS.n6542 0.00100384
R14422 VSS.n7055 VSS.n6485 0.00100384
R14423 VSS.n6423 VSS.n6318 0.00100384
R14424 VSS.n6788 VSS.n6678 0.00100384
R14425 VSS.n5997 VSS.n5993 0.00100384
R14426 VSS.n5799 VSS.n5797 0.00100384
R14427 VSS.n5618 VSS.n5616 0.00100384
R14428 VSS.n5438 VSS.n5434 0.00100384
R14429 VSS.n5258 VSS.n5256 0.00100384
R14430 VSS.n3760 VSS.n3758 0.00100384
R14431 VSS.n6078 VSS.n6077 0.00100384
R14432 VSS.n11074 VSS.n11072 0.00100384
R14433 VSS.n4451 VSS.n4450 0.00100384
R14434 VSS.n4380 VSS.n4181 0.00100384
R14435 VSS.n4268 VSS.n4249 0.00100384
R14436 VSS.n659 VSS.n658 0.00100384
R14437 VSS.n1002 VSS.n998 0.00100384
R14438 VSS.n1167 VSS.n884 0.00100384
R14439 VSS.n14306 VSS.n14302 0.00100384
R14440 VSS.n2401 VSS.n555 0.00100384
R14441 VSS.n514 VSS.n513 0.00100384
R14442 VSS.n1131 VSS.n915 0.00100384
R14443 VSS.n12389 VSS.n12387 0.00100384
R14444 VSS.n13047 VSS.n2484 0.00100384
R14445 VSS.n13094 VSS.n2357 0.00100384
R14446 VSS.n2344 VSS.n1932 0.00100384
R14447 VSS.n1524 VSS.n1522 0.00100384
R14448 VSS.n13764 VSS.n13762 0.00100384
R14449 VSS.n717 VSS.n713 0.00100384
R14450 VSS.n14112 VSS.n633 0.00100384
R14451 VSS.n1662 VSS.n1646 0.00100384
R14452 VSS.n13645 VSS.n13225 0.00100384
R14453 VSS.n1411 VSS.n843 0.00100384
R14454 VSS.n2242 VSS.n1988 0.00100384
R14455 VSS.n2177 VSS.n2063 0.00100384
R14456 VSS.n13190 VSS.n1855 0.00100384
R14457 VSS.n13928 VSS.n1778 0.00100384
R14458 VSS.n1973 VSS.n1953 0.00100384
R14459 VSS.n12982 VSS.n2567 0.00100384
R14460 VSS.n2689 VSS.n2673 0.00100384
R14461 VSS.n12905 VSS.n2748 0.00100384
R14462 VSS.n2869 VSS.n2853 0.00100384
R14463 VSS.n12723 VSS.n2956 0.00100384
R14464 VSS.n2525 VSS.n2505 0.00100384
R14465 VSS.n11576 VSS.n11575 0.00100384
R14466 VSS.n11700 VSS.n11698 0.00100384
R14467 VSS.n12053 VSS.n12051 0.00100384
R14468 VSS.n11832 VSS.n11830 0.00100384
R14469 VSS.n3457 VSS.n3455 0.00100384
R14470 VSS.n3222 VSS.n3218 0.00100384
R14471 VSS.n11628 VSS.n11627 0.00100384
R14472 VSS.n10617 VSS.n10616 0.00100381
R14473 VSS.n3326 VSS.n3322 0.00100381
R14474 VSS.n5393 VSS.n5389 0.00100381
R14475 VSS.n6132 VSS.n6128 0.00100381
R14476 VSS.n6116 VSS.n6112 0.00100381
R14477 VSS.n5950 VSS.n5946 0.00100381
R14478 VSS.n5934 VSS.n5930 0.00100381
R14479 VSS.n5769 VSS.n5765 0.00100381
R14480 VSS.n5753 VSS.n5749 0.00100381
R14481 VSS.n5589 VSS.n5585 0.00100381
R14482 VSS.n5573 VSS.n5569 0.00100381
R14483 VSS.n5409 VSS.n5405 0.00100381
R14484 VSS.n5229 VSS.n5225 0.00100381
R14485 VSS.n5213 VSS.n5209 0.00100381
R14486 VSS.n10116 VSS.n10112 0.00100381
R14487 VSS.n10161 VSS.n10157 0.00100381
R14488 VSS.n11159 VSS.n11155 0.00100381
R14489 VSS.n11175 VSS.n11171 0.00100381
R14490 VSS.n12290 VSS.n12286 0.00100381
R14491 VSS.n12318 VSS.n12314 0.00100381
R14492 VSS.n11552 VSS.n11548 0.00100381
R14493 VSS.n12477 VSS.n12476 0.00100381
R14494 VSS.n12175 VSS.n12171 0.00100381
R14495 VSS.n12193 VSS.n12189 0.00100381
R14496 VSS.n14491 VSS.n14490 0.00100381
R14497 VSS.n14482 VSS.n22 0.00100381
R14498 VSS.n3181 VSS.n3177 0.00100381
R14499 VSS.n12564 VSS.n12560 0.00100381
R14500 VSS.n3409 VSS.n3405 0.00100381
R14501 VSS.n3579 VSS.n3575 0.00100381
R14502 VSS.n11894 VSS.n11890 0.00100381
R14503 VSS.n12008 VSS.n12004 0.00100381
R14504 VSS.n12025 VSS.n12021 0.00100381
R14505 VSS.n10615 VSS.n10606 0.00100381
R14506 VSS.n6102 VSS.n6101 0.0010038
R14507 VSS.n5920 VSS.n5919 0.0010038
R14508 VSS.n5739 VSS.n5738 0.0010038
R14509 VSS.n5559 VSS.n5558 0.0010038
R14510 VSS.n5379 VSS.n5378 0.0010038
R14511 VSS.n5199 VSS.n5198 0.0010038
R14512 VSS.n10147 VSS.n10146 0.0010038
R14513 VSS.n12360 VSS.n12359 0.0010038
R14514 VSS.n12276 VSS.n12275 0.0010038
R14515 VSS.n11799 VSS.n11798 0.0010038
R14516 VSS.n11816 VSS.n11815 0.0010038
R14517 VSS.n3387 VSS.n3386 0.0010038
R14518 VSS.n3333 VSS.n3332 0.0010038
R14519 VSS.n3301 VSS.n3300 0.0010038
R14520 VSS.n7 VSS.n6 0.0010038
R14521 VSS.n6103 VSS.n6102 0.00100371
R14522 VSS.n5921 VSS.n5920 0.00100371
R14523 VSS.n5740 VSS.n5739 0.00100371
R14524 VSS.n5560 VSS.n5559 0.00100371
R14525 VSS.n5380 VSS.n5379 0.00100371
R14526 VSS.n5200 VSS.n5199 0.00100371
R14527 VSS.n10148 VSS.n10147 0.00100371
R14528 VSS.n12359 VSS.n12358 0.00100371
R14529 VSS.n12277 VSS.n12276 0.00100371
R14530 VSS.n11800 VSS.n11799 0.00100371
R14531 VSS.n11817 VSS.n11816 0.00100371
R14532 VSS.n3388 VSS.n3387 0.00100371
R14533 VSS.n3334 VSS.n3333 0.00100371
R14534 VSS.n3302 VSS.n3301 0.00100371
R14535 VSS.n8 VSS.n7 0.00100371
R14536 VSS.n12478 VSS.n12477 0.00100369
R14537 VSS.n10616 VSS.n10615 0.00100369
R14538 VSS.n11338 VSS.n11337 0.00100208
R14539 VSS.n11509 VSS.n11508 0.00100208
R14540 VSS.n11196 VSS.n11195 0.00100208
R14541 VSS.n11527 VSS.n11526 0.00100116
R14542 VSS.n1507 VSS.n1506 0.00100116
R14543 VSS.n1232 VSS.n1231 0.00100116
R14544 VSS.n6144 VSS.n6143 0.00100116
R14545 VSS.n8422 VSS.n8421 0.00100116
R14546 VSS.n8643 VSS.n8642 0.00100116
R14547 VSS.n8717 VSS.n8716 0.00100116
R14548 VSS.n9718 VSS.n9717 0.00100116
R14549 VSS.n9735 VSS.n9734 0.00100116
R14550 VSS.n7487 VSS.n7486 0.00100116
R14551 VSS.n10806 VSS.n10805 0.00100116
R14552 VSS.n9763 VSS.n9762 0.00100116
R14553 VSS.n9751 VSS.n9750 0.00100116
R14554 VSS.n5961 VSS.n5960 0.00100116
R14555 VSS.n5780 VSS.n5779 0.00100116
R14556 VSS.n5599 VSS.n5598 0.00100116
R14557 VSS.n5419 VSS.n5418 0.00100116
R14558 VSS.n5239 VSS.n5238 0.00100116
R14559 VSS.n4568 VSS.n4567 0.00100116
R14560 VSS.n3710 VSS.n3709 0.00100116
R14561 VSS.n11517 VSS.n11516 0.00100116
R14562 VSS.n10731 VSS.n10730 0.00100116
R14563 VSS.n10721 VSS.n10720 0.00100116
R14564 VSS.n986 VSS.n985 0.00100116
R14565 VSS.n14351 VSS.n14350 0.00100116
R14566 VSS.n503 VSS.n502 0.00100116
R14567 VSS.n1066 VSS.n1065 0.00100116
R14568 VSS.n1317 VSS.n1316 0.00100116
R14569 VSS.n459 VSS.n458 0.00100116
R14570 VSS.n13745 VSS.n13744 0.00100116
R14571 VSS.n13282 VSS.n13281 0.00100116
R14572 VSS.n13351 VSS.n13350 0.00100116
R14573 VSS.n13828 VSS.n13827 0.00100116
R14574 VSS.n1588 VSS.n1587 0.00100116
R14575 VSS.n12329 VSS.n12328 0.00100116
R14576 VSS.n11755 VSS.n11754 0.00100116
R14577 VSS.n12035 VSS.n12034 0.00100116
R14578 VSS.n11918 VSS.n11917 0.00100116
R14579 VSS.n3437 VSS.n3436 0.00100116
R14580 VSS.n12572 VSS.n12571 0.00100116
R14581 VSS.n13412 VSS.n13411 0.00100116
R14582 VSS.n4478 VSS.n4477 0.00100062
R14583 VSS.n4500 VSS.n4499 0.00100062
R14584 VSS.n3699 VSS.n3698 0.0010004
R14585 VSS.n3697 VSS.n3696 0.0010004
R14586 VSS.n14504 VSS.n19 0.00100037
R14587 VSS.n14479 VSS.n14478 0.00100037
R14588 VSS.n505 VSS.n504 0.00100034
R14589 VSS.n1234 VSS.n1233 0.00100034
R14590 VSS.n13747 VSS.n13746 0.00100034
R14591 VSS.n13284 VSS.n13283 0.00100034
R14592 VSS.n13414 VSS.n13413 0.00100034
R14593 VSS.n4526 VSS.n4525 0.00100033
R14594 VSS.n4467 VSS.n4466 0.00100031
R14595 VSS.n4514 VSS.n4513 0.00100031
R14596 VSS.n382 VSS.n381 0.00100031
R14597 VSS.n37 VSS.n36 0.00100031
R14598 VSS.n180 VSS.n179 0.00100031
R14599 VSS.n344 VSS.n343 0.00100031
R14600 VSS.n271 VSS.n270 0.00100031
R14601 VSS.n159 VSS.n158 0.00100031
R14602 VSS.n98 VSS.n97 0.00100031
R14603 VSS.n11524 VSS.n11522 0.00100024
R14604 VSS.n5601 VSS.n5597 0.00100022
R14605 VSS.n5421 VSS.n5417 0.00100022
R14606 VSS.n5241 VSS.n5237 0.00100022
R14607 VSS.n10106 VSS.n10104 0.00100022
R14608 VSS.n11149 VSS.n11147 0.00100022
R14609 VSS.n9757 VSS.n7489 0.00100021
R14610 VSS.n988 VSS.n984 0.00100021
R14611 VSS.n1509 VSS.n1505 0.00100021
R14612 VSS.n457 VSS.n456 0.00100021
R14613 VSS.n702 VSS.n701 0.00100021
R14614 VSS.n3297 VSS.n3184 0.00100021
R14615 VSS.n3354 VSS.n3339 0.00100021
R14616 VSS.n3394 VSS.n3393 0.00100021
R14617 VSS.n11823 VSS.n11822 0.00100021
R14618 VSS.n11806 VSS.n11805 0.00100021
R14619 VSS.n12272 VSS.n11689 0.00100021
R14620 VSS.n12355 VSS.n12351 0.00100021
R14621 VSS.n12038 VSS.n12037 0.00100021
R14622 VSS.n11925 VSS.n11924 0.00100021
R14623 VSS.n3440 VSS.n3439 0.00100021
R14624 VSS.n11288 VSS.n11287 0.00100018
R14625 VSS.n301 VSS.n300 0.00100018
R14626 VSS.n6242 VSS.n6237 0.00100017
R14627 VSS.n8844 VSS.n8843 0.00100017
R14628 VSS.n9540 VSS.n7594 0.00100017
R14629 VSS.n9852 VSS.n9851 0.00100017
R14630 VSS.n9859 VSS.n9856 0.00100017
R14631 VSS.n9851 VSS.n9850 0.00100017
R14632 VSS.n7605 VSS.n7604 0.00100017
R14633 VSS.n9532 VSS.n9531 0.00100017
R14634 VSS.n9920 VSS.n9919 0.00100017
R14635 VSS.n9912 VSS.n9911 0.00100017
R14636 VSS.n9906 VSS.n6268 0.00100017
R14637 VSS.n9912 VSS.n6261 0.00100017
R14638 VSS.n9920 VSS.n6256 0.00100017
R14639 VSS.n9928 VSS.n9927 0.00100017
R14640 VSS.n6249 VSS.n6248 0.00100017
R14641 VSS.n10036 VSS.n10033 0.00100017
R14642 VSS.n4638 VSS.n4637 0.00100017
R14643 VSS.n10022 VSS.n10021 0.00100017
R14644 VSS.n10013 VSS.n10012 0.00100017
R14645 VSS.n10004 VSS.n10003 0.00100017
R14646 VSS.n9995 VSS.n9994 0.00100017
R14647 VSS.n3783 VSS.n3782 0.00100017
R14648 VSS.n11115 VSS.n3822 0.00100017
R14649 VSS.n11117 VSS.n3822 0.00100017
R14650 VSS.n11119 VSS.n3819 0.00100017
R14651 VSS.n11121 VSS.n3819 0.00100017
R14652 VSS.n11006 VSS.n3841 0.00100017
R14653 VSS.n11004 VSS.n3841 0.00100017
R14654 VSS.n11001 VSS.n11000 0.00100017
R14655 VSS.n11000 VSS.n10999 0.00100017
R14656 VSS.n10956 VSS.n3890 0.00100017
R14657 VSS.n10958 VSS.n3890 0.00100017
R14658 VSS.n10960 VSS.n3887 0.00100017
R14659 VSS.n10962 VSS.n3887 0.00100017
R14660 VSS.n4439 VSS.n4154 0.00100017
R14661 VSS.n4352 VSS.n4207 0.00100017
R14662 VSS.n13146 VSS.n13145 0.00100017
R14663 VSS.n14149 VSS.n14148 0.00100017
R14664 VSS.n14140 VSS.n14139 0.00100017
R14665 VSS.n14053 VSS.n14044 0.00100017
R14666 VSS.n14039 VSS.n1705 0.00100017
R14667 VSS.n14053 VSS.n14052 0.00100017
R14668 VSS.n14047 VSS.n14046 0.00100017
R14669 VSS.n14131 VSS.n14130 0.00100017
R14670 VSS.n13176 VSS.n1887 0.00100017
R14671 VSS.n12703 VSS.n12700 0.00100017
R14672 VSS.n13176 VSS.n13175 0.00100017
R14673 VSS.n1890 VSS.n1889 0.00100017
R14674 VSS.n13164 VSS.n13163 0.00100017
R14675 VSS.n13155 VSS.n13154 0.00100017
R14676 VSS.n12840 VSS.n2920 0.00100017
R14677 VSS.n12845 VSS.n2915 0.00100017
R14678 VSS.n2911 VSS.n2910 0.00100017
R14679 VSS.n12922 VSS.n2735 0.00100017
R14680 VSS.n2731 VSS.n2730 0.00100017
R14681 VSS.n2555 VSS.n2554 0.00100017
R14682 VSS.n12826 VSS.n2927 0.00100017
R14683 VSS.n12828 VSS.n2927 0.00100017
R14684 VSS.n12832 VSS.n12830 0.00100017
R14685 VSS.n12832 VSS.n12831 0.00100017
R14686 VSS.n14002 VSS.n1748 0.00100017
R14687 VSS.n14000 VSS.n1748 0.00100017
R14688 VSS.n13997 VSS.n13996 0.00100017
R14689 VSS.n13996 VSS.n13995 0.00100017
R14690 VSS.n14025 VSS.n1712 0.00100017
R14691 VSS.n14027 VSS.n1712 0.00100017
R14692 VSS.n14031 VSS.n14029 0.00100017
R14693 VSS.n14031 VSS.n14030 0.00100017
R14694 VSS.n6086 VSS.n6085 0.00100017
R14695 VSS.n5904 VSS.n5903 0.00100017
R14696 VSS.n5723 VSS.n5722 0.00100017
R14697 VSS.n5543 VSS.n5542 0.00100017
R14698 VSS.n5363 VSS.n5362 0.00100017
R14699 VSS.n10097 VSS.n10096 0.00100017
R14700 VSS.n10744 VSS.n10743 0.00100017
R14701 VSS.n14370 VSS.n14369 0.00100017
R14702 VSS.n1245 VSS.n1244 0.00100017
R14703 VSS.n13426 VSS.n13425 0.00100017
R14704 VSS.n9941 VSS.n6242 0.00100017
R14705 VSS.n8843 VSS.n8842 0.00100017
R14706 VSS.n7595 VSS.n7594 0.00100017
R14707 VSS.n9601 VSS.n9600 0.00100017
R14708 VSS.n8766 VSS.n8765 0.00100017
R14709 VSS.n8523 VSS.n8522 0.00100017
R14710 VSS.n9797 VSS.n9796 0.00100017
R14711 VSS.n9463 VSS.n9462 0.00100017
R14712 VSS.n9154 VSS.n9153 0.00100017
R14713 VSS.n9857 VSS.n9856 0.00100017
R14714 VSS.n7604 VSS.n7602 0.00100017
R14715 VSS.n9533 VSS.n9532 0.00100017
R14716 VSS.n9904 VSS.n6268 0.00100017
R14717 VSS.n9927 VSS.n6254 0.00100017
R14718 VSS.n9935 VSS.n6249 0.00100017
R14719 VSS.n10034 VSS.n10033 0.00100017
R14720 VSS.n10030 VSS.n4638 0.00100017
R14721 VSS.n10021 VSS.n4642 0.00100017
R14722 VSS.n10012 VSS.n4646 0.00100017
R14723 VSS.n10003 VSS.n4650 0.00100017
R14724 VSS.n9994 VSS.n4654 0.00100017
R14725 VSS.n4155 VSS.n4154 0.00100017
R14726 VSS.n4226 VSS.n4207 0.00100017
R14727 VSS.n540 VSS.n539 0.00100017
R14728 VSS.n13145 VSS.n1902 0.00100017
R14729 VSS.n14148 VSS.n14147 0.00100017
R14730 VSS.n14139 VSS.n618 0.00100017
R14731 VSS.n1357 VSS.n1356 0.00100017
R14732 VSS.n1125 VSS.n1124 0.00100017
R14733 VSS.n13865 VSS.n13864 0.00100017
R14734 VSS.n1627 VSS.n1626 0.00100017
R14735 VSS.n807 VSS.n806 0.00100017
R14736 VSS.n1707 VSS.n1705 0.00100017
R14737 VSS.n14049 VSS.n14047 0.00100017
R14738 VSS.n14132 VSS.n14131 0.00100017
R14739 VSS.n12701 VSS.n12700 0.00100017
R14740 VSS.n13172 VSS.n1890 0.00100017
R14741 VSS.n13163 VSS.n1894 0.00100017
R14742 VSS.n13154 VSS.n1898 0.00100017
R14743 VSS.n2922 VSS.n2920 0.00100017
R14744 VSS.n2916 VSS.n2915 0.00100017
R14745 VSS.n2910 VSS.n2908 0.00100017
R14746 VSS.n2736 VSS.n2735 0.00100017
R14747 VSS.n2730 VSS.n2728 0.00100017
R14748 VSS.n12999 VSS.n2555 0.00100017
R14749 VSS.n12819 VSS.n12807 0.00100016
R14750 VSS.n12819 VSS.n12818 0.00100015
R14751 VSS.n6154 VSS.n6153 0.00100011
R14752 VSS.n4326 VSS.n4325 0.00100011
R14753 VSS.n12460 VSS.n12459 0.00100011
R14754 VSS.n9429 VSS.n9363 0.00100011
R14755 VSS.n1601 VSS.n1517 0.00100011
R14756 VSS.n14356 VSS.n14355 0.0010001
R14757 VSS.n467 VSS.n466 0.0010001
R14758 VSS.n698 VSS.n689 0.0010001
R14759 VSS.n1320 VSS.n1315 0.0010001
R14760 VSS.n11775 VSS.n11758 0.0010001
R14761 VSS.n11923 VSS.n11922 0.0010001
R14762 VSS.n3433 VSS.n3432 0.0010001
R14763 VSS.n15 VSS.n14 0.00100009
R14764 VSS.n8631 VSS.n8630 0.00100009
R14765 VSS.n8630 VSS.n8629 0.00100009
R14766 VSS.n8732 VSS.n8731 0.00100009
R14767 VSS.n8732 VSS.n8320 0.00100009
R14768 VSS.n9706 VSS.n9705 0.00100009
R14769 VSS.n9705 VSS.n9704 0.00100009
R14770 VSS.n9119 VSS.n9118 0.00100009
R14771 VSS.n9119 VSS.n9053 0.00100009
R14772 VSS.n10821 VSS.n10820 0.00100009
R14773 VSS.n10821 VSS.n3955 0.00100009
R14774 VSS.n9774 VSS.n9773 0.00100009
R14775 VSS.n9774 VSS.n7420 0.00100009
R14776 VSS.n11081 VSS.n11080 0.00100009
R14777 VSS.n14366 VSS.n14365 0.00100009
R14778 VSS.n14366 VSS.n14364 0.00100009
R14779 VSS.n1080 VSS.n1079 0.00100009
R14780 VSS.n1080 VSS.n1078 0.00100009
R14781 VSS.n1330 VSS.n1329 0.00100009
R14782 VSS.n1330 VSS.n1328 0.00100009
R14783 VSS.n772 VSS.n771 0.00100009
R14784 VSS.n772 VSS.n687 0.00100009
R14785 VSS.n13377 VSS.n13376 0.00100009
R14786 VSS.n13377 VSS.n13375 0.00100009
R14787 VSS.n13842 VSS.n13841 0.00100009
R14788 VSS.n13842 VSS.n13840 0.00100009
R14789 VSS.n12341 VSS.n12340 0.00100009
R14790 VSS.n12208 VSS.n12207 0.00100009
R14791 VSS.n12044 VSS.n12043 0.00100009
R14792 VSS.n11933 VSS.n11932 0.00100009
R14793 VSS.n3448 VSS.n3447 0.00100009
R14794 VSS.n12583 VSS.n12582 0.00100009
R14795 VSS.n12814 VSS.n12813 0.00100009
R14796 VSS.n3288 VSS.n3189 0.00100009
R14797 VSS.n10810 VSS.n10809 0.00100008
R14798 VSS.n3966 VSS.n3965 0.00100008
R14799 VSS.n9760 VSS.n9759 0.00100008
R14800 VSS.n9749 VSS.n9748 0.00100008
R14801 VSS.n9741 VSS.n9740 0.00100008
R14802 VSS.n9733 VSS.n9732 0.00100008
R14803 VSS.n9724 VSS.n9723 0.00100008
R14804 VSS.n9716 VSS.n9715 0.00100008
R14805 VSS.n7515 VSS.n7514 0.00100008
R14806 VSS.n8721 VSS.n8720 0.00100008
R14807 VSS.n8649 VSS.n8648 0.00100008
R14808 VSS.n8641 VSS.n8640 0.00100008
R14809 VSS.n8338 VSS.n8337 0.00100008
R14810 VSS.n13364 VSS.n13363 0.00100008
R14811 VSS.n12576 VSS.n12575 0.00100008
R14812 VSS.n7482 VSS.n7481 0.00100007
R14813 VSS.n9430 VSS.n9429 0.00100007
R14814 VSS.n1602 VSS.n1601 0.00100007
R14815 VSS.n13743 VSS.n13742 0.00100006
R14816 VSS.n6098 VSS.n6097 0.00100006
R14817 VSS.n5916 VSS.n5915 0.00100006
R14818 VSS.n5735 VSS.n5734 0.00100006
R14819 VSS.n5555 VSS.n5554 0.00100006
R14820 VSS.n5375 VSS.n5374 0.00100006
R14821 VSS.n5195 VSS.n5194 0.00100006
R14822 VSS.n10143 VSS.n10142 0.00100006
R14823 VSS.n11192 VSS.n3703 0.00100006
R14824 VSS.n6146 VSS.n6142 0.00100006
R14825 VSS.n5963 VSS.n5959 0.00100006
R14826 VSS.n5782 VSS.n5778 0.00100006
R14827 VSS.n18 VSS.n16 0.00100006
R14828 VSS.n1515 VSS.n1514 0.00100006
R14829 VSS.n13293 VSS.n13279 0.00100006
R14830 VSS.n13756 VSS.n13755 0.00100006
R14831 VSS.n994 VSS.n993 0.00100006
R14832 VSS.n10725 VSS.n10723 0.00100006
R14833 VSS.n8424 VSS.n8420 0.00100006
R14834 VSS.n10802 VSS.n4098 0.00100006
R14835 VSS.n11329 VSS.n11194 0.00100006
R14836 VSS.n11336 VSS.n11333 0.00100006
R14837 VSS.n13366 VSS.n13365 0.00100005
R14838 VSS.n3175 VSS.n3174 0.00100005
R14839 VSS.n11500 VSS.n11490 0.00100002
R14840 VSS.n11501 VSS.n3630 0.00100001
R14841 VSS.n8334 VSS.n8333 0.001
R14842 VSS.n8327 VSS.n8326 0.001
R14843 VSS.n7511 VSS.n7510 0.001
R14844 VSS.n7504 VSS.n7503 0.001
R14845 VSS.n3962 VSS.n3961 0.001
R14846 VSS.n3328 VSS.n3327 0.001
R14847 VSS.n4665 VSS.n4664 0.001
R14848 VSS.n11686 VSS.n11685 0.001
R14849 VSS.n12321 VSS.n12320 0.001
R14850 VSS.n11554 VSS.n11553 0.001
R14851 VSS.n12178 VSS.n12177 0.001
R14852 VSS.n12196 VSS.n12195 0.001
R14853 VSS.n14492 VSS.n14489 0.001
R14854 VSS.n14465 VSS.n14464 0.001
R14855 VSS.n3183 VSS.n3182 0.001
R14856 VSS.n3412 VSS.n3411 0.001
R14857 VSS.n3382 VSS.n3381 0.001
R14858 VSS.n11897 VSS.n11896 0.001
R14859 VSS.n11810 VSS.n11809 0.001
R14860 VSS.n9744 VSS.n9743 0.001
R14861 VSS.n694 VSS.n693 0.001
R14862 VSS.n12819 VSS.n12809 0.001
R14863 VSS.n12820 VSS.n12819 0.001
R14864 VSS.n14509 VSS.n14508 0.001
R14865 VSS.n3194 VSS.n3193 0.001
R14866 VSS.n706 VSS.n705 0.001
R14867 VSS.n10607 VSS.n4542 0.001
R14868 VSS.n4090 VSS.n4032 0.001
R14869 VSS.n7502 VSS.n7501 0.001
R14870 VSS.n10628 VSS.n10627 0.001
R14871 VSS.n3284 VSS.n3282 0.001
R14872 VSS.n3282 VSS.n3278 0.001
R14873 VSS.n9690 VSS.n9682 0.001
R14874 VSS.n9137 VSS.n9052 0.001
R14875 VSS.n8557 VSS.n8351 0.001
R14876 VSS.n8702 VSS.n8694 0.001
R14877 VSS.n9634 VSS.n9624 0.001
R14878 VSS.n8747 VSS.n8305 0.001
R14879 VSS.n8249 VSS.n8215 0.001
R14880 VSS.n6203 VSS.n6193 0.001
R14881 VSS.n9957 VSS.n6230 0.001
R14882 VSS.n8853 VSS.n7953 0.001
R14883 VSS.n8482 VSS.n8449 0.001
R14884 VSS.n9444 VSS.n9339 0.001
R14885 VSS.n9815 VSS.n7180 0.001
R14886 VSS.n7367 VSS.n7272 0.001
R14887 VSS.n7208 VSS.n7194 0.001
R14888 VSS.n9265 VSS.n9169 0.001
R14889 VSS.n8958 VSS.n7815 0.001
R14890 VSS.n7788 VSS.n7631 0.001
R14891 VSS.n7709 VSS.n7666 0.001
R14892 VSS.n7137 VSS.n7116 0.001
R14893 VSS.n9872 VSS.n7087 0.001
R14894 VSS.n8932 VSS.n7888 0.001
R14895 VSS.n7984 VSS.n7877 0.001
R14896 VSS.n6887 VSS.n6626 0.001
R14897 VSS.n6960 VSS.n6578 0.001
R14898 VSS.n7040 VSS.n6517 0.001
R14899 VSS.n6289 VSS.n6275 0.001
R14900 VSS.n6421 VSS.n6326 0.001
R14901 VSS.n6434 VSS.n6314 0.001
R14902 VSS.n6820 VSS.n6674 0.001
R14903 VSS.n6786 VSS.n6680 0.001
R14904 VSS.n5895 VSS.n5894 0.001
R14905 VSS.n5714 VSS.n5713 0.001
R14906 VSS.n5534 VSS.n5533 0.001
R14907 VSS.n5354 VSS.n5353 0.001
R14908 VSS.n10088 VSS.n10087 0.001
R14909 VSS.n3809 VSS.n3796 0.001
R14910 VSS.n4624 VSS.n4611 0.001
R14911 VSS.n6079 VSS.n5990 0.001
R14912 VSS.n11134 VSS.n3741 0.001
R14913 VSS.n11107 VSS.n11060 0.001
R14914 VSS.n6337 VSS.n3830 0.001
R14915 VSS.n11042 VSS.n3833 0.001
R14916 VSS.n10987 VSS.n3873 0.001
R14917 VSS.n10906 VSS.n3859 0.001
R14918 VSS.n7283 VSS.n3898 0.001
R14919 VSS.n10891 VSS.n3901 0.001
R14920 VSS.n4019 VSS.n4001 0.001
R14921 VSS.n4083 VSS.n4043 0.001
R14922 VSS.n4404 VSS.n4190 0.001
R14923 VSS.n4283 VSS.n4234 0.001
R14924 VSS.n4344 VSS.n4236 0.001
R14925 VSS.n10776 VSS.n4119 0.001
R14926 VSS.n10754 VSS.n4114 0.001
R14927 VSS.n1296 VSS.n1288 0.001
R14928 VSS.n790 VSS.n686 0.001
R14929 VSS.n1345 VSS.n1216 0.001
R14930 VSS.n1106 VSS.n964 0.001
R14931 VSS.n14228 VSS.n572 0.001
R14932 VSS.n14229 VSS.n556 0.001
R14933 VSS.n14275 VSS.n14265 0.001
R14934 VSS.n13045 VSS.n2492 0.001
R14935 VSS.n2478 VSS.n2465 0.001
R14936 VSS.n13101 VSS.n2364 0.001
R14937 VSS.n13113 VSS.n1928 0.001
R14938 VSS.n1616 VSS.n1485 0.001
R14939 VSS.n13658 VSS.n1661 0.001
R14940 VSS.n13643 VSS.n13233 0.001
R14941 VSS.n13883 VSS.n13221 0.001
R14942 VSS.n1435 VSS.n822 0.001
R14943 VSS.n2222 VSS.n2005 0.001
R14944 VSS.n2157 VSS.n2080 0.001
R14945 VSS.n1849 VSS.n1835 0.001
R14946 VSS.n13935 VSS.n1785 0.001
R14947 VSS.n1823 VSS.n1777 0.001
R14948 VSS.n2017 VSS.n1972 0.001
R14949 VSS.n2319 VSS.n1954 0.001
R14950 VSS.n12962 VSS.n2584 0.001
R14951 VSS.n2777 VSS.n2688 0.001
R14952 VSS.n12885 VSS.n2765 0.001
R14953 VSS.n3042 VSS.n2868 0.001
R14954 VSS.n12730 VSS.n2963 0.001
R14955 VSS.n3028 VSS.n2955 0.001
R14956 VSS.n2597 VSS.n2524 0.001
R14957 VSS.n13024 VSS.n2506 0.001
R14958 VSS.n12256 VSS.n12255 0.001
R14959 VSS.n12149 VSS.n12148 0.001
R14960 VSS.n11981 VSS.n11980 0.001
R14961 VSS.n3553 VSS.n3552 0.001
R14962 VSS.n12605 VSS.n12604 0.001
R14963 VSS.n3164 VSS.n3145 0.001
R14964 VSS.n11629 VSS.n11605 0.001
R14965 VSS.n12739 VSS.n2935 0.001
R14966 VSS.n12796 VSS.n2938 0.001
R14967 VSS.n13948 VSS.n1720 0.001
R14968 VSS.n14016 VSS.n1722 0.001
R14969 VSS.n13564 VSS.n13485 0.001
R14970 VSS.n13603 VSS.n13487 0.001
R14971 VSS.n13344 VSS.n13328 0.001
R14972 VSS.n13473 VSS.n13440 0.001
R14973 VSS.n13473 VSS.n13472 0.001
R14974 VSS.n13473 VSS.n13466 0.001
R14975 VSS.n13473 VSS.n13460 0.001
R14976 VSS.n13474 VSS.n13473 0.001
R14977 VSS.n13603 VSS.n13602 0.001
R14978 VSS.n13603 VSS.n13504 0.001
R14979 VSS.n13603 VSS.n13503 0.001
R14980 VSS.n13603 VSS.n13501 0.001
R14981 VSS.n14016 VSS.n14015 0.001
R14982 VSS.n14016 VSS.n1739 0.001
R14983 VSS.n14016 VSS.n1738 0.001
R14984 VSS.n14016 VSS.n1736 0.001
R14985 VSS.n12797 VSS.n12796 0.001
R14986 VSS.n12796 VSS.n12795 0.001
R14987 VSS.n12796 VSS.n12786 0.001
R14988 VSS.n12796 VSS.n2942 0.001
R14989 VSS.n4083 VSS.n4082 0.001
R14990 VSS.n4083 VSS.n4076 0.001
R14991 VSS.n4083 VSS.n4070 0.001
R14992 VSS.n4083 VSS.n4064 0.001
R14993 VSS.n10892 VSS.n10891 0.001
R14994 VSS.n10891 VSS.n10890 0.001
R14995 VSS.n10891 VSS.n10881 0.001
R14996 VSS.n10891 VSS.n3905 0.001
R14997 VSS.n10937 VSS.n3859 0.001
R14998 VSS.n10934 VSS.n3859 0.001
R14999 VSS.n10929 VSS.n3859 0.001
R15000 VSS.n10922 VSS.n3859 0.001
R15001 VSS.n11043 VSS.n11042 0.001
R15002 VSS.n11042 VSS.n11041 0.001
R15003 VSS.n11042 VSS.n11032 0.001
R15004 VSS.n11042 VSS.n3837 0.001
R15005 VSS.n9690 VSS.n9678 0.001
R15006 VSS.n9690 VSS.n9672 0.001
R15007 VSS.n9691 VSS.n9690 0.001
R15008 VSS.n9137 VSS.n9133 0.001
R15009 VSS.n9137 VSS.n9127 0.001
R15010 VSS.n9138 VSS.n9137 0.001
R15011 VSS.n9137 VSS.n9046 0.001
R15012 VSS.n9137 VSS.n9040 0.001
R15013 VSS.n9137 VSS.n9034 0.001
R15014 VSS.n9137 VSS.n9030 0.001
R15015 VSS.n9690 VSS.n9689 0.001
R15016 VSS.n9690 VSS.n9658 0.001
R15017 VSS.n9690 VSS.n9652 0.001
R15018 VSS.n9690 VSS.n9646 0.001
R15019 VSS.n8557 VSS.n8357 0.001
R15020 VSS.n8557 VSS.n8363 0.001
R15021 VSS.n8558 VSS.n8557 0.001
R15022 VSS.n8482 VSS.n8478 0.001
R15023 VSS.n8482 VSS.n8472 0.001
R15024 VSS.n8482 VSS.n8468 0.001
R15025 VSS.n8483 VSS.n8482 0.001
R15026 VSS.n8826 VSS.n8182 0.001
R15027 VSS.n8826 VSS.n8181 0.001
R15028 VSS.n8826 VSS.n8180 0.001
R15029 VSS.n8826 VSS.n8179 0.001
R15030 VSS.n8375 VSS.n8183 0.001
R15031 VSS.n8368 VSS.n8183 0.001
R15032 VSS.n8382 VSS.n8183 0.001
R15033 VSS.n8788 VSS.n8214 0.001
R15034 VSS.n8788 VSS.n8213 0.001
R15035 VSS.n8788 VSS.n8212 0.001
R15036 VSS.n8788 VSS.n8211 0.001
R15037 VSS.n8702 VSS.n8690 0.001
R15038 VSS.n8702 VSS.n8684 0.001
R15039 VSS.n8703 VSS.n8702 0.001
R15040 VSS.n9634 VSS.n9630 0.001
R15041 VSS.n9635 VSS.n9634 0.001
R15042 VSS.n9634 VSS.n9618 0.001
R15043 VSS.n9634 VSS.n7547 0.001
R15044 VSS.n9634 VSS.n7541 0.001
R15045 VSS.n9634 VSS.n7535 0.001
R15046 VSS.n9634 VSS.n7531 0.001
R15047 VSS.n8702 VSS.n8701 0.001
R15048 VSS.n8702 VSS.n8670 0.001
R15049 VSS.n8702 VSS.n8664 0.001
R15050 VSS.n8702 VSS.n8658 0.001
R15051 VSS.n8747 VSS.n8311 0.001
R15052 VSS.n8747 VSS.n8317 0.001
R15053 VSS.n8747 VSS.n8738 0.001
R15054 VSS.n8615 VSS.n8612 0.001
R15055 VSS.n8615 VSS.n8605 0.001
R15056 VSS.n8615 VSS.n8599 0.001
R15057 VSS.n8615 VSS.n8593 0.001
R15058 VSS.n8615 VSS.n8587 0.001
R15059 VSS.n8615 VSS.n8581 0.001
R15060 VSS.n8616 VSS.n8615 0.001
R15061 VSS.n8615 VSS.n8575 0.001
R15062 VSS.n8750 VSS.n8747 0.001
R15063 VSS.n8747 VSS.n8301 0.001
R15064 VSS.n8747 VSS.n8295 0.001
R15065 VSS.n8747 VSS.n8289 0.001
R15066 VSS.n8255 VSS.n8215 0.001
R15067 VSS.n8256 VSS.n8215 0.001
R15068 VSS.n8240 VSS.n8215 0.001
R15069 VSS.n8224 VSS.n8215 0.001
R15070 VSS.n8232 VSS.n8215 0.001
R15071 VSS.n8227 VSS.n8215 0.001
R15072 VSS.n8776 VSS.n8215 0.001
R15073 VSS.n8788 VSS.n8787 0.001
R15074 VSS.n8789 VSS.n8788 0.001
R15075 VSS.n8788 VSS.n8208 0.001
R15076 VSS.n8788 VSS.n8199 0.001
R15077 VSS.n6203 VSS.n6199 0.001
R15078 VSS.n6203 VSS.n6189 0.001
R15079 VSS.n6204 VSS.n6203 0.001
R15080 VSS.n9979 VSS.n6230 0.001
R15081 VSS.n6230 VSS.n6217 0.001
R15082 VSS.n6230 VSS.n6218 0.001
R15083 VSS.n6230 VSS.n6229 0.001
R15084 VSS.n6761 VSS.n6714 0.001
R15085 VSS.n6761 VSS.n6713 0.001
R15086 VSS.n6761 VSS.n6712 0.001
R15087 VSS.n6761 VSS.n6695 0.001
R15088 VSS.n6762 VSS.n6761 0.001
R15089 VSS.n6761 VSS.n6709 0.001
R15090 VSS.n6761 VSS.n6699 0.001
R15091 VSS.n6761 VSS.n6698 0.001
R15092 VSS.n9968 VSS.n6230 0.001
R15093 VSS.n9966 VSS.n6230 0.001
R15094 VSS.n9959 VSS.n6230 0.001
R15095 VSS.n8152 VSS.n8034 0.001
R15096 VSS.n8034 VSS.n8019 0.001
R15097 VSS.n8034 VSS.n8033 0.001
R15098 VSS.n8034 VSS.n8021 0.001
R15099 VSS.n8114 VSS.n8094 0.001
R15100 VSS.n8114 VSS.n8093 0.001
R15101 VSS.n8114 VSS.n8092 0.001
R15102 VSS.n8114 VSS.n8091 0.001
R15103 VSS.n8114 VSS.n8045 0.001
R15104 VSS.n8114 VSS.n8044 0.001
R15105 VSS.n8114 VSS.n8043 0.001
R15106 VSS.n8114 VSS.n8042 0.001
R15107 VSS.n8127 VSS.n8034 0.001
R15108 VSS.n8142 VSS.n8034 0.001
R15109 VSS.n8130 VSS.n8034 0.001
R15110 VSS.n8135 VSS.n8034 0.001
R15111 VSS.n8070 VSS.n7953 0.001
R15112 VSS.n8065 VSS.n7953 0.001
R15113 VSS.n8059 VSS.n7953 0.001
R15114 VSS.n8057 VSS.n7953 0.001
R15115 VSS.n8893 VSS.n7971 0.001
R15116 VSS.n8893 VSS.n7970 0.001
R15117 VSS.n8893 VSS.n7969 0.001
R15118 VSS.n8893 VSS.n7951 0.001
R15119 VSS.n8894 VSS.n8893 0.001
R15120 VSS.n8893 VSS.n7966 0.001
R15121 VSS.n8893 VSS.n7956 0.001
R15122 VSS.n8893 VSS.n7955 0.001
R15123 VSS.n8866 VSS.n7953 0.001
R15124 VSS.n8860 VSS.n7953 0.001
R15125 VSS.n8858 VSS.n7953 0.001
R15126 VSS.n8814 VSS.n8183 0.001
R15127 VSS.n8798 VSS.n8183 0.001
R15128 VSS.n8805 VSS.n8183 0.001
R15129 VSS.n8800 VSS.n8183 0.001
R15130 VSS.n8384 VSS.n8183 0.001
R15131 VSS.n8826 VSS.n8825 0.001
R15132 VSS.n8827 VSS.n8826 0.001
R15133 VSS.n8826 VSS.n8176 0.001
R15134 VSS.n8826 VSS.n8167 0.001
R15135 VSS.n9552 VSS.n7555 0.001
R15136 VSS.n7575 VSS.n7555 0.001
R15137 VSS.n7583 VSS.n7555 0.001
R15138 VSS.n7580 VSS.n7555 0.001
R15139 VSS.n8271 VSS.n7555 0.001
R15140 VSS.n8264 VSS.n7555 0.001
R15141 VSS.n8278 VSS.n7555 0.001
R15142 VSS.n8280 VSS.n7555 0.001
R15143 VSS.n9577 VSS.n7559 0.001
R15144 VSS.n9577 VSS.n7560 0.001
R15145 VSS.n9577 VSS.n7561 0.001
R15146 VSS.n9577 VSS.n9576 0.001
R15147 VSS.n9581 VSS.n9577 0.001
R15148 VSS.n9589 VSS.n9577 0.001
R15149 VSS.n9592 VSS.n9577 0.001
R15150 VSS.n8557 VSS.n8535 0.001
R15151 VSS.n8557 VSS.n8541 0.001
R15152 VSS.n8557 VSS.n8547 0.001
R15153 VSS.n8557 VSS.n8551 0.001
R15154 VSS.n8482 VSS.n8455 0.001
R15155 VSS.n8482 VSS.n8445 0.001
R15156 VSS.n8482 VSS.n8440 0.001
R15157 VSS.n9415 VSS.n9412 0.001
R15158 VSS.n9415 VSS.n9405 0.001
R15159 VSS.n9415 VSS.n9399 0.001
R15160 VSS.n9415 VSS.n9393 0.001
R15161 VSS.n9415 VSS.n9387 0.001
R15162 VSS.n9415 VSS.n9381 0.001
R15163 VSS.n9416 VSS.n9415 0.001
R15164 VSS.n9415 VSS.n9375 0.001
R15165 VSS.n9788 VSS.n9785 0.001
R15166 VSS.n9785 VSS.n7402 0.001
R15167 VSS.n9785 VSS.n7408 0.001
R15168 VSS.n9785 VSS.n7412 0.001
R15169 VSS.n9785 VSS.n7388 0.001
R15170 VSS.n9785 VSS.n7418 0.001
R15171 VSS.n9785 VSS.n9782 0.001
R15172 VSS.n7472 VSS.n7469 0.001
R15173 VSS.n7472 VSS.n7462 0.001
R15174 VSS.n7472 VSS.n7456 0.001
R15175 VSS.n7472 VSS.n7450 0.001
R15176 VSS.n7472 VSS.n7444 0.001
R15177 VSS.n7472 VSS.n7438 0.001
R15178 VSS.n7473 VSS.n7472 0.001
R15179 VSS.n7472 VSS.n7432 0.001
R15180 VSS.n10835 VSS.n10832 0.001
R15181 VSS.n10832 VSS.n3938 0.001
R15182 VSS.n10832 VSS.n3944 0.001
R15183 VSS.n10832 VSS.n3948 0.001
R15184 VSS.n10832 VSS.n3924 0.001
R15185 VSS.n10832 VSS.n3954 0.001
R15186 VSS.n10832 VSS.n10829 0.001
R15187 VSS.n9444 VSS.n9345 0.001
R15188 VSS.n9444 VSS.n9351 0.001
R15189 VSS.n9444 VSS.n9435 0.001
R15190 VSS.n9109 VSS.n9106 0.001
R15191 VSS.n9109 VSS.n9099 0.001
R15192 VSS.n9109 VSS.n9093 0.001
R15193 VSS.n9109 VSS.n9087 0.001
R15194 VSS.n9109 VSS.n9081 0.001
R15195 VSS.n9109 VSS.n9075 0.001
R15196 VSS.n9110 VSS.n9109 0.001
R15197 VSS.n9109 VSS.n9069 0.001
R15198 VSS.n9447 VSS.n9444 0.001
R15199 VSS.n9444 VSS.n9335 0.001
R15200 VSS.n9444 VSS.n9329 0.001
R15201 VSS.n9444 VSS.n9323 0.001
R15202 VSS.n9516 VSS.n9015 0.001
R15203 VSS.n9517 VSS.n9516 0.001
R15204 VSS.n9516 VSS.n9014 0.001
R15205 VSS.n9516 VSS.n9005 0.001
R15206 VSS.n9516 VSS.n9003 0.001
R15207 VSS.n9516 VSS.n9002 0.001
R15208 VSS.n9516 VSS.n9001 0.001
R15209 VSS.n9516 VSS.n9000 0.001
R15210 VSS.n9292 VSS.n9016 0.001
R15211 VSS.n9308 VSS.n9016 0.001
R15212 VSS.n9301 VSS.n9016 0.001
R15213 VSS.n9299 VSS.n9016 0.001
R15214 VSS.n9493 VSS.n9016 0.001
R15215 VSS.n9502 VSS.n9016 0.001
R15216 VSS.n9505 VSS.n9016 0.001
R15217 VSS.n7233 VSS.n7180 0.001
R15218 VSS.n7226 VSS.n7180 0.001
R15219 VSS.n7236 VSS.n7180 0.001
R15220 VSS.n9838 VSS.n7179 0.001
R15221 VSS.n9839 VSS.n9838 0.001
R15222 VSS.n9838 VSS.n7178 0.001
R15223 VSS.n9838 VSS.n7169 0.001
R15224 VSS.n9838 VSS.n7167 0.001
R15225 VSS.n9838 VSS.n7166 0.001
R15226 VSS.n9838 VSS.n7165 0.001
R15227 VSS.n9838 VSS.n7164 0.001
R15228 VSS.n9827 VSS.n7180 0.001
R15229 VSS.n9824 VSS.n7180 0.001
R15230 VSS.n9817 VSS.n7180 0.001
R15231 VSS.n7257 VSS.n7208 0.001
R15232 VSS.n7213 VSS.n7208 0.001
R15233 VSS.n7248 VSS.n7208 0.001
R15234 VSS.n7245 VSS.n7208 0.001
R15235 VSS.n7367 VSS.n7274 0.001
R15236 VSS.n7367 VSS.n7273 0.001
R15237 VSS.n7367 VSS.n7271 0.001
R15238 VSS.n7367 VSS.n7270 0.001
R15239 VSS.n7367 VSS.n7269 0.001
R15240 VSS.n7367 VSS.n7268 0.001
R15241 VSS.n7367 VSS.n7267 0.001
R15242 VSS.n7208 VSS.n7195 0.001
R15243 VSS.n7208 VSS.n7207 0.001
R15244 VSS.n7208 VSS.n7193 0.001
R15245 VSS.n9265 VSS.n9170 0.001
R15246 VSS.n9265 VSS.n9181 0.001
R15247 VSS.n9266 VSS.n9265 0.001
R15248 VSS.n9238 VSS.n9165 0.001
R15249 VSS.n9219 VSS.n9165 0.001
R15250 VSS.n9227 VSS.n9165 0.001
R15251 VSS.n9224 VSS.n9165 0.001
R15252 VSS.n9193 VSS.n9165 0.001
R15253 VSS.n9202 VSS.n9165 0.001
R15254 VSS.n9204 VSS.n9165 0.001
R15255 VSS.n9211 VSS.n9165 0.001
R15256 VSS.n9265 VSS.n9264 0.001
R15257 VSS.n9265 VSS.n9168 0.001
R15258 VSS.n9265 VSS.n9167 0.001
R15259 VSS.n9265 VSS.n9166 0.001
R15260 VSS.n8958 VSS.n7825 0.001
R15261 VSS.n8958 VSS.n7826 0.001
R15262 VSS.n8959 VSS.n8958 0.001
R15263 VSS.n8945 VSS.n7814 0.001
R15264 VSS.n7858 VSS.n7814 0.001
R15265 VSS.n7866 VSS.n7814 0.001
R15266 VSS.n7863 VSS.n7814 0.001
R15267 VSS.n7897 VSS.n7814 0.001
R15268 VSS.n7905 VSS.n7814 0.001
R15269 VSS.n7913 VSS.n7814 0.001
R15270 VSS.n7910 VSS.n7814 0.001
R15271 VSS.n8958 VSS.n8957 0.001
R15272 VSS.n8958 VSS.n7817 0.001
R15273 VSS.n8958 VSS.n7816 0.001
R15274 VSS.n7746 VSS.n7631 0.001
R15275 VSS.n7739 VSS.n7631 0.001
R15276 VSS.n7749 VSS.n7631 0.001
R15277 VSS.n8985 VSS.n7630 0.001
R15278 VSS.n8985 VSS.n7629 0.001
R15279 VSS.n8985 VSS.n7628 0.001
R15280 VSS.n8985 VSS.n7627 0.001
R15281 VSS.n8985 VSS.n7619 0.001
R15282 VSS.n8985 VSS.n7618 0.001
R15283 VSS.n8986 VSS.n8985 0.001
R15284 VSS.n8985 VSS.n7617 0.001
R15285 VSS.n7800 VSS.n7631 0.001
R15286 VSS.n7797 VSS.n7631 0.001
R15287 VSS.n7790 VSS.n7631 0.001
R15288 VSS.n7682 VSS.n7666 0.001
R15289 VSS.n7678 VSS.n7666 0.001
R15290 VSS.n7690 VSS.n7666 0.001
R15291 VSS.n7775 VSS.n7665 0.001
R15292 VSS.n7775 VSS.n7664 0.001
R15293 VSS.n7775 VSS.n7663 0.001
R15294 VSS.n7775 VSS.n7662 0.001
R15295 VSS.n7775 VSS.n7654 0.001
R15296 VSS.n7775 VSS.n7653 0.001
R15297 VSS.n7776 VSS.n7775 0.001
R15298 VSS.n7775 VSS.n7652 0.001
R15299 VSS.n7721 VSS.n7666 0.001
R15300 VSS.n7718 VSS.n7666 0.001
R15301 VSS.n7711 VSS.n7666 0.001
R15302 VSS.n9894 VSS.n7087 0.001
R15303 VSS.n7087 VSS.n7074 0.001
R15304 VSS.n7087 VSS.n7075 0.001
R15305 VSS.n7087 VSS.n7086 0.001
R15306 VSS.n7137 VSS.n7118 0.001
R15307 VSS.n7137 VSS.n7117 0.001
R15308 VSS.n7137 VSS.n7115 0.001
R15309 VSS.n7137 VSS.n7097 0.001
R15310 VSS.n7137 VSS.n7096 0.001
R15311 VSS.n7137 VSS.n7095 0.001
R15312 VSS.n7137 VSS.n7094 0.001
R15313 VSS.n9874 VSS.n7087 0.001
R15314 VSS.n9881 VSS.n7087 0.001
R15315 VSS.n9883 VSS.n7087 0.001
R15316 VSS.n8932 VSS.n7889 0.001
R15317 VSS.n8932 VSS.n7890 0.001
R15318 VSS.n8932 VSS.n7891 0.001
R15319 VSS.n8920 VSS.n7877 0.001
R15320 VSS.n8904 VSS.n7877 0.001
R15321 VSS.n8911 VSS.n7877 0.001
R15322 VSS.n8906 VSS.n7877 0.001
R15323 VSS.n7995 VSS.n7877 0.001
R15324 VSS.n7991 VSS.n7877 0.001
R15325 VSS.n7981 VSS.n7877 0.001
R15326 VSS.n8932 VSS.n8931 0.001
R15327 VSS.n8933 VSS.n8932 0.001
R15328 VSS.n8932 VSS.n7887 0.001
R15329 VSS.n8932 VSS.n7878 0.001
R15330 VSS.n6854 VSS.n6853 0.001
R15331 VSS.n6854 VSS.n6641 0.001
R15332 VSS.n6854 VSS.n6640 0.001
R15333 VSS.n6854 VSS.n6639 0.001
R15334 VSS.n6854 VSS.n6637 0.001
R15335 VSS.n6854 VSS.n6636 0.001
R15336 VSS.n6854 VSS.n6635 0.001
R15337 VSS.n6854 VSS.n6634 0.001
R15338 VSS.n6909 VSS.n6626 0.001
R15339 VSS.n6626 VSS.n6625 0.001
R15340 VSS.n6626 VSS.n6614 0.001
R15341 VSS.n6626 VSS.n6613 0.001
R15342 VSS.n6889 VSS.n6626 0.001
R15343 VSS.n6896 VSS.n6626 0.001
R15344 VSS.n6899 VSS.n6626 0.001
R15345 VSS.n6921 VSS.n6920 0.001
R15346 VSS.n6921 VSS.n6593 0.001
R15347 VSS.n6921 VSS.n6592 0.001
R15348 VSS.n6921 VSS.n6591 0.001
R15349 VSS.n6921 VSS.n6589 0.001
R15350 VSS.n6921 VSS.n6588 0.001
R15351 VSS.n6921 VSS.n6587 0.001
R15352 VSS.n6921 VSS.n6586 0.001
R15353 VSS.n6982 VSS.n6578 0.001
R15354 VSS.n6578 VSS.n6577 0.001
R15355 VSS.n6578 VSS.n6566 0.001
R15356 VSS.n6578 VSS.n6565 0.001
R15357 VSS.n6962 VSS.n6578 0.001
R15358 VSS.n6969 VSS.n6578 0.001
R15359 VSS.n6972 VSS.n6578 0.001
R15360 VSS.n7040 VSS.n6527 0.001
R15361 VSS.n7040 VSS.n6528 0.001
R15362 VSS.n7041 VSS.n7040 0.001
R15363 VSS.n6993 VSS.n6516 0.001
R15364 VSS.n6547 VSS.n6516 0.001
R15365 VSS.n6555 VSS.n6516 0.001
R15366 VSS.n6552 VSS.n6516 0.001
R15367 VSS.n6932 VSS.n6516 0.001
R15368 VSS.n6940 VSS.n6516 0.001
R15369 VSS.n6948 VSS.n6516 0.001
R15370 VSS.n6945 VSS.n6516 0.001
R15371 VSS.n7040 VSS.n7039 0.001
R15372 VSS.n7040 VSS.n6519 0.001
R15373 VSS.n7040 VSS.n6518 0.001
R15374 VSS.n6469 VSS.n6289 0.001
R15375 VSS.n6477 VSS.n6289 0.001
R15376 VSS.n6465 VSS.n6289 0.001
R15377 VSS.n7053 VSS.n7052 0.001
R15378 VSS.n7053 VSS.n6495 0.001
R15379 VSS.n7053 VSS.n6494 0.001
R15380 VSS.n7053 VSS.n6493 0.001
R15381 VSS.n7053 VSS.n6491 0.001
R15382 VSS.n7053 VSS.n6490 0.001
R15383 VSS.n7053 VSS.n6489 0.001
R15384 VSS.n7053 VSS.n6488 0.001
R15385 VSS.n6289 VSS.n6274 0.001
R15386 VSS.n6289 VSS.n6288 0.001
R15387 VSS.n6289 VSS.n6276 0.001
R15388 VSS.n6456 VSS.n6314 0.001
R15389 VSS.n6314 VSS.n6301 0.001
R15390 VSS.n6314 VSS.n6302 0.001
R15391 VSS.n6314 VSS.n6313 0.001
R15392 VSS.n6421 VSS.n6328 0.001
R15393 VSS.n6421 VSS.n6327 0.001
R15394 VSS.n6421 VSS.n6325 0.001
R15395 VSS.n6421 VSS.n6324 0.001
R15396 VSS.n6421 VSS.n6323 0.001
R15397 VSS.n6421 VSS.n6322 0.001
R15398 VSS.n6421 VSS.n6321 0.001
R15399 VSS.n6436 VSS.n6314 0.001
R15400 VSS.n6443 VSS.n6314 0.001
R15401 VSS.n6445 VSS.n6314 0.001
R15402 VSS.n6831 VSS.n6674 0.001
R15403 VSS.n6822 VSS.n6674 0.001
R15404 VSS.n6829 VSS.n6674 0.001
R15405 VSS.n6786 VSS.n6785 0.001
R15406 VSS.n6786 VSS.n6687 0.001
R15407 VSS.n6786 VSS.n6686 0.001
R15408 VSS.n6786 VSS.n6685 0.001
R15409 VSS.n6786 VSS.n6683 0.001
R15410 VSS.n6786 VSS.n6682 0.001
R15411 VSS.n6786 VSS.n6681 0.001
R15412 VSS.n6842 VSS.n6674 0.001
R15413 VSS.n6674 VSS.n6673 0.001
R15414 VSS.n6674 VSS.n6662 0.001
R15415 VSS.n6674 VSS.n6661 0.001
R15416 VSS.n6042 VSS.n6039 0.001
R15417 VSS.n6042 VSS.n6032 0.001
R15418 VSS.n6042 VSS.n6026 0.001
R15419 VSS.n6042 VSS.n6020 0.001
R15420 VSS.n6042 VSS.n6014 0.001
R15421 VSS.n6042 VSS.n6008 0.001
R15422 VSS.n6043 VSS.n6042 0.001
R15423 VSS.n6042 VSS.n6002 0.001
R15424 VSS.n5898 VSS.n5895 0.001
R15425 VSS.n5895 VSS.n5882 0.001
R15426 VSS.n5895 VSS.n5876 0.001
R15427 VSS.n5895 VSS.n5870 0.001
R15428 VSS.n5895 VSS.n5866 0.001
R15429 VSS.n5895 VSS.n5860 0.001
R15430 VSS.n5895 VSS.n5854 0.001
R15431 VSS.n5844 VSS.n5841 0.001
R15432 VSS.n5844 VSS.n5834 0.001
R15433 VSS.n5844 VSS.n5828 0.001
R15434 VSS.n5844 VSS.n5822 0.001
R15435 VSS.n5844 VSS.n5816 0.001
R15436 VSS.n5844 VSS.n5810 0.001
R15437 VSS.n5845 VSS.n5844 0.001
R15438 VSS.n5844 VSS.n5804 0.001
R15439 VSS.n5717 VSS.n5714 0.001
R15440 VSS.n5714 VSS.n5701 0.001
R15441 VSS.n5714 VSS.n5695 0.001
R15442 VSS.n5714 VSS.n5689 0.001
R15443 VSS.n5714 VSS.n5685 0.001
R15444 VSS.n5714 VSS.n5679 0.001
R15445 VSS.n5714 VSS.n5673 0.001
R15446 VSS.n5663 VSS.n5660 0.001
R15447 VSS.n5663 VSS.n5653 0.001
R15448 VSS.n5663 VSS.n5647 0.001
R15449 VSS.n5663 VSS.n5641 0.001
R15450 VSS.n5663 VSS.n5635 0.001
R15451 VSS.n5663 VSS.n5629 0.001
R15452 VSS.n5664 VSS.n5663 0.001
R15453 VSS.n5663 VSS.n5623 0.001
R15454 VSS.n5537 VSS.n5534 0.001
R15455 VSS.n5534 VSS.n5521 0.001
R15456 VSS.n5534 VSS.n5515 0.001
R15457 VSS.n5534 VSS.n5509 0.001
R15458 VSS.n5534 VSS.n5505 0.001
R15459 VSS.n5534 VSS.n5499 0.001
R15460 VSS.n5534 VSS.n5493 0.001
R15461 VSS.n5483 VSS.n5480 0.001
R15462 VSS.n5483 VSS.n5473 0.001
R15463 VSS.n5483 VSS.n5467 0.001
R15464 VSS.n5483 VSS.n5461 0.001
R15465 VSS.n5483 VSS.n5455 0.001
R15466 VSS.n5483 VSS.n5449 0.001
R15467 VSS.n5484 VSS.n5483 0.001
R15468 VSS.n5483 VSS.n5443 0.001
R15469 VSS.n5357 VSS.n5354 0.001
R15470 VSS.n5354 VSS.n5341 0.001
R15471 VSS.n5354 VSS.n5335 0.001
R15472 VSS.n5354 VSS.n5329 0.001
R15473 VSS.n5354 VSS.n5325 0.001
R15474 VSS.n5354 VSS.n5319 0.001
R15475 VSS.n5354 VSS.n5313 0.001
R15476 VSS.n5303 VSS.n5300 0.001
R15477 VSS.n5303 VSS.n5293 0.001
R15478 VSS.n5303 VSS.n5287 0.001
R15479 VSS.n5303 VSS.n5281 0.001
R15480 VSS.n5303 VSS.n5275 0.001
R15481 VSS.n5303 VSS.n5269 0.001
R15482 VSS.n5304 VSS.n5303 0.001
R15483 VSS.n5303 VSS.n5263 0.001
R15484 VSS.n10091 VSS.n10088 0.001
R15485 VSS.n10088 VSS.n10075 0.001
R15486 VSS.n10088 VSS.n10069 0.001
R15487 VSS.n10088 VSS.n10063 0.001
R15488 VSS.n10088 VSS.n10059 0.001
R15489 VSS.n10088 VSS.n10053 0.001
R15490 VSS.n10088 VSS.n10047 0.001
R15491 VSS.n4624 VSS.n4586 0.001
R15492 VSS.n4624 VSS.n4592 0.001
R15493 VSS.n4624 VSS.n4598 0.001
R15494 VSS.n4624 VSS.n4602 0.001
R15495 VSS.n3809 VSS.n3808 0.001
R15496 VSS.n3809 VSS.n3802 0.001
R15497 VSS.n3809 VSS.n3790 0.001
R15498 VSS.n3809 VSS.n3781 0.001
R15499 VSS.n3809 VSS.n3775 0.001
R15500 VSS.n3809 VSS.n3769 0.001
R15501 VSS.n3809 VSS.n3765 0.001
R15502 VSS.n4624 VSS.n4617 0.001
R15503 VSS.n4624 VSS.n4623 0.001
R15504 VSS.n4627 VSS.n4624 0.001
R15505 VSS.n6079 VSS.n6055 0.001
R15506 VSS.n6079 VSS.n6061 0.001
R15507 VSS.n6079 VSS.n6067 0.001
R15508 VSS.n6079 VSS.n6072 0.001
R15509 VSS.n6080 VSS.n6079 0.001
R15510 VSS.n6079 VSS.n5986 0.001
R15511 VSS.n6079 VSS.n5980 0.001
R15512 VSS.n6203 VSS.n6176 0.001
R15513 VSS.n6203 VSS.n6170 0.001
R15514 VSS.n6203 VSS.n6166 0.001
R15515 VSS.n6203 VSS.n6161 0.001
R15516 VSS.n11107 VSS.n11106 0.001
R15517 VSS.n11107 VSS.n11100 0.001
R15518 VSS.n11107 VSS.n11094 0.001
R15519 VSS.n11107 VSS.n11088 0.001
R15520 VSS.n11137 VSS.n11134 0.001
R15521 VSS.n11134 VSS.n3727 0.001
R15522 VSS.n11134 VSS.n3733 0.001
R15523 VSS.n11134 VSS.n3737 0.001
R15524 VSS.n11134 VSS.n3747 0.001
R15525 VSS.n11134 VSS.n3753 0.001
R15526 VSS.n11134 VSS.n11130 0.001
R15527 VSS.n11107 VSS.n11066 0.001
R15528 VSS.n11108 VSS.n11107 0.001
R15529 VSS.n11107 VSS.n11056 0.001
R15530 VSS.n6348 VSS.n3830 0.001
R15531 VSS.n6353 VSS.n3830 0.001
R15532 VSS.n6361 VSS.n3830 0.001
R15533 VSS.n6356 VSS.n3830 0.001
R15534 VSS.n6342 VSS.n3830 0.001
R15535 VSS.n6400 VSS.n3830 0.001
R15536 VSS.n6398 VSS.n3830 0.001
R15537 VSS.n11042 VSS.n3834 0.001
R15538 VSS.n11042 VSS.n3832 0.001
R15539 VSS.n11042 VSS.n3831 0.001
R15540 VSS.n10987 VSS.n3862 0.001
R15541 VSS.n10988 VSS.n10987 0.001
R15542 VSS.n10987 VSS.n3863 0.001
R15543 VSS.n10987 VSS.n3872 0.001
R15544 VSS.n10987 VSS.n3874 0.001
R15545 VSS.n10987 VSS.n3875 0.001
R15546 VSS.n10987 VSS.n3876 0.001
R15547 VSS.n10908 VSS.n3859 0.001
R15548 VSS.n10915 VSS.n3859 0.001
R15549 VSS.n10948 VSS.n3859 0.001
R15550 VSS.n7294 VSS.n3898 0.001
R15551 VSS.n7299 VSS.n3898 0.001
R15552 VSS.n7307 VSS.n3898 0.001
R15553 VSS.n7302 VSS.n3898 0.001
R15554 VSS.n7288 VSS.n3898 0.001
R15555 VSS.n7346 VSS.n3898 0.001
R15556 VSS.n7344 VSS.n3898 0.001
R15557 VSS.n10891 VSS.n3902 0.001
R15558 VSS.n10891 VSS.n3900 0.001
R15559 VSS.n10891 VSS.n3899 0.001
R15560 VSS.n4019 VSS.n3981 0.001
R15561 VSS.n4019 VSS.n3987 0.001
R15562 VSS.n4019 VSS.n3993 0.001
R15563 VSS.n4019 VSS.n3997 0.001
R15564 VSS.n4019 VSS.n4007 0.001
R15565 VSS.n4019 VSS.n4013 0.001
R15566 VSS.n4020 VSS.n4019 0.001
R15567 VSS.n4083 VSS.n4049 0.001
R15568 VSS.n4084 VSS.n4083 0.001
R15569 VSS.n4083 VSS.n4039 0.001
R15570 VSS.n4140 VSS.n4114 0.001
R15571 VSS.n4147 VSS.n4114 0.001
R15572 VSS.n4142 VSS.n4114 0.001
R15573 VSS.n4447 VSS.n4114 0.001
R15574 VSS.n4404 VSS.n4193 0.001
R15575 VSS.n4404 VSS.n4192 0.001
R15576 VSS.n4404 VSS.n4191 0.001
R15577 VSS.n4405 VSS.n4185 0.001
R15578 VSS.n4405 VSS.n4184 0.001
R15579 VSS.n4405 VSS.n4183 0.001
R15580 VSS.n4405 VSS.n4182 0.001
R15581 VSS.n4344 VSS.n4343 0.001
R15582 VSS.n4344 VSS.n4253 0.001
R15583 VSS.n4344 VSS.n4252 0.001
R15584 VSS.n4344 VSS.n4250 0.001
R15585 VSS.n4305 VSS.n4234 0.001
R15586 VSS.n4319 VSS.n4234 0.001
R15587 VSS.n4308 VSS.n4234 0.001
R15588 VSS.n4312 VSS.n4234 0.001
R15589 VSS.n4285 VSS.n4234 0.001
R15590 VSS.n4292 VSS.n4234 0.001
R15591 VSS.n4294 VSS.n4234 0.001
R15592 VSS.n4344 VSS.n4237 0.001
R15593 VSS.n4344 VSS.n4235 0.001
R15594 VSS.n4345 VSS.n4344 0.001
R15595 VSS.n4404 VSS.n4189 0.001
R15596 VSS.n4404 VSS.n4194 0.001
R15597 VSS.n4404 VSS.n4196 0.001
R15598 VSS.n4405 VSS.n4168 0.001
R15599 VSS.n4405 VSS.n4167 0.001
R15600 VSS.n4405 VSS.n4166 0.001
R15601 VSS.n4406 VSS.n4405 0.001
R15602 VSS.n10776 VSS.n4115 0.001
R15603 VSS.n10776 VSS.n4116 0.001
R15604 VSS.n10776 VSS.n4117 0.001
R15605 VSS.n10776 VSS.n4118 0.001
R15606 VSS.n10776 VSS.n4126 0.001
R15607 VSS.n10777 VSS.n10776 0.001
R15608 VSS.n10776 VSS.n4127 0.001
R15609 VSS.n10756 VSS.n4114 0.001
R15610 VSS.n10764 VSS.n4114 0.001
R15611 VSS.n10765 VSS.n4114 0.001
R15612 VSS.n1296 VSS.n1284 0.001
R15613 VSS.n1296 VSS.n1278 0.001
R15614 VSS.n1297 VSS.n1296 0.001
R15615 VSS.n790 VSS.n786 0.001
R15616 VSS.n790 VSS.n780 0.001
R15617 VSS.n791 VSS.n790 0.001
R15618 VSS.n790 VSS.n680 0.001
R15619 VSS.n790 VSS.n674 0.001
R15620 VSS.n790 VSS.n668 0.001
R15621 VSS.n790 VSS.n664 0.001
R15622 VSS.n1296 VSS.n1295 0.001
R15623 VSS.n1296 VSS.n1264 0.001
R15624 VSS.n1296 VSS.n1258 0.001
R15625 VSS.n1296 VSS.n1252 0.001
R15626 VSS.n1345 VSS.n1222 0.001
R15627 VSS.n1345 VSS.n1228 0.001
R15628 VSS.n1345 VSS.n1336 0.001
R15629 VSS.n1047 VSS.n1044 0.001
R15630 VSS.n1047 VSS.n1037 0.001
R15631 VSS.n1047 VSS.n1031 0.001
R15632 VSS.n1047 VSS.n1025 0.001
R15633 VSS.n1047 VSS.n1019 0.001
R15634 VSS.n1047 VSS.n1013 0.001
R15635 VSS.n1048 VSS.n1047 0.001
R15636 VSS.n1047 VSS.n1007 0.001
R15637 VSS.n1348 VSS.n1345 0.001
R15638 VSS.n1345 VSS.n1212 0.001
R15639 VSS.n1345 VSS.n1206 0.001
R15640 VSS.n1345 VSS.n1200 0.001
R15641 VSS.n1106 VSS.n970 0.001
R15642 VSS.n1106 VSS.n976 0.001
R15643 VSS.n1106 VSS.n1086 0.001
R15644 VSS.n14332 VSS.n14328 0.001
R15645 VSS.n14332 VSS.n14322 0.001
R15646 VSS.n14332 VSS.n14318 0.001
R15647 VSS.n14332 VSS.n14313 0.001
R15648 VSS.n14228 VSS.n575 0.001
R15649 VSS.n14228 VSS.n574 0.001
R15650 VSS.n14228 VSS.n573 0.001
R15651 VSS.n14229 VSS.n557 0.001
R15652 VSS.n14230 VSS.n14229 0.001
R15653 VSS.n14229 VSS.n548 0.001
R15654 VSS.n10704 VSS.n10692 0.001
R15655 VSS.n10705 VSS.n10704 0.001
R15656 VSS.n10704 VSS.n10687 0.001
R15657 VSS.n10704 VSS.n10681 0.001
R15658 VSS.n14275 VSS.n14271 0.001
R15659 VSS.n14276 VSS.n14275 0.001
R15660 VSS.n14275 VSS.n14259 0.001
R15661 VSS.n14275 VSS.n535 0.001
R15662 VSS.n14275 VSS.n529 0.001
R15663 VSS.n14275 VSS.n523 0.001
R15664 VSS.n14275 VSS.n519 0.001
R15665 VSS.n10704 VSS.n10703 0.001
R15666 VSS.n10704 VSS.n10670 0.001
R15667 VSS.n10704 VSS.n10664 0.001
R15668 VSS.n10704 VSS.n10658 0.001
R15669 VSS.n14202 VSS.n602 0.001
R15670 VSS.n602 VSS.n587 0.001
R15671 VSS.n602 VSS.n601 0.001
R15672 VSS.n602 VSS.n589 0.001
R15673 VSS.n1151 VSS.n932 0.001
R15674 VSS.n1151 VSS.n931 0.001
R15675 VSS.n1151 VSS.n930 0.001
R15676 VSS.n1151 VSS.n913 0.001
R15677 VSS.n1152 VSS.n1151 0.001
R15678 VSS.n1151 VSS.n927 0.001
R15679 VSS.n1151 VSS.n917 0.001
R15680 VSS.n1151 VSS.n916 0.001
R15681 VSS.n14177 VSS.n602 0.001
R15682 VSS.n14192 VSS.n602 0.001
R15683 VSS.n14180 VSS.n602 0.001
R15684 VSS.n14185 VSS.n602 0.001
R15685 VSS.n12453 VSS.n12450 0.001
R15686 VSS.n12453 VSS.n12444 0.001
R15687 VSS.n12453 VSS.n12438 0.001
R15688 VSS.n12453 VSS.n12394 0.001
R15689 VSS.n12416 VSS.n2478 0.001
R15690 VSS.n12412 VSS.n2478 0.001
R15691 VSS.n12406 VSS.n2478 0.001
R15692 VSS.n12404 VSS.n2478 0.001
R15693 VSS.n13045 VSS.n2494 0.001
R15694 VSS.n13045 VSS.n2493 0.001
R15695 VSS.n13045 VSS.n2491 0.001
R15696 VSS.n13045 VSS.n2490 0.001
R15697 VSS.n13045 VSS.n2489 0.001
R15698 VSS.n13045 VSS.n2488 0.001
R15699 VSS.n13045 VSS.n2487 0.001
R15700 VSS.n13055 VSS.n2478 0.001
R15701 VSS.n2478 VSS.n2477 0.001
R15702 VSS.n2478 VSS.n2466 0.001
R15703 VSS.n2451 VSS.n2356 0.001
R15704 VSS.n2441 VSS.n2356 0.001
R15705 VSS.n2440 VSS.n2356 0.001
R15706 VSS.n2432 VSS.n2356 0.001
R15707 VSS.n13102 VSS.n13101 0.001
R15708 VSS.n13101 VSS.n2370 0.001
R15709 VSS.n13101 VSS.n2362 0.001
R15710 VSS.n13101 VSS.n2361 0.001
R15711 VSS.n13101 VSS.n2360 0.001
R15712 VSS.n13101 VSS.n2359 0.001
R15713 VSS.n13101 VSS.n2358 0.001
R15714 VSS.n13071 VSS.n2356 0.001
R15715 VSS.n13086 VSS.n2356 0.001
R15716 VSS.n13074 VSS.n2356 0.001
R15717 VSS.n13079 VSS.n2356 0.001
R15718 VSS.n13135 VSS.n1928 0.001
R15719 VSS.n1928 VSS.n1915 0.001
R15720 VSS.n1928 VSS.n1916 0.001
R15721 VSS.n1928 VSS.n1927 0.001
R15722 VSS.n2342 VSS.n1942 0.001
R15723 VSS.n2342 VSS.n1941 0.001
R15724 VSS.n2342 VSS.n1940 0.001
R15725 VSS.n2342 VSS.n1939 0.001
R15726 VSS.n2342 VSS.n1938 0.001
R15727 VSS.n2342 VSS.n1937 0.001
R15728 VSS.n2342 VSS.n1936 0.001
R15729 VSS.n2342 VSS.n1935 0.001
R15730 VSS.n13124 VSS.n1928 0.001
R15731 VSS.n13122 VSS.n1928 0.001
R15732 VSS.n13115 VSS.n1928 0.001
R15733 VSS.n14228 VSS.n571 0.001
R15734 VSS.n14228 VSS.n576 0.001
R15735 VSS.n14228 VSS.n578 0.001
R15736 VSS.n14229 VSS.n553 0.001
R15737 VSS.n14229 VSS.n552 0.001
R15738 VSS.n14229 VSS.n551 0.001
R15739 VSS.n14229 VSS.n550 0.001
R15740 VSS.n1165 VSS.n1164 0.001
R15741 VSS.n1165 VSS.n894 0.001
R15742 VSS.n1165 VSS.n893 0.001
R15743 VSS.n1165 VSS.n892 0.001
R15744 VSS.n1165 VSS.n890 0.001
R15745 VSS.n1165 VSS.n889 0.001
R15746 VSS.n1165 VSS.n888 0.001
R15747 VSS.n1165 VSS.n887 0.001
R15748 VSS.n1397 VSS.n879 0.001
R15749 VSS.n879 VSS.n866 0.001
R15750 VSS.n879 VSS.n867 0.001
R15751 VSS.n879 VSS.n878 0.001
R15752 VSS.n1375 VSS.n879 0.001
R15753 VSS.n1384 VSS.n879 0.001
R15754 VSS.n1387 VSS.n879 0.001
R15755 VSS.n1109 VSS.n1106 0.001
R15756 VSS.n1106 VSS.n1092 0.001
R15757 VSS.n1106 VSS.n1098 0.001
R15758 VSS.n1106 VSS.n1102 0.001
R15759 VSS.n14332 VSS.n14299 0.001
R15760 VSS.n14332 VSS.n14293 0.001
R15761 VSS.n14333 VSS.n14332 0.001
R15762 VSS.n14332 VSS.n14287 0.001
R15763 VSS.n1569 VSS.n1566 0.001
R15764 VSS.n1569 VSS.n1559 0.001
R15765 VSS.n1569 VSS.n1553 0.001
R15766 VSS.n1569 VSS.n1547 0.001
R15767 VSS.n1569 VSS.n1541 0.001
R15768 VSS.n1569 VSS.n1535 0.001
R15769 VSS.n1570 VSS.n1569 0.001
R15770 VSS.n1569 VSS.n1529 0.001
R15771 VSS.n13856 VSS.n13853 0.001
R15772 VSS.n13853 VSS.n13725 0.001
R15773 VSS.n13853 VSS.n13731 0.001
R15774 VSS.n13853 VSS.n13735 0.001
R15775 VSS.n13853 VSS.n13711 0.001
R15776 VSS.n13853 VSS.n13741 0.001
R15777 VSS.n13853 VSS.n13850 0.001
R15778 VSS.n13809 VSS.n13806 0.001
R15779 VSS.n13809 VSS.n13799 0.001
R15780 VSS.n13809 VSS.n13793 0.001
R15781 VSS.n13809 VSS.n13787 0.001
R15782 VSS.n13809 VSS.n13781 0.001
R15783 VSS.n13809 VSS.n13775 0.001
R15784 VSS.n13810 VSS.n13809 0.001
R15785 VSS.n13809 VSS.n13769 0.001
R15786 VSS.n13391 VSS.n13388 0.001
R15787 VSS.n13388 VSS.n13262 0.001
R15788 VSS.n13388 VSS.n13268 0.001
R15789 VSS.n13388 VSS.n13272 0.001
R15790 VSS.n13388 VSS.n13248 0.001
R15791 VSS.n13388 VSS.n13278 0.001
R15792 VSS.n13388 VSS.n13385 0.001
R15793 VSS.n1616 VSS.n1491 0.001
R15794 VSS.n1616 VSS.n1497 0.001
R15795 VSS.n1616 VSS.n1607 0.001
R15796 VSS.n762 VSS.n759 0.001
R15797 VSS.n762 VSS.n752 0.001
R15798 VSS.n762 VSS.n746 0.001
R15799 VSS.n762 VSS.n740 0.001
R15800 VSS.n762 VSS.n734 0.001
R15801 VSS.n762 VSS.n728 0.001
R15802 VSS.n763 VSS.n762 0.001
R15803 VSS.n762 VSS.n722 0.001
R15804 VSS.n1619 VSS.n1616 0.001
R15805 VSS.n1616 VSS.n1481 0.001
R15806 VSS.n1616 VSS.n1475 0.001
R15807 VSS.n1616 VSS.n1469 0.001
R15808 VSS.n14115 VSS.n649 0.001
R15809 VSS.n14116 VSS.n14115 0.001
R15810 VSS.n14115 VSS.n648 0.001
R15811 VSS.n14115 VSS.n639 0.001
R15812 VSS.n14115 VSS.n637 0.001
R15813 VSS.n14115 VSS.n636 0.001
R15814 VSS.n14115 VSS.n635 0.001
R15815 VSS.n14115 VSS.n634 0.001
R15816 VSS.n1689 VSS.n650 0.001
R15817 VSS.n1692 VSS.n650 0.001
R15818 VSS.n1682 VSS.n650 0.001
R15819 VSS.n1677 VSS.n650 0.001
R15820 VSS.n14092 VSS.n650 0.001
R15821 VSS.n14101 VSS.n650 0.001
R15822 VSS.n14104 VSS.n650 0.001
R15823 VSS.n13682 VSS.n1661 0.001
R15824 VSS.n13690 VSS.n1661 0.001
R15825 VSS.n13678 VSS.n1661 0.001
R15826 VSS.n14079 VSS.n1660 0.001
R15827 VSS.n14079 VSS.n1659 0.001
R15828 VSS.n14079 VSS.n1658 0.001
R15829 VSS.n14079 VSS.n1657 0.001
R15830 VSS.n14079 VSS.n1649 0.001
R15831 VSS.n14079 VSS.n1648 0.001
R15832 VSS.n14080 VSS.n14079 0.001
R15833 VSS.n14079 VSS.n1647 0.001
R15834 VSS.n13669 VSS.n1661 0.001
R15835 VSS.n13666 VSS.n1661 0.001
R15836 VSS.n13660 VSS.n1661 0.001
R15837 VSS.n13905 VSS.n13221 0.001
R15838 VSS.n13221 VSS.n13208 0.001
R15839 VSS.n13221 VSS.n13209 0.001
R15840 VSS.n13221 VSS.n13220 0.001
R15841 VSS.n13643 VSS.n13235 0.001
R15842 VSS.n13643 VSS.n13234 0.001
R15843 VSS.n13643 VSS.n13232 0.001
R15844 VSS.n13643 VSS.n13231 0.001
R15845 VSS.n13643 VSS.n13230 0.001
R15846 VSS.n13643 VSS.n13229 0.001
R15847 VSS.n13643 VSS.n13228 0.001
R15848 VSS.n13885 VSS.n13221 0.001
R15849 VSS.n13892 VSS.n13221 0.001
R15850 VSS.n13894 VSS.n13221 0.001
R15851 VSS.n1435 VSS.n823 0.001
R15852 VSS.n1435 VSS.n834 0.001
R15853 VSS.n1436 VSS.n1435 0.001
R15854 VSS.n1408 VSS.n818 0.001
R15855 VSS.n848 VSS.n818 0.001
R15856 VSS.n856 VSS.n818 0.001
R15857 VSS.n853 VSS.n818 0.001
R15858 VSS.n1182 VSS.n818 0.001
R15859 VSS.n1175 VSS.n818 0.001
R15860 VSS.n1189 VSS.n818 0.001
R15861 VSS.n1191 VSS.n818 0.001
R15862 VSS.n1435 VSS.n1434 0.001
R15863 VSS.n1435 VSS.n821 0.001
R15864 VSS.n1435 VSS.n820 0.001
R15865 VSS.n1435 VSS.n819 0.001
R15866 VSS.n2198 VSS.n2005 0.001
R15867 VSS.n2191 VSS.n2005 0.001
R15868 VSS.n2201 VSS.n2005 0.001
R15869 VSS.n2245 VSS.n2004 0.001
R15870 VSS.n2246 VSS.n2245 0.001
R15871 VSS.n2245 VSS.n2003 0.001
R15872 VSS.n2245 VSS.n1994 0.001
R15873 VSS.n2245 VSS.n1992 0.001
R15874 VSS.n2245 VSS.n1991 0.001
R15875 VSS.n2245 VSS.n1990 0.001
R15876 VSS.n2245 VSS.n1989 0.001
R15877 VSS.n2234 VSS.n2005 0.001
R15878 VSS.n2231 VSS.n2005 0.001
R15879 VSS.n2224 VSS.n2005 0.001
R15880 VSS.n2110 VSS.n2080 0.001
R15881 VSS.n2106 VSS.n2080 0.001
R15882 VSS.n2118 VSS.n2080 0.001
R15883 VSS.n2180 VSS.n2079 0.001
R15884 VSS.n2181 VSS.n2180 0.001
R15885 VSS.n2180 VSS.n2078 0.001
R15886 VSS.n2180 VSS.n2069 0.001
R15887 VSS.n2180 VSS.n2067 0.001
R15888 VSS.n2180 VSS.n2066 0.001
R15889 VSS.n2180 VSS.n2065 0.001
R15890 VSS.n2180 VSS.n2064 0.001
R15891 VSS.n2169 VSS.n2080 0.001
R15892 VSS.n2166 VSS.n2080 0.001
R15893 VSS.n2159 VSS.n2080 0.001
R15894 VSS.n12661 VSS.n1849 0.001
R15895 VSS.n12654 VSS.n1849 0.001
R15896 VSS.n12664 VSS.n1849 0.001
R15897 VSS.n13188 VSS.n13187 0.001
R15898 VSS.n13188 VSS.n1865 0.001
R15899 VSS.n13188 VSS.n1864 0.001
R15900 VSS.n13188 VSS.n1863 0.001
R15901 VSS.n13188 VSS.n1861 0.001
R15902 VSS.n13188 VSS.n1860 0.001
R15903 VSS.n13188 VSS.n1859 0.001
R15904 VSS.n13188 VSS.n1858 0.001
R15905 VSS.n1849 VSS.n1834 0.001
R15906 VSS.n1849 VSS.n1848 0.001
R15907 VSS.n1849 VSS.n1836 0.001
R15908 VSS.n12689 VSS.n1777 0.001
R15909 VSS.n12684 VSS.n1777 0.001
R15910 VSS.n12678 VSS.n1777 0.001
R15911 VSS.n12676 VSS.n1777 0.001
R15912 VSS.n13936 VSS.n13935 0.001
R15913 VSS.n13935 VSS.n1791 0.001
R15914 VSS.n13935 VSS.n1783 0.001
R15915 VSS.n13935 VSS.n1782 0.001
R15916 VSS.n13935 VSS.n1781 0.001
R15917 VSS.n13935 VSS.n1780 0.001
R15918 VSS.n13935 VSS.n1779 0.001
R15919 VSS.n1826 VSS.n1777 0.001
R15920 VSS.n1819 VSS.n1777 0.001
R15921 VSS.n13921 VSS.n1777 0.001
R15922 VSS.n2030 VSS.n1972 0.001
R15923 VSS.n2019 VSS.n1972 0.001
R15924 VSS.n2025 VSS.n1972 0.001
R15925 VSS.n2319 VSS.n1971 0.001
R15926 VSS.n2319 VSS.n1970 0.001
R15927 VSS.n2319 VSS.n1969 0.001
R15928 VSS.n2319 VSS.n1968 0.001
R15929 VSS.n2320 VSS.n2319 0.001
R15930 VSS.n2319 VSS.n1966 0.001
R15931 VSS.n2319 VSS.n1955 0.001
R15932 VSS.n2272 VSS.n1972 0.001
R15933 VSS.n2269 VSS.n1972 0.001
R15934 VSS.n2262 VSS.n1972 0.001
R15935 VSS.n2260 VSS.n1972 0.001
R15936 VSS.n12985 VSS.n2583 0.001
R15937 VSS.n12986 VSS.n12985 0.001
R15938 VSS.n12985 VSS.n2582 0.001
R15939 VSS.n12985 VSS.n2573 0.001
R15940 VSS.n12985 VSS.n2571 0.001
R15941 VSS.n12985 VSS.n2570 0.001
R15942 VSS.n12985 VSS.n2569 0.001
R15943 VSS.n12985 VSS.n2568 0.001
R15944 VSS.n2719 VSS.n2584 0.001
R15945 VSS.n2714 VSS.n2584 0.001
R15946 VSS.n2708 VSS.n2584 0.001
R15947 VSS.n2706 VSS.n2584 0.001
R15948 VSS.n12964 VSS.n2584 0.001
R15949 VSS.n12971 VSS.n2584 0.001
R15950 VSS.n12974 VSS.n2584 0.001
R15951 VSS.n12949 VSS.n2687 0.001
R15952 VSS.n12949 VSS.n2686 0.001
R15953 VSS.n12949 VSS.n2685 0.001
R15954 VSS.n12949 VSS.n2684 0.001
R15955 VSS.n12949 VSS.n2676 0.001
R15956 VSS.n12949 VSS.n2675 0.001
R15957 VSS.n12950 VSS.n12949 0.001
R15958 VSS.n12949 VSS.n2674 0.001
R15959 VSS.n2808 VSS.n2688 0.001
R15960 VSS.n2791 VSS.n2688 0.001
R15961 VSS.n2799 VSS.n2688 0.001
R15962 VSS.n2796 VSS.n2688 0.001
R15963 VSS.n2774 VSS.n2688 0.001
R15964 VSS.n2784 VSS.n2688 0.001
R15965 VSS.n2816 VSS.n2688 0.001
R15966 VSS.n12908 VSS.n2764 0.001
R15967 VSS.n12909 VSS.n12908 0.001
R15968 VSS.n12908 VSS.n2763 0.001
R15969 VSS.n12908 VSS.n2754 0.001
R15970 VSS.n12908 VSS.n2752 0.001
R15971 VSS.n12908 VSS.n2751 0.001
R15972 VSS.n12908 VSS.n2750 0.001
R15973 VSS.n12908 VSS.n2749 0.001
R15974 VSS.n2899 VSS.n2765 0.001
R15975 VSS.n2894 VSS.n2765 0.001
R15976 VSS.n2888 VSS.n2765 0.001
R15977 VSS.n2886 VSS.n2765 0.001
R15978 VSS.n12887 VSS.n2765 0.001
R15979 VSS.n12894 VSS.n2765 0.001
R15980 VSS.n12897 VSS.n2765 0.001
R15981 VSS.n12623 VSS.n2868 0.001
R15982 VSS.n12631 VSS.n2868 0.001
R15983 VSS.n12619 VSS.n2868 0.001
R15984 VSS.n12872 VSS.n2867 0.001
R15985 VSS.n12872 VSS.n2866 0.001
R15986 VSS.n12872 VSS.n2865 0.001
R15987 VSS.n12872 VSS.n2864 0.001
R15988 VSS.n12872 VSS.n2856 0.001
R15989 VSS.n12872 VSS.n2855 0.001
R15990 VSS.n12873 VSS.n12872 0.001
R15991 VSS.n12872 VSS.n2854 0.001
R15992 VSS.n3053 VSS.n2868 0.001
R15993 VSS.n3050 VSS.n2868 0.001
R15994 VSS.n3044 VSS.n2868 0.001
R15995 VSS.n3080 VSS.n2955 0.001
R15996 VSS.n3075 VSS.n2955 0.001
R15997 VSS.n3069 VSS.n2955 0.001
R15998 VSS.n3067 VSS.n2955 0.001
R15999 VSS.n12731 VSS.n12730 0.001
R16000 VSS.n12730 VSS.n2969 0.001
R16001 VSS.n12730 VSS.n2961 0.001
R16002 VSS.n12730 VSS.n2960 0.001
R16003 VSS.n12730 VSS.n2959 0.001
R16004 VSS.n12730 VSS.n2958 0.001
R16005 VSS.n12730 VSS.n2957 0.001
R16006 VSS.n3031 VSS.n2955 0.001
R16007 VSS.n3024 VSS.n2955 0.001
R16008 VSS.n12716 VSS.n2955 0.001
R16009 VSS.n2637 VSS.n2524 0.001
R16010 VSS.n2599 VSS.n2524 0.001
R16011 VSS.n2605 VSS.n2524 0.001
R16012 VSS.n13024 VSS.n2523 0.001
R16013 VSS.n13024 VSS.n2522 0.001
R16014 VSS.n13024 VSS.n2521 0.001
R16015 VSS.n13024 VSS.n2520 0.001
R16016 VSS.n13025 VSS.n13024 0.001
R16017 VSS.n13024 VSS.n2518 0.001
R16018 VSS.n13024 VSS.n2507 0.001
R16019 VSS.n2627 VSS.n2524 0.001
R16020 VSS.n2624 VSS.n2524 0.001
R16021 VSS.n2617 VSS.n2524 0.001
R16022 VSS.n2615 VSS.n2524 0.001
R16023 VSS.n11677 VSS.n11676 0.001
R16024 VSS.n11676 VSS.n11673 0.001
R16025 VSS.n11676 VSS.n11667 0.001
R16026 VSS.n11676 VSS.n11661 0.001
R16027 VSS.n11676 VSS.n11655 0.001
R16028 VSS.n11676 VSS.n11649 0.001
R16029 VSS.n11676 VSS.n11643 0.001
R16030 VSS.n11676 VSS.n11581 0.001
R16031 VSS.n12259 VSS.n12256 0.001
R16032 VSS.n12256 VSS.n12243 0.001
R16033 VSS.n12256 VSS.n12237 0.001
R16034 VSS.n12256 VSS.n12231 0.001
R16035 VSS.n12256 VSS.n12227 0.001
R16036 VSS.n12256 VSS.n12221 0.001
R16037 VSS.n12256 VSS.n12215 0.001
R16038 VSS.n11746 VSS.n11745 0.001
R16039 VSS.n11745 VSS.n11742 0.001
R16040 VSS.n11745 VSS.n11736 0.001
R16041 VSS.n11745 VSS.n11730 0.001
R16042 VSS.n11745 VSS.n11724 0.001
R16043 VSS.n11745 VSS.n11718 0.001
R16044 VSS.n11745 VSS.n11712 0.001
R16045 VSS.n11745 VSS.n11705 0.001
R16046 VSS.n12152 VSS.n12149 0.001
R16047 VSS.n12149 VSS.n12136 0.001
R16048 VSS.n12149 VSS.n12130 0.001
R16049 VSS.n12149 VSS.n12124 0.001
R16050 VSS.n12149 VSS.n12120 0.001
R16051 VSS.n12149 VSS.n12114 0.001
R16052 VSS.n12149 VSS.n12108 0.001
R16053 VSS.n12098 VSS.n12095 0.001
R16054 VSS.n12098 VSS.n12088 0.001
R16055 VSS.n12098 VSS.n12082 0.001
R16056 VSS.n12098 VSS.n12076 0.001
R16057 VSS.n12098 VSS.n12070 0.001
R16058 VSS.n12098 VSS.n12064 0.001
R16059 VSS.n12099 VSS.n12098 0.001
R16060 VSS.n12098 VSS.n12058 0.001
R16061 VSS.n11984 VSS.n11981 0.001
R16062 VSS.n11981 VSS.n11968 0.001
R16063 VSS.n11981 VSS.n11962 0.001
R16064 VSS.n11981 VSS.n11956 0.001
R16065 VSS.n11981 VSS.n11952 0.001
R16066 VSS.n11981 VSS.n11946 0.001
R16067 VSS.n11981 VSS.n11940 0.001
R16068 VSS.n11878 VSS.n11877 0.001
R16069 VSS.n11877 VSS.n11874 0.001
R16070 VSS.n11877 VSS.n11868 0.001
R16071 VSS.n11877 VSS.n11862 0.001
R16072 VSS.n11877 VSS.n11856 0.001
R16073 VSS.n11877 VSS.n11850 0.001
R16074 VSS.n11877 VSS.n11844 0.001
R16075 VSS.n11877 VSS.n11837 0.001
R16076 VSS.n3556 VSS.n3553 0.001
R16077 VSS.n3553 VSS.n3540 0.001
R16078 VSS.n3553 VSS.n3534 0.001
R16079 VSS.n3553 VSS.n3528 0.001
R16080 VSS.n3553 VSS.n3524 0.001
R16081 VSS.n3553 VSS.n3518 0.001
R16082 VSS.n3553 VSS.n3512 0.001
R16083 VSS.n3502 VSS.n3499 0.001
R16084 VSS.n3502 VSS.n3492 0.001
R16085 VSS.n3502 VSS.n3486 0.001
R16086 VSS.n3502 VSS.n3480 0.001
R16087 VSS.n3502 VSS.n3474 0.001
R16088 VSS.n3502 VSS.n3468 0.001
R16089 VSS.n3503 VSS.n3502 0.001
R16090 VSS.n3502 VSS.n3462 0.001
R16091 VSS.n12605 VSS.n12592 0.001
R16092 VSS.n12605 VSS.n3115 0.001
R16093 VSS.n12605 VSS.n3109 0.001
R16094 VSS.n12605 VSS.n3103 0.001
R16095 VSS.n12605 VSS.n3099 0.001
R16096 VSS.n12605 VSS.n3093 0.001
R16097 VSS.n12606 VSS.n12605 0.001
R16098 VSS.n3167 VSS.n3164 0.001
R16099 VSS.n3164 VSS.n3126 0.001
R16100 VSS.n3164 VSS.n3132 0.001
R16101 VSS.n3164 VSS.n3136 0.001
R16102 VSS.n3267 VSS.n3264 0.001
R16103 VSS.n3267 VSS.n3258 0.001
R16104 VSS.n3268 VSS.n3267 0.001
R16105 VSS.n3267 VSS.n3250 0.001
R16106 VSS.n3267 VSS.n3243 0.001
R16107 VSS.n3267 VSS.n3237 0.001
R16108 VSS.n3267 VSS.n3231 0.001
R16109 VSS.n3267 VSS.n3227 0.001
R16110 VSS.n3164 VSS.n3151 0.001
R16111 VSS.n3164 VSS.n3157 0.001
R16112 VSS.n3164 VSS.n3163 0.001
R16113 VSS.n11632 VSS.n11629 0.001
R16114 VSS.n11629 VSS.n11611 0.001
R16115 VSS.n11629 VSS.n11617 0.001
R16116 VSS.n11629 VSS.n11622 0.001
R16117 VSS.n11629 VSS.n11601 0.001
R16118 VSS.n11629 VSS.n11595 0.001
R16119 VSS.n11629 VSS.n11589 0.001
R16120 VSS.n12453 VSS.n12381 0.001
R16121 VSS.n12453 VSS.n12375 0.001
R16122 VSS.n12453 VSS.n12371 0.001
R16123 VSS.n12454 VSS.n12453 0.001
R16124 VSS.n2979 VSS.n2935 0.001
R16125 VSS.n2993 VSS.n2935 0.001
R16126 VSS.n2982 VSS.n2935 0.001
R16127 VSS.n2986 VSS.n2935 0.001
R16128 VSS.n12744 VSS.n2935 0.001
R16129 VSS.n12746 VSS.n2935 0.001
R16130 VSS.n12754 VSS.n2935 0.001
R16131 VSS.n12796 VSS.n2939 0.001
R16132 VSS.n12796 VSS.n2937 0.001
R16133 VSS.n12796 VSS.n2936 0.001
R16134 VSS.n13970 VSS.n1720 0.001
R16135 VSS.n13984 VSS.n1720 0.001
R16136 VSS.n13973 VSS.n1720 0.001
R16137 VSS.n13977 VSS.n1720 0.001
R16138 VSS.n13950 VSS.n1720 0.001
R16139 VSS.n13957 VSS.n1720 0.001
R16140 VSS.n13959 VSS.n1720 0.001
R16141 VSS.n14016 VSS.n1723 0.001
R16142 VSS.n14016 VSS.n1721 0.001
R16143 VSS.n14017 VSS.n14016 0.001
R16144 VSS.n13512 VSS.n13485 0.001
R16145 VSS.n13517 VSS.n13485 0.001
R16146 VSS.n13525 VSS.n13485 0.001
R16147 VSS.n13520 VSS.n13485 0.001
R16148 VSS.n13567 VSS.n13485 0.001
R16149 VSS.n13560 VSS.n13485 0.001
R16150 VSS.n13577 VSS.n13485 0.001
R16151 VSS.n13603 VSS.n13488 0.001
R16152 VSS.n13603 VSS.n13486 0.001
R16153 VSS.n13604 VSS.n13603 0.001
R16154 VSS.n13344 VSS.n13308 0.001
R16155 VSS.n13344 VSS.n13314 0.001
R16156 VSS.n13344 VSS.n13320 0.001
R16157 VSS.n13344 VSS.n13324 0.001
R16158 VSS.n13344 VSS.n13334 0.001
R16159 VSS.n13344 VSS.n13340 0.001
R16160 VSS.n13345 VSS.n13344 0.001
R16161 VSS.n13473 VSS.n13446 0.001
R16162 VSS.n13473 VSS.n13436 0.001
R16163 VSS.n13473 VSS.n13409 0.001
R16164 VSS.n4541 VSS.n4540 0.001
R16165 VSS.n10635 VSS.n10634 0.001
R16166 VSS.n3367 VSS.n3366 0.001
R16167 VSS.n5388 VSS.n5387 0.001
R16168 VSS.n6127 VSS.n6126 0.001
R16169 VSS.n6111 VSS.n6110 0.001
R16170 VSS.n5945 VSS.n5944 0.001
R16171 VSS.n5929 VSS.n5928 0.001
R16172 VSS.n5764 VSS.n5763 0.001
R16173 VSS.n5748 VSS.n5747 0.001
R16174 VSS.n5584 VSS.n5583 0.001
R16175 VSS.n5568 VSS.n5567 0.001
R16176 VSS.n5404 VSS.n5403 0.001
R16177 VSS.n5224 VSS.n5223 0.001
R16178 VSS.n5208 VSS.n5207 0.001
R16179 VSS.n10119 VSS.n10118 0.001
R16180 VSS.n10156 VSS.n10155 0.001
R16181 VSS.n11162 VSS.n11161 0.001
R16182 VSS.n11178 VSS.n11177 0.001
R16183 VSS.n12285 VSS.n12284 0.001
R16184 VSS.n12313 VSS.n12312 0.001
R16185 VSS.n11562 VSS.n11561 0.001
R16186 VSS.n3611 VSS.n3610 0.001
R16187 VSS.n11485 VSS.n11470 0.001
R16188 VSS.n11485 VSS.n11465 0.001
R16189 VSS.n11485 VSS.n11460 0.001
R16190 VSS.n12170 VSS.n12169 0.001
R16191 VSS.n12188 VSS.n12187 0.001
R16192 VSS.n14499 VSS.n14498 0.001
R16193 VSS.n14467 VSS.n14466 0.001
R16194 VSS.n3312 VSS.n3311 0.001
R16195 VSS.n12558 VSS.n12557 0.001
R16196 VSS.n3404 VSS.n3403 0.001
R16197 VSS.n3574 VSS.n3573 0.001
R16198 VSS.n11889 VSS.n11888 0.001
R16199 VSS.n12003 VSS.n12002 0.001
R16200 VSS.n12020 VSS.n12019 0.001
R16201 VSS.n9690 VSS.n9666 0.001
R16202 VSS.n9690 VSS.n9661 0.001
R16203 VSS.n9137 VSS.n9025 0.001
R16204 VSS.n8702 VSS.n8678 0.001
R16205 VSS.n8702 VSS.n8673 0.001
R16206 VSS.n9634 VSS.n7526 0.001
R16207 VSS.n8747 VSS.n8741 0.001
R16208 VSS.n8615 VSS.n8570 0.001
R16209 VSS.n8747 VSS.n8746 0.001
R16210 VSS.n8778 VSS.n8215 0.001
R16211 VSS.n8788 VSS.n8209 0.001
R16212 VSS.n9976 VSS.n6230 0.001
R16213 VSS.n9974 VSS.n6230 0.001
R16214 VSS.n6761 VSS.n6697 0.001
R16215 VSS.n8114 VSS.n8039 0.001
R16216 VSS.n8035 VSS.n8034 0.001
R16217 VSS.n8067 VSS.n7953 0.001
R16218 VSS.n8868 VSS.n7953 0.001
R16219 VSS.n8893 VSS.n7954 0.001
R16220 VSS.n8189 VSS.n8183 0.001
R16221 VSS.n8826 VSS.n8177 0.001
R16222 VSS.n7570 VSS.n7555 0.001
R16223 VSS.n9577 VSS.n7556 0.001
R16224 VSS.n9577 VSS.n7558 0.001
R16225 VSS.n8557 VSS.n8347 0.001
R16226 VSS.n8557 VSS.n8556 0.001
R16227 VSS.n8482 VSS.n8463 0.001
R16228 VSS.n9415 VSS.n9370 0.001
R16229 VSS.n9785 VSS.n7391 0.001
R16230 VSS.n9785 VSS.n7396 0.001
R16231 VSS.n7472 VSS.n7427 0.001
R16232 VSS.n10832 VSS.n3932 0.001
R16233 VSS.n10832 VSS.n3929 0.001
R16234 VSS.n9444 VSS.n9438 0.001
R16235 VSS.n9109 VSS.n9064 0.001
R16236 VSS.n9444 VSS.n9443 0.001
R16237 VSS.n9516 VSS.n8999 0.001
R16238 VSS.n9315 VSS.n9016 0.001
R16239 VSS.n9318 VSS.n9016 0.001
R16240 VSS.n7220 VSS.n7180 0.001
R16241 VSS.n7187 VSS.n7180 0.001
R16242 VSS.n9838 VSS.n7163 0.001
R16243 VSS.n7209 VSS.n7208 0.001
R16244 VSS.n7374 VSS.n7208 0.001
R16245 VSS.n7367 VSS.n7264 0.001
R16246 VSS.n9265 VSS.n9183 0.001
R16247 VSS.n9214 VSS.n9165 0.001
R16248 VSS.n9265 VSS.n9184 0.001
R16249 VSS.n8958 VSS.n7819 0.001
R16250 VSS.n8958 VSS.n7828 0.001
R16251 VSS.n7853 VSS.n7814 0.001
R16252 VSS.n7733 VSS.n7631 0.001
R16253 VSS.n7643 VSS.n7631 0.001
R16254 VSS.n8985 VSS.n7616 0.001
R16255 VSS.n7699 VSS.n7666 0.001
R16256 VSS.n7702 VSS.n7666 0.001
R16257 VSS.n7775 VSS.n7651 0.001
R16258 VSS.n9891 VSS.n7087 0.001
R16259 VSS.n9889 VSS.n7087 0.001
R16260 VSS.n7137 VSS.n7091 0.001
R16261 VSS.n9851 VSS.n7150 0.001
R16262 VSS.n8932 VSS.n7892 0.001
R16263 VSS.n8932 VSS.n8928 0.001
R16264 VSS.n7943 VSS.n7877 0.001
R16265 VSS.n6854 VSS.n6631 0.001
R16266 VSS.n6627 VSS.n6626 0.001
R16267 VSS.n6906 VSS.n6626 0.001
R16268 VSS.n6921 VSS.n6583 0.001
R16269 VSS.n6579 VSS.n6578 0.001
R16270 VSS.n6979 VSS.n6578 0.001
R16271 VSS.n7040 VSS.n6521 0.001
R16272 VSS.n7040 VSS.n6530 0.001
R16273 VSS.n6542 VSS.n6516 0.001
R16274 VSS.n6290 VSS.n6289 0.001
R16275 VSS.n7060 VSS.n6289 0.001
R16276 VSS.n7053 VSS.n6485 0.001
R16277 VSS.n6453 VSS.n6314 0.001
R16278 VSS.n6451 VSS.n6314 0.001
R16279 VSS.n6421 VSS.n6318 0.001
R16280 VSS.n9913 VSS.n9912 0.001
R16281 VSS.n9921 VSS.n9920 0.001
R16282 VSS.n6837 VSS.n6674 0.001
R16283 VSS.n6839 VSS.n6674 0.001
R16284 VSS.n6786 VSS.n6678 0.001
R16285 VSS.n6042 VSS.n5997 0.001
R16286 VSS.n5895 VSS.n5887 0.001
R16287 VSS.n5895 VSS.n5890 0.001
R16288 VSS.n5844 VSS.n5799 0.001
R16289 VSS.n5714 VSS.n5706 0.001
R16290 VSS.n5714 VSS.n5709 0.001
R16291 VSS.n5663 VSS.n5618 0.001
R16292 VSS.n5534 VSS.n5526 0.001
R16293 VSS.n5534 VSS.n5529 0.001
R16294 VSS.n5483 VSS.n5438 0.001
R16295 VSS.n5354 VSS.n5346 0.001
R16296 VSS.n5354 VSS.n5349 0.001
R16297 VSS.n5303 VSS.n5258 0.001
R16298 VSS.n10088 VSS.n10080 0.001
R16299 VSS.n10088 VSS.n10083 0.001
R16300 VSS.n4624 VSS.n4580 0.001
R16301 VSS.n4624 VSS.n4607 0.001
R16302 VSS.n3809 VSS.n3760 0.001
R16303 VSS.n6079 VSS.n6075 0.001
R16304 VSS.n6203 VSS.n6184 0.001
R16305 VSS.n11134 VSS.n3721 0.001
R16306 VSS.n11134 VSS.n11133 0.001
R16307 VSS.n11107 VSS.n11074 0.001
R16308 VSS.n11113 VSS.n3822 0.001
R16309 VSS.n3820 VSS.n3819 0.001
R16310 VSS.n6391 VSS.n3830 0.001
R16311 VSS.n6392 VSS.n3830 0.001
R16312 VSS.n11042 VSS.n3836 0.001
R16313 VSS.n3844 VSS.n3841 0.001
R16314 VSS.n11000 VSS.n3845 0.001
R16315 VSS.n10987 VSS.n3858 0.001
R16316 VSS.n10987 VSS.n10986 0.001
R16317 VSS.n10945 VSS.n3859 0.001
R16318 VSS.n10954 VSS.n3890 0.001
R16319 VSS.n3888 VSS.n3887 0.001
R16320 VSS.n7337 VSS.n3898 0.001
R16321 VSS.n7338 VSS.n3898 0.001
R16322 VSS.n10891 VSS.n3904 0.001
R16323 VSS.n10852 VSS.n10851 0.001
R16324 VSS.n3911 VSS.n3910 0.001
R16325 VSS.n4019 VSS.n3974 0.001
R16326 VSS.n4019 VSS.n4018 0.001
R16327 VSS.n4083 VSS.n4057 0.001
R16328 VSS.n4302 VSS.n4234 0.001
R16329 VSS.n4300 VSS.n4234 0.001
R16330 VSS.n4344 VSS.n4249 0.001
R16331 VSS.n4404 VSS.n4188 0.001
R16332 VSS.n4404 VSS.n4403 0.001
R16333 VSS.n4405 VSS.n4181 0.001
R16334 VSS.n10776 VSS.n4113 0.001
R16335 VSS.n10776 VSS.n10775 0.001
R16336 VSS.n4451 VSS.n4114 0.001
R16337 VSS.n1296 VSS.n1272 0.001
R16338 VSS.n1296 VSS.n1269 0.001
R16339 VSS.n790 VSS.n659 0.001
R16340 VSS.n1345 VSS.n1341 0.001
R16341 VSS.n1047 VSS.n1002 0.001
R16342 VSS.n1345 VSS.n1344 0.001
R16343 VSS.n14275 VSS.n514 0.001
R16344 VSS.n10704 VSS.n10673 0.001
R16345 VSS.n1151 VSS.n915 0.001
R16346 VSS.n603 VSS.n602 0.001
R16347 VSS.n2479 VSS.n2478 0.001
R16348 VSS.n13052 VSS.n2478 0.001
R16349 VSS.n13045 VSS.n2484 0.001
R16350 VSS.n13101 VSS.n2357 0.001
R16351 VSS.n2456 VSS.n2356 0.001
R16352 VSS.n13132 VSS.n1928 0.001
R16353 VSS.n13130 VSS.n1928 0.001
R16354 VSS.n2342 VSS.n1932 0.001
R16355 VSS.n14228 VSS.n570 0.001
R16356 VSS.n14228 VSS.n14227 0.001
R16357 VSS.n14229 VSS.n555 0.001
R16358 VSS.n1165 VSS.n884 0.001
R16359 VSS.n1394 VSS.n879 0.001
R16360 VSS.n880 VSS.n879 0.001
R16361 VSS.n1106 VSS.n960 0.001
R16362 VSS.n1106 VSS.n1105 0.001
R16363 VSS.n14332 VSS.n14306 0.001
R16364 VSS.n1569 VSS.n1524 0.001
R16365 VSS.n13853 VSS.n13716 0.001
R16366 VSS.n13853 VSS.n13719 0.001
R16367 VSS.n13809 VSS.n13764 0.001
R16368 VSS.n13388 VSS.n13256 0.001
R16369 VSS.n13388 VSS.n13251 0.001
R16370 VSS.n1616 VSS.n1612 0.001
R16371 VSS.n762 VSS.n717 0.001
R16372 VSS.n1616 VSS.n1615 0.001
R16373 VSS.n14115 VSS.n633 0.001
R16374 VSS.n1685 VSS.n650 0.001
R16375 VSS.n1464 VSS.n650 0.001
R16376 VSS.n13670 VSS.n1661 0.001
R16377 VSS.n13697 VSS.n1661 0.001
R16378 VSS.n14079 VSS.n1646 0.001
R16379 VSS.n13902 VSS.n13221 0.001
R16380 VSS.n13900 VSS.n13221 0.001
R16381 VSS.n13643 VSS.n13225 0.001
R16382 VSS.n1435 VSS.n836 0.001
R16383 VSS.n843 VSS.n818 0.001
R16384 VSS.n1435 VSS.n837 0.001
R16385 VSS.n2211 VSS.n2005 0.001
R16386 VSS.n2214 VSS.n2005 0.001
R16387 VSS.n2245 VSS.n1988 0.001
R16388 VSS.n2127 VSS.n2080 0.001
R16389 VSS.n2130 VSS.n2080 0.001
R16390 VSS.n2180 VSS.n2063 0.001
R16391 VSS.n1850 VSS.n1849 0.001
R16392 VSS.n13195 VSS.n1849 0.001
R16393 VSS.n13188 VSS.n1855 0.001
R16394 VSS.n12686 VSS.n1777 0.001
R16395 VSS.n13923 VSS.n1777 0.001
R16396 VSS.n13935 VSS.n1778 0.001
R16397 VSS.n14054 VSS.n14053 0.001
R16398 VSS.n2027 VSS.n1972 0.001
R16399 VSS.n1979 VSS.n1972 0.001
R16400 VSS.n2319 VSS.n1953 0.001
R16401 VSS.n12985 VSS.n2567 0.001
R16402 VSS.n2664 VSS.n2584 0.001
R16403 VSS.n2716 VSS.n2584 0.001
R16404 VSS.n12949 VSS.n2673 0.001
R16405 VSS.n2814 VSS.n2688 0.001
R16406 VSS.n2787 VSS.n2688 0.001
R16407 VSS.n12908 VSS.n2748 0.001
R16408 VSS.n2845 VSS.n2765 0.001
R16409 VSS.n2896 VSS.n2765 0.001
R16410 VSS.n3054 VSS.n2868 0.001
R16411 VSS.n12638 VSS.n2868 0.001
R16412 VSS.n12872 VSS.n2853 0.001
R16413 VSS.n3077 VSS.n2955 0.001
R16414 VSS.n12718 VSS.n2955 0.001
R16415 VSS.n12730 VSS.n2956 0.001
R16416 VSS.n13177 VSS.n13176 0.001
R16417 VSS.n2634 VSS.n2524 0.001
R16418 VSS.n2607 VSS.n2524 0.001
R16419 VSS.n13024 VSS.n2505 0.001
R16420 VSS.n11676 VSS.n11576 0.001
R16421 VSS.n12256 VSS.n12248 0.001
R16422 VSS.n12256 VSS.n12251 0.001
R16423 VSS.n11745 VSS.n11700 0.001
R16424 VSS.n12149 VSS.n12141 0.001
R16425 VSS.n12149 VSS.n12144 0.001
R16426 VSS.n12098 VSS.n12053 0.001
R16427 VSS.n11981 VSS.n11973 0.001
R16428 VSS.n11981 VSS.n11976 0.001
R16429 VSS.n11877 VSS.n11832 0.001
R16430 VSS.n3553 VSS.n3545 0.001
R16431 VSS.n3553 VSS.n3548 0.001
R16432 VSS.n3502 VSS.n3457 0.001
R16433 VSS.n12605 VSS.n12597 0.001
R16434 VSS.n12605 VSS.n12600 0.001
R16435 VSS.n3164 VSS.n3120 0.001
R16436 VSS.n3164 VSS.n3141 0.001
R16437 VSS.n3267 VSS.n3222 0.001
R16438 VSS.n11629 VSS.n11625 0.001
R16439 VSS.n12453 VSS.n12389 0.001
R16440 VSS.n12824 VSS.n2927 0.001
R16441 VSS.n12833 VSS.n12832 0.001
R16442 VSS.n2945 VSS.n2935 0.001
R16443 VSS.n12757 VSS.n2935 0.001
R16444 VSS.n12796 VSS.n2941 0.001
R16445 VSS.n1750 VSS.n1748 0.001
R16446 VSS.n13996 VSS.n1751 0.001
R16447 VSS.n13967 VSS.n1720 0.001
R16448 VSS.n13965 VSS.n1720 0.001
R16449 VSS.n14016 VSS.n1735 0.001
R16450 VSS.n14023 VSS.n1712 0.001
R16451 VSS.n14032 VSS.n14031 0.001
R16452 VSS.n13556 VSS.n13485 0.001
R16453 VSS.n13580 VSS.n13485 0.001
R16454 VSS.n13603 VSS.n13500 0.001
R16455 VSS.n13400 VSS.n13399 0.001
R16456 VSS.n13623 VSS.n13622 0.001
R16457 VSS.n13344 VSS.n13301 0.001
R16458 VSS.n13344 VSS.n13343 0.001
R16459 VSS.n13473 VSS.n13454 0.001
R16460 VSS.n3431 VSS 0.000820819
R16461 VSS.n11314 VSS.n11313 0.000801468
R16462 VSS.n6087 VSS.n4671 0.000760417
R16463 VSS.n5905 VSS.n4680 0.000760417
R16464 VSS.n5724 VSS.n4689 0.000760417
R16465 VSS.n5544 VSS.n4700 0.000760417
R16466 VSS.n5364 VSS.n4712 0.000760417
R16467 VSS.n10098 VSS.n4575 0.000760417
R16468 VSS.n3716 VSS.n3715 0.000760417
R16469 VSS.n12342 VSS.n11569 0.000760417
R16470 VSS.n12265 VSS.n11693 0.000760417
R16471 VSS.n12158 VSS.n11779 0.000760417
R16472 VSS.n11990 VSS.n11825 0.000760417
R16473 VSS.n3562 VSS.n3397 0.000760417
R16474 VSS.n12584 VSS.n3117 0.000760417
R16475 VSS.n3289 VSS.n3187 0.000760417
R16476 VSS.n11313 VSS.n11305 0.00073829
R16477 VSS.n11313 VSS.n11312 0.00073829
R16478 VSS.n11312 VSS.n11311 0.00073829
R16479 VSS.n4817 VSS.n4811 0.000712971
R16480 VSS.n4819 VSS.n4818 0.000712971
R16481 VSS.n4927 VSS.n4926 0.000712971
R16482 VSS.n4925 VSS.n4824 0.000712971
R16483 VSS.n4914 VSS.n4860 0.000712971
R16484 VSS.n4913 VSS.n4861 0.000712971
R16485 VSS.n4948 VSS.n4947 0.000712971
R16486 VSS.n5095 VSS.n5094 0.000712971
R16487 VSS.n4816 VSS.n4812 0.000712971
R16488 VSS.n4815 VSS.n4814 0.000712971
R16489 VSS.n4944 VSS.n4943 0.000712971
R16490 VSS.n4946 VSS.n4945 0.000712971
R16491 VSS.n4935 VSS.n4821 0.000712971
R16492 VSS.n4934 VSS.n4822 0.000712971
R16493 VSS.n4923 VSS.n4834 0.000712971
R16494 VSS.n4922 VSS.n4835 0.000712971
R16495 VSS.n4920 VSS.n4841 0.000712971
R16496 VSS.n4919 VSS.n4842 0.000712971
R16497 VSS.n4917 VSS.n4852 0.000712971
R16498 VSS.n4916 VSS.n4853 0.000712971
R16499 VSS.n4911 VSS.n4862 0.000712971
R16500 VSS.n4910 VSS.n4863 0.000712971
R16501 VSS.n10177 VSS.n10176 0.000712971
R16502 VSS.n10176 VSS.n4552 0.000712971
R16503 VSS.n5098 VSS.n5097 0.000712971
R16504 VSS.n5100 VSS.n5099 0.000712971
R16505 VSS.n5107 VSS.n5106 0.000712971
R16506 VSS.n5109 VSS.n5108 0.000712971
R16507 VSS.n12483 VSS.n12482 0.000712971
R16508 VSS.n12482 VSS.n12481 0.000712971
R16509 VSS.n5155 VSS.n5154 0.000712971
R16510 VSS.n10413 VSS.n10410 0.000712971
R16511 VSS.n10412 VSS.n10411 0.000712971
R16512 VSS.n10507 VSS.n10506 0.000712971
R16513 VSS.n10509 VSS.n10508 0.000712971
R16514 VSS.n10513 VSS.n10253 0.000712971
R16515 VSS.n10515 VSS.n10514 0.000712971
R16516 VSS.n10520 VSS.n10519 0.000712971
R16517 VSS.n10523 VSS.n10522 0.000712971
R16518 VSS.n10532 VSS.n10524 0.000712971
R16519 VSS.n10531 VSS.n10530 0.000712971
R16520 VSS.n12549 VSS.n12548 0.000712971
R16521 VSS.n10424 VSS.n10396 0.000712971
R16522 VSS.n10425 VSS.n10395 0.000712971
R16523 VSS.n10389 VSS.n10388 0.000712971
R16524 VSS.n10386 VSS.n10385 0.000712971
R16525 VSS.n10378 VSS.n10377 0.000712971
R16526 VSS.n10376 VSS.n10375 0.000712971
R16527 VSS.n10381 VSS.n10380 0.000712971
R16528 VSS.n10383 VSS.n10382 0.000712971
R16529 VSS.n10391 VSS.n10272 0.000712971
R16530 VSS.n10393 VSS.n10392 0.000712971
R16531 VSS.n10422 VSS.n10401 0.000712971
R16532 VSS.n10421 VSS.n10402 0.000712971
R16533 VSS.n10418 VSS.n10404 0.000712971
R16534 VSS.n10417 VSS.n10405 0.000712971
R16535 VSS.n10415 VSS.n10408 0.000712971
R16536 VSS.n10414 VSS.n10409 0.000712971
R16537 VSS.n10200 VSS.n10199 0.000712971
R16538 VSS.n10197 VSS.n4550 0.000712971
R16539 VSS.n10192 VSS.n3683 0.000712971
R16540 VSS.n10194 VSS.n10193 0.000712971
R16541 VSS.n10198 VSS.n4549 0.000712971
R16542 VSS.n4905 VSS.n4548 0.000712971
R16543 VSS.n4906 VSS.n4864 0.000712971
R16544 VSS.n4908 VSS.n4907 0.000712971
R16545 VSS.n12491 VSS.n3602 0.000712971
R16546 VSS.n12490 VSS.n3602 0.000712971
R16547 VSS.n10596 VSS.n10594 0.000712971
R16548 VSS.n10593 VSS.n3680 0.000712971
R16549 VSS.n10374 VSS.n10372 0.000712971
R16550 VSS.n10373 VSS.n10204 0.000712971
R16551 VSS.n11443 VSS.n11442 0.000712971
R16552 VSS.n11445 VSS.n11444 0.000712971
R16553 VSS.n10600 VSS.n10599 0.000712971
R16554 VSS.n10371 VSS.n4543 0.000712971
R16555 VSS.n11432 VSS.n3682 0.000712971
R16556 VSS.n11431 VSS.n11430 0.000712971
R16557 VSS.n11452 VSS.n11451 0.000712971
R16558 VSS.n11450 VSS.n3677 0.000712971
R16559 VSS.n11449 VSS.n11448 0.000712971
R16560 VSS.n3681 VSS.n3678 0.000712971
R16561 VSS.n11439 VSS.n11438 0.000712971
R16562 VSS.n10595 VSS.n10203 0.000712971
R16563 VSS.n10604 VSS.n4547 0.000712971
R16564 VSS.n10605 VSS.n4546 0.000712971
R16565 VSS.n10793 VSS.n10791 0.000684314
R16566 VSS.n10800 VSS.n10797 0.000684314
R16567 VSS.n10789 VSS.n4103 0.000684314
R16568 VSS.n10738 VSS.n10736 0.000684314
R16569 VSS.n10645 VSS.n10642 0.000684314
R16570 VSS.n10740 VSS.n4456 0.000684314
R16571 VSS.n12160 VSS.n11778 0.000672891
R16572 VSS.n3206 VSS 0.00066041
R16573 VSS.n3353 VSS 0.00066041
R16574 VSS.n11916 VSS 0.00066041
R16575 VSS.n11772 VSS 0.00066041
R16576 VSS.n11547 VSS 0.00066041
R16577 VSS.n4940 VSS.n4801 0.000606486
R16578 VSS.n4941 VSS.n4809 0.000606486
R16579 VSS.n4951 VSS.n4950 0.000606486
R16580 VSS.n4954 VSS.n4953 0.000606486
R16581 VSS.n4805 VSS.n4804 0.000606486
R16582 VSS.n4962 VSS.n4961 0.000606486
R16583 VSS.n4830 VSS.n4784 0.000606486
R16584 VSS.n4829 VSS.n4828 0.000606486
R16585 VSS.n4964 VSS.n4963 0.000606486
R16586 VSS.n5017 VSS.n5016 0.000606486
R16587 VSS.n4975 VSS.n4974 0.000606486
R16588 VSS.n4972 VSS.n4971 0.000606486
R16589 VSS.n5014 VSS.n5013 0.000606486
R16590 VSS.n5023 VSS.n5022 0.000606486
R16591 VSS.n4894 VSS.n4893 0.000606486
R16592 VSS.n4892 VSS.n4891 0.000606486
R16593 VSS.n5056 VSS.n5055 0.000606486
R16594 VSS.n5054 VSS.n5053 0.000606486
R16595 VSS.n4848 VSS.n4776 0.000606486
R16596 VSS.n4847 VSS.n4846 0.000606486
R16597 VSS.n5025 VSS.n5024 0.000606486
R16598 VSS.n5036 VSS.n5035 0.000606486
R16599 VSS.n5033 VSS.n5032 0.000606486
R16600 VSS.n5048 VSS.n5047 0.000606486
R16601 VSS.n5045 VSS.n5043 0.000606486
R16602 VSS.n4869 VSS.n4773 0.000606486
R16603 VSS.n4872 VSS.n4871 0.000606486
R16604 VSS.n4878 VSS.n4877 0.000606486
R16605 VSS.n4875 VSS.n4874 0.000606486
R16606 VSS.n4900 VSS.n4899 0.000606486
R16607 VSS.n4904 VSS.n4903 0.000606486
R16608 VSS.n4873 VSS.n4551 0.000606486
R16609 VSS.n10191 VSS.n3684 0.000606486
R16610 VSS.n10190 VSS.n10189 0.000606486
R16611 VSS.n10178 VSS.n4560 0.000606486
R16612 VSS.n10180 VSS.n4559 0.000606486
R16613 VSS.n4897 VSS.n4896 0.000606486
R16614 VSS.n4889 VSS.n4888 0.000606486
R16615 VSS.n10184 VSS.n4556 0.000606486
R16616 VSS.n10182 VSS.n4557 0.000606486
R16617 VSS.n4882 VSS.n4879 0.000606486
R16618 VSS.n4881 VSS.n4880 0.000606486
R16619 VSS.n4885 VSS.n4865 0.000606486
R16620 VSS.n4884 VSS.n4866 0.000606486
R16621 VSS.n10165 VSS.n10164 0.000606486
R16622 VSS.n4724 VSS.n4723 0.000606486
R16623 VSS.n4725 VSS.n4721 0.000606486
R16624 VSS.n5068 VSS.n4763 0.000606486
R16625 VSS.n10187 VSS.n10186 0.000606486
R16626 VSS.n4770 VSS.n4555 0.000606486
R16627 VSS.n4856 VSS.n4855 0.000606486
R16628 VSS.n4858 VSS.n4854 0.000606486
R16629 VSS.n5173 VSS.n5172 0.000606486
R16630 VSS.n4768 VSS.n4765 0.000606486
R16631 VSS.n4767 VSS.n4766 0.000606486
R16632 VSS.n5064 VSS.n5063 0.000606486
R16633 VSS.n5066 VSS.n5065 0.000606486
R16634 VSS.n5059 VSS.n5058 0.000606486
R16635 VSS.n5061 VSS.n5060 0.000606486
R16636 VSS.n5170 VSS.n5169 0.000606486
R16637 VSS.n5168 VSS.n5167 0.000606486
R16638 VSS.n4849 VSS.n4777 0.000606486
R16639 VSS.n4850 VSS.n4843 0.000606486
R16640 VSS.n4762 VSS.n4728 0.000606486
R16641 VSS.n5165 VSS.n5164 0.000606486
R16642 VSS.n5041 VSS.n5037 0.000606486
R16643 VSS.n5040 VSS.n5039 0.000606486
R16644 VSS.n5051 VSS.n4778 0.000606486
R16645 VSS.n5050 VSS.n4779 0.000606486
R16646 VSS.n5162 VSS.n5161 0.000606486
R16647 VSS.n4987 VSS.n4729 0.000606486
R16648 VSS.n4988 VSS.n4986 0.000606486
R16649 VSS.n5076 VSS.n4756 0.000606486
R16650 VSS.n5071 VSS.n4761 0.000606486
R16651 VSS.n5073 VSS.n4760 0.000606486
R16652 VSS.n4838 VSS.n4837 0.000606486
R16653 VSS.n4839 VSS.n4836 0.000606486
R16654 VSS.n4984 VSS.n4733 0.000606486
R16655 VSS.n4996 VSS.n4995 0.000606486
R16656 VSS.n4999 VSS.n4998 0.000606486
R16657 VSS.n4992 VSS.n4991 0.000606486
R16658 VSS.n4993 VSS.n4759 0.000606486
R16659 VSS.n5029 VSS.n5028 0.000606486
R16660 VSS.n5030 VSS.n4781 0.000606486
R16661 VSS.n5000 VSS.n4983 0.000606486
R16662 VSS.n5001 VSS.n4982 0.000606486
R16663 VSS.n5019 VSS.n4787 0.000606486
R16664 VSS.n5020 VSS.n4786 0.000606486
R16665 VSS.n4832 VSS.n4825 0.000606486
R16666 VSS.n4831 VSS.n4785 0.000606486
R16667 VSS.n5007 VSS.n4755 0.000606486
R16668 VSS.n5006 VSS.n4977 0.000606486
R16669 VSS.n5011 VSS.n4976 0.000606486
R16670 VSS.n5010 VSS.n5009 0.000606486
R16671 VSS.n4980 VSS.n4736 0.000606486
R16672 VSS.n5004 VSS.n5003 0.000606486
R16673 VSS.n4979 VSS.n4978 0.000606486
R16674 VSS.n5083 VSS.n4750 0.000606486
R16675 VSS.n5079 VSS.n4754 0.000606486
R16676 VSS.n5081 VSS.n4753 0.000606486
R16677 VSS.n4793 VSS.n4752 0.000606486
R16678 VSS.n4796 VSS.n4794 0.000606486
R16679 VSS.n4968 VSS.n4967 0.000606486
R16680 VSS.n4969 VSS.n4798 0.000606486
R16681 VSS.n4930 VSS.n4929 0.000606486
R16682 VSS.n4932 VSS.n4928 0.000606486
R16683 VSS.n4791 VSS.n4788 0.000606486
R16684 VSS.n4790 VSS.n4789 0.000606486
R16685 VSS.n5133 VSS.n5132 0.000606486
R16686 VSS.n5092 VSS.n4746 0.000606486
R16687 VSS.n5130 VSS.n5129 0.000606486
R16688 VSS.n5128 VSS.n5127 0.000606486
R16689 VSS.n5125 VSS.n5124 0.000606486
R16690 VSS.n5086 VSS.n4742 0.000606486
R16691 VSS.n4955 VSS.n4748 0.000606486
R16692 VSS.n5089 VSS.n5088 0.000606486
R16693 VSS.n4958 VSS.n4957 0.000606486
R16694 VSS.n4959 VSS.n4803 0.000606486
R16695 VSS.n4938 VSS.n4937 0.000606486
R16696 VSS.n4939 VSS.n4802 0.000606486
R16697 VSS.n5122 VSS.n5121 0.000606486
R16698 VSS.n5103 VSS.n4743 0.000606486
R16699 VSS.n5104 VSS.n5102 0.000606486
R16700 VSS.n5120 VSS.n4744 0.000606486
R16701 VSS.n5137 VSS.n5136 0.000606486
R16702 VSS.n5144 VSS.n5143 0.000606486
R16703 VSS.n5151 VSS.n5150 0.000606486
R16704 VSS.n5160 VSS.n4730 0.000606486
R16705 VSS.n5174 VSS.n4719 0.000606486
R16706 VSS.n10168 VSS.n10167 0.000606486
R16707 VSS.n10363 VSS.n10362 0.000606486
R16708 VSS.n10281 VSS.n10280 0.000606486
R16709 VSS.n12495 VSS.n3599 0.000606486
R16710 VSS.n12494 VSS.n12493 0.000606486
R16711 VSS.n10358 VSS.n10357 0.000606486
R16712 VSS.n10588 VSS.n10209 0.000606486
R16713 VSS.n10586 VSS.n10210 0.000606486
R16714 VSS.n10584 VSS.n10213 0.000606486
R16715 VSS.n10582 VSS.n10214 0.000606486
R16716 VSS.n10580 VSS.n10217 0.000606486
R16717 VSS.n10578 VSS.n10218 0.000606486
R16718 VSS.n10432 VSS.n10431 0.000606486
R16719 VSS.n10460 VSS.n10257 0.000606486
R16720 VSS.n10461 VSS.n10264 0.000606486
R16721 VSS.n10459 VSS.n10263 0.000606486
R16722 VSS.n10458 VSS.n10457 0.000606486
R16723 VSS.n10433 VSS.n10268 0.000606486
R16724 VSS.n10438 VSS.n10437 0.000606486
R16725 VSS.n10442 VSS.n10441 0.000606486
R16726 VSS.n10440 VSS.n10439 0.000606486
R16727 VSS.n10574 VSS.n10573 0.000606486
R16728 VSS.n10571 VSS.n10570 0.000606486
R16729 VSS.n10297 VSS.n10224 0.000606486
R16730 VSS.n10299 VSS.n10298 0.000606486
R16731 VSS.n10356 VSS.n10282 0.000606486
R16732 VSS.n10479 VSS.n10478 0.000606486
R16733 VSS.n10483 VSS.n10482 0.000606486
R16734 VSS.n10485 VSS.n10484 0.000606486
R16735 VSS.n10252 VSS.n10251 0.000606486
R16736 VSS.n10339 VSS.n10319 0.000606486
R16737 VSS.n10566 VSS.n10227 0.000606486
R16738 VSS.n10568 VSS.n10567 0.000606486
R16739 VSS.n10295 VSS.n10294 0.000606486
R16740 VSS.n10296 VSS.n10225 0.000606486
R16741 VSS.n10292 VSS.n10216 0.000606486
R16742 VSS.n10291 VSS.n10273 0.000606486
R16743 VSS.n10345 VSS.n10313 0.000606486
R16744 VSS.n10344 VSS.n10314 0.000606486
R16745 VSS.n10562 VSS.n10230 0.000606486
R16746 VSS.n10564 VSS.n10229 0.000606486
R16747 VSS.n10558 VSS.n10234 0.000606486
R16748 VSS.n10560 VSS.n10233 0.000606486
R16749 VSS.n10575 VSS.n10220 0.000606486
R16750 VSS.n10576 VSS.n10219 0.000606486
R16751 VSS.n10427 VSS.n10271 0.000606486
R16752 VSS.n10429 VSS.n10428 0.000606486
R16753 VSS.n10334 VSS.n10331 0.000606486
R16754 VSS.n10330 VSS.n10329 0.000606486
R16755 VSS.n10337 VSS.n10336 0.000606486
R16756 VSS.n10326 VSS.n10325 0.000606486
R16757 VSS.n10327 VSS.n10232 0.000606486
R16758 VSS.n12536 VSS.n12535 0.000606486
R16759 VSS.n10323 VSS.n10322 0.000606486
R16760 VSS.n12542 VSS.n12541 0.000606486
R16761 VSS.n12540 VSS.n12539 0.000606486
R16762 VSS.n10398 VSS.n10269 0.000606486
R16763 VSS.n10399 VSS.n10397 0.000606486
R16764 VSS.n12533 VSS.n3377 0.000606486
R16765 VSS.n10446 VSS.n10445 0.000606486
R16766 VSS.n10444 VSS.n3378 0.000606486
R16767 VSS.n10450 VSS.n10449 0.000606486
R16768 VSS.n10448 VSS.n10236 0.000606486
R16769 VSS.n10455 VSS.n10435 0.000606486
R16770 VSS.n10454 VSS.n10453 0.000606486
R16771 VSS.n10554 VSS.n10238 0.000606486
R16772 VSS.n10556 VSS.n10237 0.000606486
R16773 VSS.n10550 VSS.n10241 0.000606486
R16774 VSS.n10551 VSS.n10240 0.000606486
R16775 VSS.n10464 VSS.n10463 0.000606486
R16776 VSS.n10419 VSS.n10265 0.000606486
R16777 VSS.n12545 VSS.n12544 0.000606486
R16778 VSS.n10473 VSS.n10239 0.000606486
R16779 VSS.n10472 VSS.n10471 0.000606486
R16780 VSS.n10476 VSS.n10261 0.000606486
R16781 VSS.n10475 VSS.n10470 0.000606486
R16782 VSS.n10467 VSS.n10466 0.000606486
R16783 VSS.n10469 VSS.n10468 0.000606486
R16784 VSS.n10248 VSS.n10247 0.000606486
R16785 VSS.n10246 VSS.n10245 0.000606486
R16786 VSS.n10534 VSS.n10249 0.000606486
R16787 VSS.n10543 VSS.n10536 0.000606486
R16788 VSS.n10548 VSS.n10243 0.000606486
R16789 VSS.n10546 VSS.n10244 0.000606486
R16790 VSS.n10491 VSS.n10487 0.000606486
R16791 VSS.n10490 VSS.n10489 0.000606486
R16792 VSS.n10497 VSS.n10496 0.000606486
R16793 VSS.n10495 VSS.n10259 0.000606486
R16794 VSS.n10502 VSS.n10255 0.000606486
R16795 VSS.n10500 VSS.n10499 0.000606486
R16796 VSS.n10406 VSS.n10256 0.000606486
R16797 VSS.n10504 VSS.n10503 0.000606486
R16798 VSS.n10512 VSS.n10511 0.000606486
R16799 VSS.n10518 VSS.n10517 0.000606486
R16800 VSS.n10533 VSS.n10250 0.000606486
R16801 VSS.n10542 VSS.n10537 0.000606486
R16802 VSS.n12546 VSS.n3321 0.000606486
R16803 VSS.n12532 VSS.n3379 0.000606486
R16804 VSS.n10333 VSS.n3587 0.000606486
R16805 VSS.n12520 VSS.n12519 0.000606486
R16806 VSS.n10317 VSS.n3591 0.000606486
R16807 VSS.n10342 VSS.n10341 0.000606486
R16808 VSS.n10316 VSS.n10315 0.000606486
R16809 VSS.n10303 VSS.n3600 0.000606486
R16810 VSS.n10350 VSS.n10312 0.000606486
R16811 VSS.n10348 VSS.n10347 0.000606486
R16812 VSS.n10308 VSS.n10307 0.000606486
R16813 VSS.n10310 VSS.n10309 0.000606486
R16814 VSS.n10354 VSS.n10301 0.000606486
R16815 VSS.n10352 VSS.n10302 0.000606486
R16816 VSS.n10289 VSS.n10288 0.000606486
R16817 VSS.n10287 VSS.n10286 0.000606486
R16818 VSS.n10283 VSS.n10275 0.000606486
R16819 VSS.n10284 VSS.n10212 0.000606486
R16820 VSS.n12510 VSS.n12509 0.000606486
R16821 VSS.n12513 VSS.n12512 0.000606486
R16822 VSS.n12486 VSS.n12485 0.000606486
R16823 VSS.n12488 VSS.n12484 0.000606486
R16824 VSS.n12505 VSS.n12504 0.000606486
R16825 VSS.n12507 VSS.n12506 0.000606486
R16826 VSS.n12307 VSS.n12306 0.000606486
R16827 VSS.n12301 VSS.n12300 0.000606486
R16828 VSS.n12500 VSS.n12499 0.000606486
R16829 VSS.n12502 VSS.n12501 0.000606486
R16830 VSS.n12497 VSS.n12496 0.000606486
R16831 VSS.n10360 VSS.n10359 0.000606486
R16832 VSS.n10366 VSS.n10365 0.000606486
R16833 VSS.n10364 VSS.n10277 0.000606486
R16834 VSS.n10368 VSS.n10208 0.000606486
R16835 VSS.n10370 VSS.n10369 0.000606486
R16836 VSS.n10591 VSS.n10205 0.000606486
R16837 VSS.n10590 VSS.n10206 0.000606486
R16838 VSS.n11435 VSS.n11434 0.000606486
R16839 VSS.n11437 VSS.n11436 0.000606486
R16840 VSS.n10601 VSS.n10202 0.000606486
R16841 VSS.n10602 VSS.n10201 0.000606486
R16842 VSS.n11290 VSS.n11289 0.000594191
R16843 VSS.n11294 VSS.n11291 0.000593164
R16844 VSS.n11493 VSS.n11492 0.000578781
R16845 VSS.n11492 VSS.n11491 0.000578781
R16846 VSS.n11284 VSS.n11283 0.000578781
R16847 VSS.n11283 VSS.n11282 0.000578781
R16848 VSS.n11287 VSS.n11286 0.000560257
R16849 VSS.n11286 VSS.n11285 0.000560257
R16850 VSS.n11484 VSS.n11483 0.000539391
R16851 VSS.n11485 VSS.n11484 0.000539391
R16852 VSS.n11457 VSS.n11456 0.000539391
R16853 VSS.n11459 VSS.n11458 0.000539391
R16854 VSS.n11462 VSS.n11461 0.000539391
R16855 VSS.n11469 VSS.n11468 0.000539391
R16856 VSS.n11467 VSS.n11466 0.000539391
R16857 VSS.n11464 VSS.n11463 0.000539391
R16858 VSS.n11472 VSS.n11471 0.000539391
R16859 VSS.n11474 VSS.n11473 0.000539391
R16860 VSS.n11227 VSS.n11226 0.000539391
R16861 VSS.n11226 VSS.n11225 0.000539391
R16862 VSS.n11230 VSS.n11229 0.000539391
R16863 VSS.n11229 VSS.n11228 0.000539391
R16864 VSS.n11224 VSS.n11223 0.000539391
R16865 VSS.n11223 VSS.n11222 0.000539391
R16866 VSS.n11221 VSS.n11220 0.000539391
R16867 VSS.n11210 VSS.n11209 0.000539391
R16868 VSS.n11205 VSS.n11204 0.000539391
R16869 VSS.n11207 VSS.n11206 0.000539391
R16870 VSS.n11263 VSS.n11262 0.000539391
R16871 VSS.n11262 VSS.n11261 0.000539391
R16872 VSS.n11265 VSS.n11264 0.000539391
R16873 VSS.n11267 VSS.n11266 0.000539391
R16874 VSS.n11270 VSS.n11269 0.000539391
R16875 VSS.n11272 VSS.n11271 0.000539391
R16876 VSS.n11203 VSS.n11202 0.000539391
R16877 VSS.n11202 VSS.n11201 0.000539391
R16878 VSS.n11301 VSS.n11300 0.000539391
R16879 VSS.n11300 VSS.n11299 0.000539391
R16880 VSS.n11298 VSS.n11297 0.000539391
R16881 VSS.n11297 VSS.n11296 0.000539391
R16882 VSS.n3633 VSS.n3632 0.000539391
R16883 VSS.n3632 VSS.n3631 0.000539391
R16884 VSS.n3636 VSS.n3635 0.000539391
R16885 VSS.n3635 VSS.n3634 0.000539391
R16886 VSS.n11482 VSS.n11481 0.000539391
R16887 VSS.n11481 VSS.n11480 0.000539391
R16888 VSS.n11420 VSS.n11419 0.000539391
R16889 VSS.n11417 VSS.n11416 0.000539391
R16890 VSS.n11455 VSS.n11454 0.000539391
R16891 VSS.n11454 VSS.n11453 0.000539391
R16892 VSS.n11424 VSS.n11423 0.000539391
R16893 VSS.n11423 VSS.n11422 0.000539391
R16894 VSS.n11426 VSS.n11425 0.000539391
R16895 VSS.n11427 VSS.n11426 0.000539391
R16896 VSS.n14374 VSS.n507 0.000533349
R16897 VSS.n10726 VSS.n10725 0.000533349
R16898 VSS.n14374 VSS.n14373 0.000533349
R16899 VSS.n10729 VSS.n10650 0.000533349
R16900 VSS.n10732 VSS.n10729 0.000533349
R16901 VSS.n10802 VSS.n4099 0.000533349
R16902 VSS.n8420 VSS.n8419 0.000533349
R16903 VSS.n8638 VSS.n8335 0.000533349
R16904 VSS.n8638 VSS.n8637 0.000533349
R16905 VSS.n8723 VSS.n8328 0.000533349
R16906 VSS.n8724 VSS.n8723 0.000533349
R16907 VSS.n9713 VSS.n7512 0.000533349
R16908 VSS.n9713 VSS.n9712 0.000533349
R16909 VSS.n9730 VSS.n7505 0.000533349
R16910 VSS.n9730 VSS.n9729 0.000533349
R16911 VSS.n9746 VSS.n9745 0.000533349
R16912 VSS.n9746 VSS.n7493 0.000533349
R16913 VSS.n9757 VSS.n9756 0.000533349
R16914 VSS.n10812 VSS.n3963 0.000533349
R16915 VSS.n10813 VSS.n10812 0.000533349
R16916 VSS.n10808 VSS.n10807 0.000533349
R16917 VSS.n10808 VSS.n4031 0.000533349
R16918 VSS.n9765 VSS.n9764 0.000533349
R16919 VSS.n9766 VSS.n9765 0.000533349
R16920 VSS.n9753 VSS.n9752 0.000533349
R16921 VSS.n9753 VSS.n7491 0.000533349
R16922 VSS.n9737 VSS.n9736 0.000533349
R16923 VSS.n9737 VSS.n7495 0.000533349
R16924 VSS.n9720 VSS.n9719 0.000533349
R16925 VSS.n9720 VSS.n7507 0.000533349
R16926 VSS.n8719 VSS.n8718 0.000533349
R16927 VSS.n8719 VSS.n8714 0.000533349
R16928 VSS.n8645 VSS.n8644 0.000533349
R16929 VSS.n8645 VSS.n8330 0.000533349
R16930 VSS.n14339 VSS.n14338 0.000533349
R16931 VSS.n984 VSS.n983 0.000533349
R16932 VSS.n1239 VSS.n1236 0.000533349
R16933 VSS.n1068 VSS.n1053 0.000533349
R16934 VSS.n1241 VSS.n1239 0.000533349
R16935 VSS.n1241 VSS.n1240 0.000533349
R16936 VSS.n1068 VSS.n1067 0.000533349
R16937 VSS.n13751 VSS.n13748 0.000533349
R16938 VSS.n1590 VSS.n1575 0.000533349
R16939 VSS.n13752 VSS.n13751 0.000533349
R16940 VSS.n1590 VSS.n1589 0.000533349
R16941 VSS.n13289 VSS.n13286 0.000533349
R16942 VSS.n13830 VSS.n13815 0.000533349
R16943 VSS.n13830 VSS.n13829 0.000533349
R16944 VSS.n13290 VSS.n13289 0.000533349
R16945 VSS.n13421 VSS.n13416 0.000533349
R16946 VSS.n13422 VSS.n13421 0.000533349
R16947 VSS.n456 VSS.n455 0.000533349
R16948 VSS.n1505 VSS.n1504 0.000533349
R16949 VSS.n703 VSS.n702 0.000533349
R16950 VSS.n1303 VSS.n1302 0.000533349
R16951 VSS.n3441 VSS.n3440 0.000533349
R16952 VSS.n11926 VSS.n11925 0.000533349
R16953 VSS.n12039 VSS.n12038 0.000533349
R16954 VSS.n12203 VSS.n12202 0.000533349
R16955 VSS.n14504 VSS.n14503 0.000533349
R16956 VSS.n12467 VSS.n12466 0.000533349
R16957 VSS.n3360 VSS.n3354 0.000533349
R16958 VSS.n3567 VSS.n3394 0.000533349
R16959 VSS.n11996 VSS.n11823 0.000533349
R16960 VSS.n11689 VSS.n11688 0.000533349
R16961 VSS.n12351 VSS.n12350 0.000533349
R16962 VSS.n12336 VSS.n12327 0.000533349
R16963 VSS.n12574 VSS.n12573 0.000533349
R16964 VSS.n12574 VSS.n3176 0.000533349
R16965 VSS.n11515 VSS.n11514 0.000533349
R16966 VSS.n11524 VSS.n11515 0.000533349
R16967 VSS.n10130 VSS.n3708 0.000533349
R16968 VSS.n11149 VSS.n3708 0.000533349
R16969 VSS.n6142 VSS.n6141 0.000533349
R16970 VSS.n10149 VSS.n10143 0.000533349
R16971 VSS.n5201 VSS.n5195 0.000533349
R16972 VSS.n5381 VSS.n5375 0.000533349
R16973 VSS.n5561 VSS.n5555 0.000533349
R16974 VSS.n5741 VSS.n5735 0.000533349
R16975 VSS.n5922 VSS.n5916 0.000533349
R16976 VSS.n6104 VSS.n6098 0.000533349
R16977 VSS.n5959 VSS.n5958 0.000533349
R16978 VSS.n5778 VSS.n5777 0.000533349
R16979 VSS.n4692 VSS.n4686 0.000533349
R16980 VSS.n5597 VSS.n4692 0.000533349
R16981 VSS.n4703 VSS.n4697 0.000533349
R16982 VSS.n5417 VSS.n4703 0.000533349
R16983 VSS.n4715 VSS.n4709 0.000533349
R16984 VSS.n5237 VSS.n4715 0.000533349
R16985 VSS.n5183 VSS.n4566 0.000533349
R16986 VSS.n10106 VSS.n4566 0.000533349
R16987 VSS.n11192 VSS.n11191 0.000533349
R16988 VSS.n10739 VSS.n10645 0.000516685
R16989 VSS.n10740 VSS.n10739 0.000516685
R16990 VSS.n10801 VSS.n10800 0.000516685
R16991 VSS.n10797 VSS.n10794 0.000516685
R16992 VSS.n10794 VSS.n10789 0.000516685
R16993 VSS.n10794 VSS.n10793 0.000516685
R16994 VSS.n10642 VSS.n10639 0.000516685
R16995 VSS.n10739 VSS.n10738 0.000516685
R16996 VSS.n11294 VSS.n11293 0.000516018
R16997 VSS.n11313 VSS.n11295 0.000516018
R16998 VSS.n11500 VSS.n11495 0.000513139
R16999 VSS.n10638 VSS.n10637 0.000511116
R17000 VSS.n10619 VSS.n10618 0.000511116
R17001 VSS.n10613 VSS.n10612 0.000511116
R17002 VSS.n10611 VSS.n10610 0.000511116
R17003 VSS.n4538 VSS.n4537 0.000511116
R17004 VSS.n6124 VSS.n6123 0.000511116
R17005 VSS.n6122 VSS.n6121 0.000511116
R17006 VSS.n6108 VSS.n6107 0.000511116
R17007 VSS.n5956 VSS.n5955 0.000511116
R17008 VSS.n5942 VSS.n5941 0.000511116
R17009 VSS.n5940 VSS.n5939 0.000511116
R17010 VSS.n5926 VSS.n5925 0.000511116
R17011 VSS.n5775 VSS.n5774 0.000511116
R17012 VSS.n5761 VSS.n5760 0.000511116
R17013 VSS.n5759 VSS.n5758 0.000511116
R17014 VSS.n5745 VSS.n5744 0.000511116
R17015 VSS.n5595 VSS.n5594 0.000511116
R17016 VSS.n5581 VSS.n5580 0.000511116
R17017 VSS.n5579 VSS.n5578 0.000511116
R17018 VSS.n5565 VSS.n5564 0.000511116
R17019 VSS.n5415 VSS.n5414 0.000511116
R17020 VSS.n5401 VSS.n5400 0.000511116
R17021 VSS.n5399 VSS.n5398 0.000511116
R17022 VSS.n5385 VSS.n5384 0.000511116
R17023 VSS.n5235 VSS.n5234 0.000511116
R17024 VSS.n5221 VSS.n5220 0.000511116
R17025 VSS.n5219 VSS.n5218 0.000511116
R17026 VSS.n5205 VSS.n5204 0.000511116
R17027 VSS.n10108 VSS.n10107 0.000511116
R17028 VSS.n10122 VSS.n10121 0.000511116
R17029 VSS.n10124 VSS.n10123 0.000511116
R17030 VSS.n10153 VSS.n10152 0.000511116
R17031 VSS.n11151 VSS.n11150 0.000511116
R17032 VSS.n11165 VSS.n11164 0.000511116
R17033 VSS.n11167 VSS.n11166 0.000511116
R17034 VSS.n11181 VSS.n11180 0.000511116
R17035 VSS.n3193 VSS.n3192 0.000511116
R17036 VSS.n3208 VSS.n3207 0.000511116
R17037 VSS.n12472 VSS.n12471 0.000511116
R17038 VSS.n11565 VSS.n11564 0.000511116
R17039 VSS.n11556 VSS.n11555 0.000511116
R17040 VSS.n3309 VSS.n3308 0.000511116
R17041 VSS.n3314 VSS.n3313 0.000511116
R17042 VSS.n12555 VSS.n12554 0.000511116
R17043 VSS.n12570 VSS.n12569 0.000511116
R17044 VSS.n3364 VSS.n3363 0.000511116
R17045 VSS.n3369 VSS.n3368 0.000511116
R17046 VSS.n3401 VSS.n3400 0.000511116
R17047 VSS.n3417 VSS.n3416 0.000511116
R17048 VSS.n3571 VSS.n3570 0.000511116
R17049 VSS.n3581 VSS.n3580 0.000511116
R17050 VSS.n11886 VSS.n11885 0.000511116
R17051 VSS.n11902 VSS.n11901 0.000511116
R17052 VSS.n12000 VSS.n11999 0.000511116
R17053 VSS.n12015 VSS.n12014 0.000511116
R17054 VSS.n12017 VSS.n12016 0.000511116
R17055 VSS.n12031 VSS.n12030 0.000511116
R17056 VSS.n12167 VSS.n12166 0.000511116
R17057 VSS.n12183 VSS.n12182 0.000511116
R17058 VSS.n12185 VSS.n12184 0.000511116
R17059 VSS.n12201 VSS.n12200 0.000511116
R17060 VSS.n12282 VSS.n12281 0.000511116
R17061 VSS.n12292 VSS.n12291 0.000511116
R17062 VSS.n12310 VSS.n12309 0.000511116
R17063 VSS.n12326 VSS.n12325 0.000511116
R17064 VSS.n12469 VSS.n12468 0.000511116
R17065 VSS.n14510 VSS.n14509 0.000511116
R17066 VSS.n14506 VSS.n14505 0.000511116
R17067 VSS.n6138 VSS.n6137 0.000511116
R17068 VSS.n10624 VSS.n10623 0.000511116
R17069 VSS.n6130 VSS.n6129 0.000511116
R17070 VSS.n6114 VSS.n6113 0.000511116
R17071 VSS.n5948 VSS.n5947 0.000511116
R17072 VSS.n5932 VSS.n5931 0.000511116
R17073 VSS.n5767 VSS.n5766 0.000511116
R17074 VSS.n5751 VSS.n5750 0.000511116
R17075 VSS.n5587 VSS.n5586 0.000511116
R17076 VSS.n5571 VSS.n5570 0.000511116
R17077 VSS.n5407 VSS.n5406 0.000511116
R17078 VSS.n5391 VSS.n5390 0.000511116
R17079 VSS.n5227 VSS.n5226 0.000511116
R17080 VSS.n5211 VSS.n5210 0.000511116
R17081 VSS.n10114 VSS.n10113 0.000511116
R17082 VSS.n10159 VSS.n10158 0.000511116
R17083 VSS.n11157 VSS.n11156 0.000511116
R17084 VSS.n11173 VSS.n11172 0.000511116
R17085 VSS.n3179 VSS.n3178 0.000511116
R17086 VSS.n12562 VSS.n12561 0.000511116
R17087 VSS.n3324 VSS.n3323 0.000511116
R17088 VSS.n3407 VSS.n3406 0.000511116
R17089 VSS.n3577 VSS.n3576 0.000511116
R17090 VSS.n11892 VSS.n11891 0.000511116
R17091 VSS.n12006 VSS.n12005 0.000511116
R17092 VSS.n12023 VSS.n12022 0.000511116
R17093 VSS.n12173 VSS.n12172 0.000511116
R17094 VSS.n12191 VSS.n12190 0.000511116
R17095 VSS.n12288 VSS.n12287 0.000511116
R17096 VSS.n12316 VSS.n12315 0.000511116
R17097 VSS.n11550 VSS.n11549 0.000511116
R17098 VSS.n3608 VSS.n3607 0.000511116
R17099 VSS.n11478 VSS.n3630 0.000509989
R17100 VSS.n14481 VSS.n14480 0.000509339
R17101 VSS.n14480 VSS.n14473 0.000509339
R17102 VSS.n18 VSS.n17 0.000509339
R17103 VSS.n3208 VSS.n3196 0.000509339
R17104 VSS.n3208 VSS.n3197 0.000509339
R17105 VSS.n14503 VSS.n14500 0.000509339
R17106 VSS.n14473 VSS.n14472 0.000509339
R17107 VSS.n14475 VSS.n14474 0.000509339
R17108 VSS.n14507 VSS.n14506 0.000509339
R17109 VSS.n8494 VSS.n8178 0.000507923
R17110 VSS.n8826 VSS.n8178 0.000507923
R17111 VSS.n8372 VSS.n8370 0.000507923
R17112 VSS.n8370 VSS.n8183 0.000507923
R17113 VSS.n8393 VSS.n8210 0.000507923
R17114 VSS.n8788 VSS.n8210 0.000507923
R17115 VSS.n8589 VSS.n8588 0.000507923
R17116 VSS.n8615 VSS.n8589 0.000507923
R17117 VSS.n6760 VSS.n6759 0.000507923
R17118 VSS.n6761 VSS.n6760 0.000507923
R17119 VSS.n8026 VSS.n8020 0.000507923
R17120 VSS.n8034 VSS.n8020 0.000507923
R17121 VSS.n8113 VSS.n8112 0.000507923
R17122 VSS.n8114 VSS.n8113 0.000507923
R17123 VSS.n8892 VSS.n8891 0.000507923
R17124 VSS.n8893 VSS.n8892 0.000507923
R17125 VSS.n8268 VSS.n8266 0.000507923
R17126 VSS.n8266 VSS.n7555 0.000507923
R17127 VSS.n9584 VSS.n9583 0.000507923
R17128 VSS.n9583 VSS.n9577 0.000507923
R17129 VSS.n9389 VSS.n9388 0.000507923
R17130 VSS.n9415 VSS.n9389 0.000507923
R17131 VSS.n9784 VSS.n9783 0.000507923
R17132 VSS.n9785 VSS.n9784 0.000507923
R17133 VSS.n7446 VSS.n7445 0.000507923
R17134 VSS.n7472 VSS.n7446 0.000507923
R17135 VSS.n10831 VSS.n10830 0.000507923
R17136 VSS.n10832 VSS.n10831 0.000507923
R17137 VSS.n9083 VSS.n9082 0.000507923
R17138 VSS.n9109 VSS.n9083 0.000507923
R17139 VSS.n9273 VSS.n9004 0.000507923
R17140 VSS.n9516 VSS.n9004 0.000507923
R17141 VSS.n9496 VSS.n9495 0.000507923
R17142 VSS.n9495 VSS.n9016 0.000507923
R17143 VSS.n9470 VSS.n7168 0.000507923
R17144 VSS.n9838 VSS.n7168 0.000507923
R17145 VSS.n9196 VSS.n9195 0.000507923
R17146 VSS.n9195 VSS.n9165 0.000507923
R17147 VSS.n7899 VSS.n7898 0.000507923
R17148 VSS.n7899 VSS.n7814 0.000507923
R17149 VSS.n7626 VSS.n7625 0.000507923
R17150 VSS.n8985 VSS.n7626 0.000507923
R17151 VSS.n7661 VSS.n7660 0.000507923
R17152 VSS.n7775 VSS.n7661 0.000507923
R17153 VSS.n6796 VSS.n6638 0.000507923
R17154 VSS.n6854 VSS.n6638 0.000507923
R17155 VSS.n6864 VSS.n6590 0.000507923
R17156 VSS.n6921 VSS.n6590 0.000507923
R17157 VSS.n6934 VSS.n6933 0.000507923
R17158 VSS.n6934 VSS.n6516 0.000507923
R17159 VSS.n7017 VSS.n6492 0.000507923
R17160 VSS.n7053 VSS.n6492 0.000507923
R17161 VSS.n6016 VSS.n6015 0.000507923
R17162 VSS.n6042 VSS.n6016 0.000507923
R17163 VSS.n5818 VSS.n5817 0.000507923
R17164 VSS.n5844 VSS.n5818 0.000507923
R17165 VSS.n5637 VSS.n5636 0.000507923
R17166 VSS.n5663 VSS.n5637 0.000507923
R17167 VSS.n5457 VSS.n5456 0.000507923
R17168 VSS.n5483 VSS.n5457 0.000507923
R17169 VSS.n5277 VSS.n5276 0.000507923
R17170 VSS.n5303 VSS.n5277 0.000507923
R17171 VSS.n4180 VSS.n4179 0.000507923
R17172 VSS.n4405 VSS.n4180 0.000507923
R17173 VSS.n1021 VSS.n1020 0.000507923
R17174 VSS.n1047 VSS.n1021 0.000507923
R17175 VSS.n10675 VSS.n10674 0.000507923
R17176 VSS.n10704 VSS.n10675 0.000507923
R17177 VSS.n594 VSS.n588 0.000507923
R17178 VSS.n602 VSS.n588 0.000507923
R17179 VSS.n1150 VSS.n1149 0.000507923
R17180 VSS.n1151 VSS.n1150 0.000507923
R17181 VSS.n12452 VSS.n12451 0.000507923
R17182 VSS.n12453 VSS.n12452 0.000507923
R17183 VSS.n2434 VSS.n2433 0.000507923
R17184 VSS.n2434 VSS.n2356 0.000507923
R17185 VSS.n2341 VSS.n2340 0.000507923
R17186 VSS.n2342 VSS.n2341 0.000507923
R17187 VSS.n940 VSS.n891 0.000507923
R17188 VSS.n1165 VSS.n891 0.000507923
R17189 VSS.n1378 VSS.n1377 0.000507923
R17190 VSS.n1377 VSS.n879 0.000507923
R17191 VSS.n14301 VSS.n14300 0.000507923
R17192 VSS.n14332 VSS.n14301 0.000507923
R17193 VSS.n1543 VSS.n1542 0.000507923
R17194 VSS.n1569 VSS.n1543 0.000507923
R17195 VSS.n13852 VSS.n13851 0.000507923
R17196 VSS.n13853 VSS.n13852 0.000507923
R17197 VSS.n13783 VSS.n13782 0.000507923
R17198 VSS.n13809 VSS.n13783 0.000507923
R17199 VSS.n13387 VSS.n13386 0.000507923
R17200 VSS.n13388 VSS.n13387 0.000507923
R17201 VSS.n736 VSS.n735 0.000507923
R17202 VSS.n762 VSS.n736 0.000507923
R17203 VSS.n1443 VSS.n638 0.000507923
R17204 VSS.n14115 VSS.n638 0.000507923
R17205 VSS.n14095 VSS.n14094 0.000507923
R17206 VSS.n14094 VSS.n650 0.000507923
R17207 VSS.n1656 VSS.n1655 0.000507923
R17208 VSS.n14079 VSS.n1656 0.000507923
R17209 VSS.n1179 VSS.n1177 0.000507923
R17210 VSS.n1177 VSS.n818 0.000507923
R17211 VSS.n2037 VSS.n1993 0.000507923
R17212 VSS.n2245 VSS.n1993 0.000507923
R17213 VSS.n2086 VSS.n2068 0.000507923
R17214 VSS.n2180 VSS.n2068 0.000507923
R17215 VSS.n2134 VSS.n1862 0.000507923
R17216 VSS.n13188 VSS.n1862 0.000507923
R17217 VSS.n2644 VSS.n2572 0.000507923
R17218 VSS.n12985 VSS.n2572 0.000507923
R17219 VSS.n2683 VSS.n2682 0.000507923
R17220 VSS.n12949 VSS.n2683 0.000507923
R17221 VSS.n2825 VSS.n2753 0.000507923
R17222 VSS.n12908 VSS.n2753 0.000507923
R17223 VSS.n2863 VSS.n2862 0.000507923
R17224 VSS.n12872 VSS.n2863 0.000507923
R17225 VSS.n11657 VSS.n11656 0.000507923
R17226 VSS.n11676 VSS.n11657 0.000507923
R17227 VSS.n11726 VSS.n11725 0.000507923
R17228 VSS.n11745 VSS.n11726 0.000507923
R17229 VSS.n12072 VSS.n12071 0.000507923
R17230 VSS.n12098 VSS.n12072 0.000507923
R17231 VSS.n11858 VSS.n11857 0.000507923
R17232 VSS.n11877 VSS.n11858 0.000507923
R17233 VSS.n3476 VSS.n3475 0.000507923
R17234 VSS.n3502 VSS.n3476 0.000507923
R17235 VSS.n3266 VSS.n3265 0.000507923
R17236 VSS.n3267 VSS.n3266 0.000507923
R17237 VSS.n3630 VSS.n3629 0.000507583
R17238 VSS.n8569 VSS.n8568 0.00050746
R17239 VSS.n8780 VSS.n8779 0.00050746
R17240 VSS.n8788 VSS.n8784 0.00050746
R17241 VSS.n6743 VSS.n6742 0.00050746
R17242 VSS.n8150 VSS.n8034 0.00050746
R17243 VSS.n8117 VSS.n8038 0.00050746
R17244 VSS.n8875 VSS.n8874 0.00050746
R17245 VSS.n8826 VSS.n8822 0.00050746
R17246 VSS.n8818 VSS.n8188 0.00050746
R17247 VSS.n9556 VSS.n7569 0.00050746
R17248 VSS.n9369 VSS.n9368 0.00050746
R17249 VSS.n9512 VSS.n9017 0.00050746
R17250 VSS.n9834 VSS.n7181 0.00050746
R17251 VSS.n7370 VSS.n7263 0.00050746
R17252 VSS.n9242 VSS.n9213 0.00050746
R17253 VSS.n8949 VSS.n7852 0.00050746
R17254 VSS.n7639 VSS.n7638 0.00050746
R17255 VSS.n7674 VSS.n7673 0.00050746
R17256 VSS.n7140 VSS.n7090 0.00050746
R17257 VSS.n8924 VSS.n7942 0.00050746
R17258 VSS.n6857 VSS.n6630 0.00050746
R17259 VSS.n6924 VSS.n6582 0.00050746
R17260 VSS.n6997 VSS.n6541 0.00050746
R17261 VSS.n7056 VSS.n6484 0.00050746
R17262 VSS.n6424 VSS.n6317 0.00050746
R17263 VSS.n6789 VSS.n6677 0.00050746
R17264 VSS.n5996 VSS.n5995 0.00050746
R17265 VSS.n5437 VSS.n5436 0.00050746
R17266 VSS.n11028 VSS.n11027 0.00050746
R17267 VSS.n10946 VSS.n10917 0.00050746
R17268 VSS.n10877 VSS.n10876 0.00050746
R17269 VSS.n4269 VSS.n4267 0.00050746
R17270 VSS.n4381 VSS.n4378 0.00050746
R17271 VSS.n4452 VSS.n4133 0.00050746
R17272 VSS.n657 VSS.n656 0.00050746
R17273 VSS.n1001 VSS.n1000 0.00050746
R17274 VSS.n10704 VSS.n10695 0.00050746
R17275 VSS.n14200 VSS.n602 0.00050746
R17276 VSS.n1133 VSS.n1132 0.00050746
R17277 VSS.n13048 VSS.n2483 0.00050746
R17278 VSS.n2453 VSS.n2356 0.00050746
R17279 VSS.n13095 VSS.n13093 0.00050746
R17280 VSS.n2345 VSS.n1931 0.00050746
R17281 VSS.n2400 VSS.n2399 0.00050746
R17282 VSS.n1168 VSS.n883 0.00050746
R17283 VSS.n14305 VSS.n14304 0.00050746
R17284 VSS.n716 VSS.n715 0.00050746
R17285 VSS.n14111 VSS.n651 0.00050746
R17286 VSS.n1669 VSS.n1668 0.00050746
R17287 VSS.n13646 VSS.n13224 0.00050746
R17288 VSS.n1412 VSS.n842 0.00050746
R17289 VSS.n2241 VSS.n2006 0.00050746
R17290 VSS.n2176 VSS.n2081 0.00050746
R17291 VSS.n13191 VSS.n1854 0.00050746
R17292 VSS.n13929 VSS.n13927 0.00050746
R17293 VSS.n1976 VSS.n1975 0.00050746
R17294 VSS.n12981 VSS.n2585 0.00050746
R17295 VSS.n2696 VSS.n2695 0.00050746
R17296 VSS.n12904 VSS.n2766 0.00050746
R17297 VSS.n2876 VSS.n2875 0.00050746
R17298 VSS.n12724 VSS.n12722 0.00050746
R17299 VSS.n2528 VSS.n2527 0.00050746
R17300 VSS.n11574 VSS.n11572 0.00050746
R17301 VSS.n3221 VSS.n3220 0.00050746
R17302 VSS.n12782 VSS.n12781 0.00050746
R17303 VSS.n1766 VSS.n1764 0.00050746
R17304 VSS.n13585 VSS.n13583 0.00050746
R17305 VSS.n13469 VSS.n13468 0.000507003
R17306 VSS.n13463 VSS.n13462 0.000507003
R17307 VSS.n13456 VSS.n13455 0.000507003
R17308 VSS.n13473 VSS.n13456 0.000507003
R17309 VSS.n13476 VSS.n13475 0.000507003
R17310 VSS.n13599 VSS.n13505 0.000507003
R17311 VSS.n13596 VSS.n13593 0.000507003
R17312 VSS.n13589 VSS.n13502 0.000507003
R17313 VSS.n13603 VSS.n13502 0.000507003
R17314 VSS.n13507 VSS.n13506 0.000507003
R17315 VSS.n14012 VSS.n1740 0.000507003
R17316 VSS.n14009 VSS.n14006 0.000507003
R17317 VSS.n1763 VSS.n1737 0.000507003
R17318 VSS.n14016 VSS.n1737 0.000507003
R17319 VSS.n1742 VSS.n1741 0.000507003
R17320 VSS.n2934 VSS.n2933 0.000507003
R17321 VSS.n12792 VSS.n12787 0.000507003
R17322 VSS.n12785 VSS.n2930 0.000507003
R17323 VSS.n12796 VSS.n12785 0.000507003
R17324 VSS.n12800 VSS.n2932 0.000507003
R17325 VSS.n4079 VSS.n4078 0.000507003
R17326 VSS.n4073 VSS.n4072 0.000507003
R17327 VSS.n4066 VSS.n4065 0.000507003
R17328 VSS.n4083 VSS.n4066 0.000507003
R17329 VSS.n4061 VSS.n4060 0.000507003
R17330 VSS.n3897 VSS.n3896 0.000507003
R17331 VSS.n10887 VSS.n10882 0.000507003
R17332 VSS.n10880 VSS.n3893 0.000507003
R17333 VSS.n10891 VSS.n10880 0.000507003
R17334 VSS.n10895 VSS.n3895 0.000507003
R17335 VSS.n10936 VSS.n10924 0.000507003
R17336 VSS.n10933 VSS.n10932 0.000507003
R17337 VSS.n10943 VSS.n10942 0.000507003
R17338 VSS.n10943 VSS.n3859 0.000507003
R17339 VSS.n10940 VSS.n10923 0.000507003
R17340 VSS.n3829 VSS.n3828 0.000507003
R17341 VSS.n11038 VSS.n11033 0.000507003
R17342 VSS.n11031 VSS.n3825 0.000507003
R17343 VSS.n11042 VSS.n11031 0.000507003
R17344 VSS.n11046 VSS.n3827 0.000507003
R17345 VSS.n9677 VSS.n9676 0.000507003
R17346 VSS.n9671 VSS.n9670 0.000507003
R17347 VSS.n9693 VSS.n9692 0.000507003
R17348 VSS.n9665 VSS.n9664 0.000507003
R17349 VSS.n9136 VSS.n9135 0.000507003
R17350 VSS.n9137 VSS.n9136 0.000507003
R17351 VSS.n9130 VSS.n9129 0.000507003
R17352 VSS.n9124 VSS.n9123 0.000507003
R17353 VSS.n9048 VSS.n9047 0.000507003
R17354 VSS.n9137 VSS.n9048 0.000507003
R17355 VSS.n9140 VSS.n9139 0.000507003
R17356 VSS.n9043 VSS.n9042 0.000507003
R17357 VSS.n9037 VSS.n9036 0.000507003
R17358 VSS.n9027 VSS.n9026 0.000507003
R17359 VSS.n9655 VSS.n9654 0.000507003
R17360 VSS.n9649 VSS.n9648 0.000507003
R17361 VSS.n9660 VSS.n9659 0.000507003
R17362 VSS.n9686 VSS.n9685 0.000507003
R17363 VSS.n8356 VSS.n8355 0.000507003
R17364 VSS.n8362 VSS.n8361 0.000507003
R17365 VSS.n8560 VSS.n8559 0.000507003
R17366 VSS.n8481 VSS.n8480 0.000507003
R17367 VSS.n8482 VSS.n8481 0.000507003
R17368 VSS.n8475 VSS.n8474 0.000507003
R17369 VSS.n8465 VSS.n8464 0.000507003
R17370 VSS.n8485 VSS.n8484 0.000507003
R17371 VSS.n8185 VSS.n8184 0.000507003
R17372 VSS.n8507 VSS.n8506 0.000507003
R17373 VSS.n8501 VSS.n8500 0.000507003
R17374 VSS.n8497 VSS.n8496 0.000507003
R17375 VSS.n8376 VSS.n8369 0.000507003
R17376 VSS.n8380 VSS.n8379 0.000507003
R17377 VSS.n8387 VSS.n8386 0.000507003
R17378 VSS.n8217 VSS.n8216 0.000507003
R17379 VSS.n8406 VSS.n8405 0.000507003
R17380 VSS.n8400 VSS.n8399 0.000507003
R17381 VSS.n8396 VSS.n8395 0.000507003
R17382 VSS.n8689 VSS.n8688 0.000507003
R17383 VSS.n8683 VSS.n8682 0.000507003
R17384 VSS.n8705 VSS.n8704 0.000507003
R17385 VSS.n8677 VSS.n8676 0.000507003
R17386 VSS.n9633 VSS.n9632 0.000507003
R17387 VSS.n9634 VSS.n9633 0.000507003
R17388 VSS.n9627 VSS.n9626 0.000507003
R17389 VSS.n9637 VSS.n9636 0.000507003
R17390 VSS.n9620 VSS.n9619 0.000507003
R17391 VSS.n9634 VSS.n9620 0.000507003
R17392 VSS.n9615 VSS.n9614 0.000507003
R17393 VSS.n7544 VSS.n7543 0.000507003
R17394 VSS.n7538 VSS.n7537 0.000507003
R17395 VSS.n7528 VSS.n7527 0.000507003
R17396 VSS.n8667 VSS.n8666 0.000507003
R17397 VSS.n8661 VSS.n8660 0.000507003
R17398 VSS.n8672 VSS.n8671 0.000507003
R17399 VSS.n8698 VSS.n8697 0.000507003
R17400 VSS.n8310 VSS.n8309 0.000507003
R17401 VSS.n8316 VSS.n8315 0.000507003
R17402 VSS.n8737 VSS.n8736 0.000507003
R17403 VSS.n8740 VSS.n8739 0.000507003
R17404 VSS.n8614 VSS.n8613 0.000507003
R17405 VSS.n8615 VSS.n8614 0.000507003
R17406 VSS.n8609 VSS.n8608 0.000507003
R17407 VSS.n8602 VSS.n8601 0.000507003
R17408 VSS.n8596 VSS.n8595 0.000507003
R17409 VSS.n8584 VSS.n8583 0.000507003
R17410 VSS.n8578 VSS.n8577 0.000507003
R17411 VSS.n8618 VSS.n8617 0.000507003
R17412 VSS.n8572 VSS.n8571 0.000507003
R17413 VSS.n8298 VSS.n8297 0.000507003
R17414 VSS.n8292 VSS.n8291 0.000507003
R17415 VSS.n8743 VSS.n8742 0.000507003
R17416 VSS.n8752 VSS.n8751 0.000507003
R17417 VSS.n8253 VSS.n8252 0.000507003
R17418 VSS.n8253 VSS.n8215 0.000507003
R17419 VSS.n8259 VSS.n8258 0.000507003
R17420 VSS.n8773 VSS.n8244 0.000507003
R17421 VSS.n8242 VSS.n8218 0.000507003
R17422 VSS.n8242 VSS.n8215 0.000507003
R17423 VSS.n8239 VSS.n8238 0.000507003
R17424 VSS.n8235 VSS.n8234 0.000507003
R17425 VSS.n8231 VSS.n8230 0.000507003
R17426 VSS.n8777 VSS.n8219 0.000507003
R17427 VSS.n8198 VSS.n8197 0.000507003
R17428 VSS.n8205 VSS.n8200 0.000507003
R17429 VSS.n8785 VSS.n8194 0.000507003
R17430 VSS.n8792 VSS.n8196 0.000507003
R17431 VSS.n6202 VSS.n6201 0.000507003
R17432 VSS.n6203 VSS.n6202 0.000507003
R17433 VSS.n6196 VSS.n6195 0.000507003
R17434 VSS.n6186 VSS.n6185 0.000507003
R17435 VSS.n6206 VSS.n6205 0.000507003
R17436 VSS.n9977 VSS.n6213 0.000507003
R17437 VSS.n9981 VSS.n9980 0.000507003
R17438 VSS.n6222 VSS.n6221 0.000507003
R17439 VSS.n6226 VSS.n6220 0.000507003
R17440 VSS.n6757 VSS.n6756 0.000507003
R17441 VSS.n6753 VSS.n6752 0.000507003
R17442 VSS.n6749 VSS.n6748 0.000507003
R17443 VSS.n6711 VSS.n6692 0.000507003
R17444 VSS.n6761 VSS.n6711 0.000507003
R17445 VSS.n6765 VSS.n6764 0.000507003
R17446 VSS.n6701 VSS.n6696 0.000507003
R17447 VSS.n6706 VSS.n6700 0.000507003
R17448 VSS.n6745 VSS.n6744 0.000507003
R17449 VSS.n9965 VSS.n9964 0.000507003
R17450 VSS.n9961 VSS.n9960 0.000507003
R17451 VSS.n9973 VSS.n9972 0.000507003
R17452 VSS.n9970 VSS.n9969 0.000507003
R17453 VSS.n8151 VSS.n8016 0.000507003
R17454 VSS.n8155 VSS.n8154 0.000507003
R17455 VSS.n8032 VSS.n8031 0.000507003
R17456 VSS.n8029 VSS.n8028 0.000507003
R17457 VSS.n8110 VSS.n8109 0.000507003
R17458 VSS.n8106 VSS.n8105 0.000507003
R17459 VSS.n8102 VSS.n8101 0.000507003
R17460 VSS.n8115 VSS.n8036 0.000507003
R17461 VSS.n8115 VSS.n8114 0.000507003
R17462 VSS.n8090 VSS.n8089 0.000507003
R17463 VSS.n8085 VSS.n8084 0.000507003
R17464 VSS.n8081 VSS.n8080 0.000507003
R17465 VSS.n8041 VSS.n8037 0.000507003
R17466 VSS.n8141 VSS.n8129 0.000507003
R17467 VSS.n8138 VSS.n8137 0.000507003
R17468 VSS.n8147 VSS.n8120 0.000507003
R17469 VSS.n8145 VSS.n8128 0.000507003
R17470 VSS.n8068 VSS.n8001 0.000507003
R17471 VSS.n8072 VSS.n8071 0.000507003
R17472 VSS.n8064 VSS.n8063 0.000507003
R17473 VSS.n8061 VSS.n8060 0.000507003
R17474 VSS.n8889 VSS.n8888 0.000507003
R17475 VSS.n8885 VSS.n8884 0.000507003
R17476 VSS.n8881 VSS.n8880 0.000507003
R17477 VSS.n7968 VSS.n7948 0.000507003
R17478 VSS.n8893 VSS.n7968 0.000507003
R17479 VSS.n8897 VSS.n8896 0.000507003
R17480 VSS.n7958 VSS.n7952 0.000507003
R17481 VSS.n7963 VSS.n7957 0.000507003
R17482 VSS.n8877 VSS.n8876 0.000507003
R17483 VSS.n8862 VSS.n8861 0.000507003
R17484 VSS.n8857 VSS.n8856 0.000507003
R17485 VSS.n8870 VSS.n8869 0.000507003
R17486 VSS.n8865 VSS.n8864 0.000507003
R17487 VSS.n8816 VSS.n8186 0.000507003
R17488 VSS.n8816 VSS.n8183 0.000507003
R17489 VSS.n8813 VSS.n8812 0.000507003
R17490 VSS.n8808 VSS.n8807 0.000507003
R17491 VSS.n8804 VSS.n8803 0.000507003
R17492 VSS.n8383 VSS.n8187 0.000507003
R17493 VSS.n8166 VSS.n8165 0.000507003
R17494 VSS.n8173 VSS.n8168 0.000507003
R17495 VSS.n8823 VSS.n8162 0.000507003
R17496 VSS.n8830 VSS.n8164 0.000507003
R17497 VSS.n9554 VSS.n7567 0.000507003
R17498 VSS.n9554 VSS.n7555 0.000507003
R17499 VSS.n9551 VSS.n9550 0.000507003
R17500 VSS.n7586 VSS.n7576 0.000507003
R17501 VSS.n7582 VSS.n7577 0.000507003
R17502 VSS.n8272 VSS.n8265 0.000507003
R17503 VSS.n8276 VSS.n8275 0.000507003
R17504 VSS.n8283 VSS.n8282 0.000507003
R17505 VSS.n8279 VSS.n7568 0.000507003
R17506 VSS.n9562 VSS.n9561 0.000507003
R17507 VSS.n9565 VSS.n9564 0.000507003
R17508 VSS.n9570 VSS.n9569 0.000507003
R17509 VSS.n9573 VSS.n7563 0.000507003
R17510 VSS.n9586 VSS.n9579 0.000507003
R17511 VSS.n9590 VSS.n9578 0.000507003
R17512 VSS.n9594 VSS.n9593 0.000507003
R17513 VSS.n7557 VSS.n7551 0.000507003
R17514 VSS.n8346 VSS.n8345 0.000507003
R17515 VSS.n8532 VSS.n8531 0.000507003
R17516 VSS.n8538 VSS.n8537 0.000507003
R17517 VSS.n8544 VSS.n8543 0.000507003
R17518 VSS.n8555 VSS.n8554 0.000507003
R17519 VSS.n8458 VSS.n8457 0.000507003
R17520 VSS.n8482 VSS.n8458 0.000507003
R17521 VSS.n8452 VSS.n8451 0.000507003
R17522 VSS.n8442 VSS.n8441 0.000507003
R17523 VSS.n8437 VSS.n8436 0.000507003
R17524 VSS.n9414 VSS.n9413 0.000507003
R17525 VSS.n9415 VSS.n9414 0.000507003
R17526 VSS.n9409 VSS.n9408 0.000507003
R17527 VSS.n9402 VSS.n9401 0.000507003
R17528 VSS.n9396 VSS.n9395 0.000507003
R17529 VSS.n9384 VSS.n9383 0.000507003
R17530 VSS.n9378 VSS.n9377 0.000507003
R17531 VSS.n9418 VSS.n9417 0.000507003
R17532 VSS.n9372 VSS.n9371 0.000507003
R17533 VSS.n7390 VSS.n7389 0.000507003
R17534 VSS.n9790 VSS.n9789 0.000507003
R17535 VSS.n7399 VSS.n7398 0.000507003
R17536 VSS.n7405 VSS.n7404 0.000507003
R17537 VSS.n7387 VSS.n7386 0.000507003
R17538 VSS.n7415 VSS.n7414 0.000507003
R17539 VSS.n9779 VSS.n9778 0.000507003
R17540 VSS.n7393 VSS.n7392 0.000507003
R17541 VSS.n7471 VSS.n7470 0.000507003
R17542 VSS.n7472 VSS.n7471 0.000507003
R17543 VSS.n7466 VSS.n7465 0.000507003
R17544 VSS.n7459 VSS.n7458 0.000507003
R17545 VSS.n7453 VSS.n7452 0.000507003
R17546 VSS.n7441 VSS.n7440 0.000507003
R17547 VSS.n7435 VSS.n7434 0.000507003
R17548 VSS.n7475 VSS.n7474 0.000507003
R17549 VSS.n7429 VSS.n7428 0.000507003
R17550 VSS.n10837 VSS.n10836 0.000507003
R17551 VSS.n3935 VSS.n3934 0.000507003
R17552 VSS.n3941 VSS.n3940 0.000507003
R17553 VSS.n3931 VSS.n3930 0.000507003
R17554 VSS.n3923 VSS.n3922 0.000507003
R17555 VSS.n3951 VSS.n3950 0.000507003
R17556 VSS.n10826 VSS.n10825 0.000507003
R17557 VSS.n3926 VSS.n3925 0.000507003
R17558 VSS.n9344 VSS.n9343 0.000507003
R17559 VSS.n9350 VSS.n9349 0.000507003
R17560 VSS.n9434 VSS.n9433 0.000507003
R17561 VSS.n9437 VSS.n9436 0.000507003
R17562 VSS.n9108 VSS.n9107 0.000507003
R17563 VSS.n9109 VSS.n9108 0.000507003
R17564 VSS.n9103 VSS.n9102 0.000507003
R17565 VSS.n9096 VSS.n9095 0.000507003
R17566 VSS.n9090 VSS.n9089 0.000507003
R17567 VSS.n9078 VSS.n9077 0.000507003
R17568 VSS.n9072 VSS.n9071 0.000507003
R17569 VSS.n9112 VSS.n9111 0.000507003
R17570 VSS.n9066 VSS.n9065 0.000507003
R17571 VSS.n9332 VSS.n9331 0.000507003
R17572 VSS.n9326 VSS.n9325 0.000507003
R17573 VSS.n9440 VSS.n9439 0.000507003
R17574 VSS.n9449 VSS.n9448 0.000507003
R17575 VSS.n9515 VSS.n8994 0.000507003
R17576 VSS.n9516 VSS.n9515 0.000507003
R17577 VSS.n9520 VSS.n8996 0.000507003
R17578 VSS.n8998 VSS.n8997 0.000507003
R17579 VSS.n9011 VSS.n9006 0.000507003
R17580 VSS.n9278 VSS.n9277 0.000507003
R17581 VSS.n9282 VSS.n9281 0.000507003
R17582 VSS.n9287 VSS.n9286 0.000507003
R17583 VSS.n9290 VSS.n9289 0.000507003
R17584 VSS.n9311 VSS.n9310 0.000507003
R17585 VSS.n9307 VSS.n9306 0.000507003
R17586 VSS.n9303 VSS.n9302 0.000507003
R17587 VSS.n9314 VSS.n9291 0.000507003
R17588 VSS.n9499 VSS.n9491 0.000507003
R17589 VSS.n9503 VSS.n9490 0.000507003
R17590 VSS.n9507 VSS.n9506 0.000507003
R17591 VSS.n9509 VSS.n9319 0.000507003
R17592 VSS.n7221 VSS.n7184 0.000507003
R17593 VSS.n7225 VSS.n7224 0.000507003
R17594 VSS.n7238 VSS.n7237 0.000507003
R17595 VSS.n7234 VSS.n7228 0.000507003
R17596 VSS.n7230 VSS.n7229 0.000507003
R17597 VSS.n7229 VSS.n7180 0.000507003
R17598 VSS.n9837 VSS.n7158 0.000507003
R17599 VSS.n9838 VSS.n9837 0.000507003
R17600 VSS.n9842 VSS.n7160 0.000507003
R17601 VSS.n7162 VSS.n7161 0.000507003
R17602 VSS.n7175 VSS.n7170 0.000507003
R17603 VSS.n9474 VSS.n9473 0.000507003
R17604 VSS.n9484 VSS.n9477 0.000507003
R17605 VSS.n9481 VSS.n9478 0.000507003
R17606 VSS.n7183 VSS.n7182 0.000507003
R17607 VSS.n9823 VSS.n9822 0.000507003
R17608 VSS.n9819 VSS.n9818 0.000507003
R17609 VSS.n9829 VSS.n9828 0.000507003
R17610 VSS.n9831 VSS.n7188 0.000507003
R17611 VSS.n7260 VSS.n7259 0.000507003
R17612 VSS.n7256 VSS.n7255 0.000507003
R17613 VSS.n7253 VSS.n7214 0.000507003
R17614 VSS.n7250 VSS.n7249 0.000507003
R17615 VSS.n7366 VSS.n7365 0.000507003
R17616 VSS.n7367 VSS.n7366 0.000507003
R17617 VSS.n7361 VSS.n7360 0.000507003
R17618 VSS.n7357 VSS.n7356 0.000507003
R17619 VSS.n7368 VSS.n7261 0.000507003
R17620 VSS.n7368 VSS.n7367 0.000507003
R17621 VSS.n7316 VSS.n7315 0.000507003
R17622 VSS.n7327 VSS.n7326 0.000507003
R17623 VSS.n7323 VSS.n7319 0.000507003
R17624 VSS.n7266 VSS.n7262 0.000507003
R17625 VSS.n7203 VSS.n7200 0.000507003
R17626 VSS.n7206 VSS.n7205 0.000507003
R17627 VSS.n7378 VSS.n7192 0.000507003
R17628 VSS.n7375 VSS.n7190 0.000507003
R17629 VSS.n9177 VSS.n9176 0.000507003
R17630 VSS.n9180 VSS.n9179 0.000507003
R17631 VSS.n9268 VSS.n9267 0.000507003
R17632 VSS.n9182 VSS.n9160 0.000507003
R17633 VSS.n9240 VSS.n9187 0.000507003
R17634 VSS.n9240 VSS.n9165 0.000507003
R17635 VSS.n9237 VSS.n9236 0.000507003
R17636 VSS.n9230 VSS.n9220 0.000507003
R17637 VSS.n9226 VSS.n9221 0.000507003
R17638 VSS.n9199 VSS.n9191 0.000507003
R17639 VSS.n9203 VSS.n9190 0.000507003
R17640 VSS.n9208 VSS.n9189 0.000507003
R17641 VSS.n9212 VSS.n9188 0.000507003
R17642 VSS.n9257 VSS.n9256 0.000507003
R17643 VSS.n9252 VSS.n9251 0.000507003
R17644 VSS.n9246 VSS.n9186 0.000507003
R17645 VSS.n9261 VSS.n9185 0.000507003
R17646 VSS.n7849 VSS.n7848 0.000507003
R17647 VSS.n7846 VSS.n7845 0.000507003
R17648 VSS.n8961 VSS.n8960 0.000507003
R17649 VSS.n7821 VSS.n7820 0.000507003
R17650 VSS.n7822 VSS.n7818 0.000507003
R17651 VSS.n8958 VSS.n7818 0.000507003
R17652 VSS.n8947 VSS.n7850 0.000507003
R17653 VSS.n8947 VSS.n7814 0.000507003
R17654 VSS.n8944 VSS.n8943 0.000507003
R17655 VSS.n7869 VSS.n7859 0.000507003
R17656 VSS.n7865 VSS.n7860 0.000507003
R17657 VSS.n7903 VSS.n7902 0.000507003
R17658 VSS.n7916 VSS.n7906 0.000507003
R17659 VSS.n7912 VSS.n7907 0.000507003
R17660 VSS.n7909 VSS.n7851 0.000507003
R17661 VSS.n7841 VSS.n7840 0.000507003
R17662 VSS.n7836 VSS.n7835 0.000507003
R17663 VSS.n7844 VSS.n7829 0.000507003
R17664 VSS.n8954 VSS.n7830 0.000507003
R17665 VSS.n7734 VSS.n7640 0.000507003
R17666 VSS.n7738 VSS.n7737 0.000507003
R17667 VSS.n7751 VSS.n7750 0.000507003
R17668 VSS.n7747 VSS.n7741 0.000507003
R17669 VSS.n7743 VSS.n7742 0.000507003
R17670 VSS.n7742 VSS.n7631 0.000507003
R17671 VSS.n8984 VSS.n8983 0.000507003
R17672 VSS.n8985 VSS.n8984 0.000507003
R17673 VSS.n8981 VSS.n8967 0.000507003
R17674 VSS.n8978 VSS.n8968 0.000507003
R17675 VSS.n8975 VSS.n8972 0.000507003
R17676 VSS.n7623 VSS.n7622 0.000507003
R17677 VSS.n8989 VSS.n7613 0.000507003
R17678 VSS.n7615 VSS.n7614 0.000507003
R17679 VSS.n7637 VSS.n7636 0.000507003
R17680 VSS.n7796 VSS.n7795 0.000507003
R17681 VSS.n7792 VSS.n7791 0.000507003
R17682 VSS.n7802 VSS.n7801 0.000507003
R17683 VSS.n7804 VSS.n7644 0.000507003
R17684 VSS.n7698 VSS.n7675 0.000507003
R17685 VSS.n7695 VSS.n7676 0.000507003
R17686 VSS.n7691 VSS.n7677 0.000507003
R17687 VSS.n7687 VSS.n7679 0.000507003
R17688 VSS.n7685 VSS.n7684 0.000507003
R17689 VSS.n7684 VSS.n7666 0.000507003
R17690 VSS.n7774 VSS.n7773 0.000507003
R17691 VSS.n7775 VSS.n7774 0.000507003
R17692 VSS.n7771 VSS.n7757 0.000507003
R17693 VSS.n7768 VSS.n7758 0.000507003
R17694 VSS.n7765 VSS.n7762 0.000507003
R17695 VSS.n7658 VSS.n7657 0.000507003
R17696 VSS.n7779 VSS.n7648 0.000507003
R17697 VSS.n7650 VSS.n7649 0.000507003
R17698 VSS.n7672 VSS.n7671 0.000507003
R17699 VSS.n7717 VSS.n7716 0.000507003
R17700 VSS.n7713 VSS.n7712 0.000507003
R17701 VSS.n7723 VSS.n7722 0.000507003
R17702 VSS.n7725 VSS.n7703 0.000507003
R17703 VSS.n9892 VSS.n7070 0.000507003
R17704 VSS.n9896 VSS.n9895 0.000507003
R17705 VSS.n7079 VSS.n7078 0.000507003
R17706 VSS.n7083 VSS.n7077 0.000507003
R17707 VSS.n7136 VSS.n7135 0.000507003
R17708 VSS.n7137 VSS.n7136 0.000507003
R17709 VSS.n7131 VSS.n7130 0.000507003
R17710 VSS.n7126 VSS.n7125 0.000507003
R17711 VSS.n7138 VSS.n7088 0.000507003
R17712 VSS.n7138 VSS.n7137 0.000507003
R17713 VSS.n7114 VSS.n7113 0.000507003
R17714 VSS.n7110 VSS.n7109 0.000507003
R17715 VSS.n7105 VSS.n7102 0.000507003
R17716 VSS.n7093 VSS.n7089 0.000507003
R17717 VSS.n9876 VSS.n9875 0.000507003
R17718 VSS.n9880 VSS.n9879 0.000507003
R17719 VSS.n9885 VSS.n9884 0.000507003
R17720 VSS.n9888 VSS.n9887 0.000507003
R17721 VSS.n7926 VSS.n7925 0.000507003
R17722 VSS.n7931 VSS.n7930 0.000507003
R17723 VSS.n7935 VSS.n7934 0.000507003
R17724 VSS.n7939 VSS.n7938 0.000507003
R17725 VSS.n8922 VSS.n7940 0.000507003
R17726 VSS.n8922 VSS.n7877 0.000507003
R17727 VSS.n8919 VSS.n8918 0.000507003
R17728 VSS.n8914 VSS.n8913 0.000507003
R17729 VSS.n8910 VSS.n8909 0.000507003
R17730 VSS.n7993 VSS.n7941 0.000507003
R17731 VSS.n7993 VSS.n7877 0.000507003
R17732 VSS.n7997 VSS.n7996 0.000507003
R17733 VSS.n7990 VSS.n7989 0.000507003
R17734 VSS.n7987 VSS.n7982 0.000507003
R17735 VSS.n7876 VSS.n7875 0.000507003
R17736 VSS.n7884 VSS.n7879 0.000507003
R17737 VSS.n8936 VSS.n7874 0.000507003
R17738 VSS.n8929 VSS.n7872 0.000507003
R17739 VSS.n6855 VSS.n6628 0.000507003
R17740 VSS.n6855 VSS.n6854 0.000507003
R17741 VSS.n6852 VSS.n6851 0.000507003
R17742 VSS.n6654 VSS.n6646 0.000507003
R17743 VSS.n6651 VSS.n6647 0.000507003
R17744 VSS.n6800 VSS.n6799 0.000507003
R17745 VSS.n6810 VSS.n6803 0.000507003
R17746 VSS.n6807 VSS.n6804 0.000507003
R17747 VSS.n6633 VSS.n6629 0.000507003
R17748 VSS.n6907 VSS.n6609 0.000507003
R17749 VSS.n6911 VSS.n6910 0.000507003
R17750 VSS.n6624 VSS.n6623 0.000507003
R17751 VSS.n6621 VSS.n6620 0.000507003
R17752 VSS.n6891 VSS.n6890 0.000507003
R17753 VSS.n6895 VSS.n6894 0.000507003
R17754 VSS.n6901 VSS.n6900 0.000507003
R17755 VSS.n6903 VSS.n6860 0.000507003
R17756 VSS.n6922 VSS.n6580 0.000507003
R17757 VSS.n6922 VSS.n6921 0.000507003
R17758 VSS.n6919 VSS.n6918 0.000507003
R17759 VSS.n6606 VSS.n6598 0.000507003
R17760 VSS.n6603 VSS.n6599 0.000507003
R17761 VSS.n6868 VSS.n6867 0.000507003
R17762 VSS.n6878 VSS.n6871 0.000507003
R17763 VSS.n6875 VSS.n6872 0.000507003
R17764 VSS.n6585 VSS.n6581 0.000507003
R17765 VSS.n6980 VSS.n6561 0.000507003
R17766 VSS.n6984 VSS.n6983 0.000507003
R17767 VSS.n6576 VSS.n6575 0.000507003
R17768 VSS.n6573 VSS.n6572 0.000507003
R17769 VSS.n6964 VSS.n6963 0.000507003
R17770 VSS.n6968 VSS.n6967 0.000507003
R17771 VSS.n6974 VSS.n6973 0.000507003
R17772 VSS.n6976 VSS.n6927 0.000507003
R17773 VSS.n6538 VSS.n6537 0.000507003
R17774 VSS.n6535 VSS.n6534 0.000507003
R17775 VSS.n7043 VSS.n7042 0.000507003
R17776 VSS.n6523 VSS.n6522 0.000507003
R17777 VSS.n6524 VSS.n6520 0.000507003
R17778 VSS.n7040 VSS.n6520 0.000507003
R17779 VSS.n6995 VSS.n6539 0.000507003
R17780 VSS.n6995 VSS.n6516 0.000507003
R17781 VSS.n6992 VSS.n6991 0.000507003
R17782 VSS.n6558 VSS.n6548 0.000507003
R17783 VSS.n6554 VSS.n6549 0.000507003
R17784 VSS.n6938 VSS.n6937 0.000507003
R17785 VSS.n6951 VSS.n6941 0.000507003
R17786 VSS.n6947 VSS.n6942 0.000507003
R17787 VSS.n6944 VSS.n6540 0.000507003
R17788 VSS.n7012 VSS.n7011 0.000507003
R17789 VSS.n7006 VSS.n7005 0.000507003
R17790 VSS.n6533 VSS.n6531 0.000507003
R17791 VSS.n7036 VSS.n6532 0.000507003
R17792 VSS.n6481 VSS.n6480 0.000507003
R17793 VSS.n6478 VSS.n6293 0.000507003
R17794 VSS.n6474 VSS.n6294 0.000507003
R17795 VSS.n6471 VSS.n6470 0.000507003
R17796 VSS.n6467 VSS.n6463 0.000507003
R17797 VSS.n6467 VSS.n6289 0.000507003
R17798 VSS.n7054 VSS.n6482 0.000507003
R17799 VSS.n7054 VSS.n7053 0.000507003
R17800 VSS.n7051 VSS.n7050 0.000507003
R17801 VSS.n6508 VSS.n6500 0.000507003
R17802 VSS.n6505 VSS.n6501 0.000507003
R17803 VSS.n7021 VSS.n7020 0.000507003
R17804 VSS.n7031 VSS.n7024 0.000507003
R17805 VSS.n7028 VSS.n7025 0.000507003
R17806 VSS.n6487 VSS.n6483 0.000507003
R17807 VSS.n6286 VSS.n6285 0.000507003
R17808 VSS.n6283 VSS.n6282 0.000507003
R17809 VSS.n7064 VSS.n6273 0.000507003
R17810 VSS.n7061 VSS.n6271 0.000507003
R17811 VSS.n6454 VSS.n6297 0.000507003
R17812 VSS.n6458 VSS.n6457 0.000507003
R17813 VSS.n6306 VSS.n6305 0.000507003
R17814 VSS.n6310 VSS.n6304 0.000507003
R17815 VSS.n6420 VSS.n6419 0.000507003
R17816 VSS.n6421 VSS.n6420 0.000507003
R17817 VSS.n6415 VSS.n6414 0.000507003
R17818 VSS.n6411 VSS.n6410 0.000507003
R17819 VSS.n6422 VSS.n6315 0.000507003
R17820 VSS.n6422 VSS.n6421 0.000507003
R17821 VSS.n6370 VSS.n6369 0.000507003
R17822 VSS.n6381 VSS.n6380 0.000507003
R17823 VSS.n6377 VSS.n6373 0.000507003
R17824 VSS.n6320 VSS.n6316 0.000507003
R17825 VSS.n6438 VSS.n6437 0.000507003
R17826 VSS.n6442 VSS.n6441 0.000507003
R17827 VSS.n6447 VSS.n6446 0.000507003
R17828 VSS.n6450 VSS.n6449 0.000507003
R17829 VSS.n6824 VSS.n6823 0.000507003
R17830 VSS.n6828 VSS.n6827 0.000507003
R17831 VSS.n6833 VSS.n6832 0.000507003
R17832 VSS.n6836 VSS.n6835 0.000507003
R17833 VSS.n6787 VSS.n6675 0.000507003
R17834 VSS.n6787 VSS.n6786 0.000507003
R17835 VSS.n6784 VSS.n6783 0.000507003
R17836 VSS.n6779 VSS.n6778 0.000507003
R17837 VSS.n6775 VSS.n6774 0.000507003
R17838 VSS.n6684 VSS.n6676 0.000507003
R17839 VSS.n6786 VSS.n6684 0.000507003
R17840 VSS.n6735 VSS.n6734 0.000507003
R17841 VSS.n6729 VSS.n6728 0.000507003
R17842 VSS.n6725 VSS.n6722 0.000507003
R17843 VSS.n6672 VSS.n6671 0.000507003
R17844 VSS.n6669 VSS.n6668 0.000507003
R17845 VSS.n6840 VSS.n6657 0.000507003
R17846 VSS.n6844 VSS.n6843 0.000507003
R17847 VSS.n6041 VSS.n6040 0.000507003
R17848 VSS.n6042 VSS.n6041 0.000507003
R17849 VSS.n6036 VSS.n6035 0.000507003
R17850 VSS.n6029 VSS.n6028 0.000507003
R17851 VSS.n6023 VSS.n6022 0.000507003
R17852 VSS.n6011 VSS.n6010 0.000507003
R17853 VSS.n6005 VSS.n6004 0.000507003
R17854 VSS.n6045 VSS.n6044 0.000507003
R17855 VSS.n5999 VSS.n5998 0.000507003
R17856 VSS.n5889 VSS.n5888 0.000507003
R17857 VSS.n5900 VSS.n5899 0.000507003
R17858 VSS.n5879 VSS.n5878 0.000507003
R17859 VSS.n5873 VSS.n5872 0.000507003
R17860 VSS.n5863 VSS.n5862 0.000507003
R17861 VSS.n5859 VSS.n5858 0.000507003
R17862 VSS.n5853 VSS.n5852 0.000507003
R17863 VSS.n5884 VSS.n5883 0.000507003
R17864 VSS.n5843 VSS.n5842 0.000507003
R17865 VSS.n5844 VSS.n5843 0.000507003
R17866 VSS.n5838 VSS.n5837 0.000507003
R17867 VSS.n5831 VSS.n5830 0.000507003
R17868 VSS.n5825 VSS.n5824 0.000507003
R17869 VSS.n5813 VSS.n5812 0.000507003
R17870 VSS.n5807 VSS.n5806 0.000507003
R17871 VSS.n5847 VSS.n5846 0.000507003
R17872 VSS.n5801 VSS.n5800 0.000507003
R17873 VSS.n5708 VSS.n5707 0.000507003
R17874 VSS.n5719 VSS.n5718 0.000507003
R17875 VSS.n5698 VSS.n5697 0.000507003
R17876 VSS.n5692 VSS.n5691 0.000507003
R17877 VSS.n5682 VSS.n5681 0.000507003
R17878 VSS.n5678 VSS.n5677 0.000507003
R17879 VSS.n5672 VSS.n5671 0.000507003
R17880 VSS.n5703 VSS.n5702 0.000507003
R17881 VSS.n5662 VSS.n5661 0.000507003
R17882 VSS.n5663 VSS.n5662 0.000507003
R17883 VSS.n5657 VSS.n5656 0.000507003
R17884 VSS.n5650 VSS.n5649 0.000507003
R17885 VSS.n5644 VSS.n5643 0.000507003
R17886 VSS.n5632 VSS.n5631 0.000507003
R17887 VSS.n5626 VSS.n5625 0.000507003
R17888 VSS.n5666 VSS.n5665 0.000507003
R17889 VSS.n5620 VSS.n5619 0.000507003
R17890 VSS.n5528 VSS.n5527 0.000507003
R17891 VSS.n5539 VSS.n5538 0.000507003
R17892 VSS.n5518 VSS.n5517 0.000507003
R17893 VSS.n5512 VSS.n5511 0.000507003
R17894 VSS.n5502 VSS.n5501 0.000507003
R17895 VSS.n5498 VSS.n5497 0.000507003
R17896 VSS.n5492 VSS.n5491 0.000507003
R17897 VSS.n5523 VSS.n5522 0.000507003
R17898 VSS.n5482 VSS.n5481 0.000507003
R17899 VSS.n5483 VSS.n5482 0.000507003
R17900 VSS.n5477 VSS.n5476 0.000507003
R17901 VSS.n5470 VSS.n5469 0.000507003
R17902 VSS.n5464 VSS.n5463 0.000507003
R17903 VSS.n5452 VSS.n5451 0.000507003
R17904 VSS.n5446 VSS.n5445 0.000507003
R17905 VSS.n5486 VSS.n5485 0.000507003
R17906 VSS.n5440 VSS.n5439 0.000507003
R17907 VSS.n5348 VSS.n5347 0.000507003
R17908 VSS.n5359 VSS.n5358 0.000507003
R17909 VSS.n5338 VSS.n5337 0.000507003
R17910 VSS.n5332 VSS.n5331 0.000507003
R17911 VSS.n5322 VSS.n5321 0.000507003
R17912 VSS.n5318 VSS.n5317 0.000507003
R17913 VSS.n5312 VSS.n5311 0.000507003
R17914 VSS.n5343 VSS.n5342 0.000507003
R17915 VSS.n5302 VSS.n5301 0.000507003
R17916 VSS.n5303 VSS.n5302 0.000507003
R17917 VSS.n5297 VSS.n5296 0.000507003
R17918 VSS.n5290 VSS.n5289 0.000507003
R17919 VSS.n5284 VSS.n5283 0.000507003
R17920 VSS.n5272 VSS.n5271 0.000507003
R17921 VSS.n5266 VSS.n5265 0.000507003
R17922 VSS.n5306 VSS.n5305 0.000507003
R17923 VSS.n5260 VSS.n5259 0.000507003
R17924 VSS.n10082 VSS.n10081 0.000507003
R17925 VSS.n10093 VSS.n10092 0.000507003
R17926 VSS.n10072 VSS.n10071 0.000507003
R17927 VSS.n10066 VSS.n10065 0.000507003
R17928 VSS.n10056 VSS.n10055 0.000507003
R17929 VSS.n10052 VSS.n10051 0.000507003
R17930 VSS.n10046 VSS.n10045 0.000507003
R17931 VSS.n10077 VSS.n10076 0.000507003
R17932 VSS.n4579 VSS.n4578 0.000507003
R17933 VSS.n4583 VSS.n4582 0.000507003
R17934 VSS.n4589 VSS.n4588 0.000507003
R17935 VSS.n4595 VSS.n4594 0.000507003
R17936 VSS.n3811 VSS.n3810 0.000507003
R17937 VSS.n3810 VSS.n3809 0.000507003
R17938 VSS.n3805 VSS.n3804 0.000507003
R17939 VSS.n3799 VSS.n3798 0.000507003
R17940 VSS.n3792 VSS.n3791 0.000507003
R17941 VSS.n3809 VSS.n3792 0.000507003
R17942 VSS.n3787 VSS.n3786 0.000507003
R17943 VSS.n3778 VSS.n3777 0.000507003
R17944 VSS.n3772 VSS.n3771 0.000507003
R17945 VSS.n3762 VSS.n3761 0.000507003
R17946 VSS.n4616 VSS.n4615 0.000507003
R17947 VSS.n4622 VSS.n4621 0.000507003
R17948 VSS.n4629 VSS.n4628 0.000507003
R17949 VSS.n4604 VSS.n4603 0.000507003
R17950 VSS.n6058 VSS.n6057 0.000507003
R17951 VSS.n6066 VSS.n6065 0.000507003
R17952 VSS.n6052 VSS.n6051 0.000507003
R17953 VSS.n6069 VSS.n6068 0.000507003
R17954 VSS.n6082 VSS.n6081 0.000507003
R17955 VSS.n5985 VSS.n5984 0.000507003
R17956 VSS.n5979 VSS.n5978 0.000507003
R17957 VSS.n5974 VSS.n5973 0.000507003
R17958 VSS.n6079 VSS.n5974 0.000507003
R17959 VSS.n6074 VSS.n6073 0.000507003
R17960 VSS.n6179 VSS.n6178 0.000507003
R17961 VSS.n6203 VSS.n6179 0.000507003
R17962 VSS.n6173 VSS.n6172 0.000507003
R17963 VSS.n6163 VSS.n6162 0.000507003
R17964 VSS.n6158 VSS.n6157 0.000507003
R17965 VSS.n11103 VSS.n11102 0.000507003
R17966 VSS.n11097 VSS.n11096 0.000507003
R17967 VSS.n11090 VSS.n11089 0.000507003
R17968 VSS.n11107 VSS.n11090 0.000507003
R17969 VSS.n11085 VSS.n11084 0.000507003
R17970 VSS.n3720 VSS.n3719 0.000507003
R17971 VSS.n11139 VSS.n11138 0.000507003
R17972 VSS.n3724 VSS.n3723 0.000507003
R17973 VSS.n3730 VSS.n3729 0.000507003
R17974 VSS.n3746 VSS.n3745 0.000507003
R17975 VSS.n3752 VSS.n3751 0.000507003
R17976 VSS.n11129 VSS.n11128 0.000507003
R17977 VSS.n11132 VSS.n11131 0.000507003
R17978 VSS.n11069 VSS.n11068 0.000507003
R17979 VSS.n11107 VSS.n11069 0.000507003
R17980 VSS.n11063 VSS.n11062 0.000507003
R17981 VSS.n11110 VSS.n11109 0.000507003
R17982 VSS.n11053 VSS.n11052 0.000507003
R17983 VSS.n6390 VSS.n6347 0.000507003
R17984 VSS.n6387 VSS.n6349 0.000507003
R17985 VSS.n6364 VSS.n6354 0.000507003
R17986 VSS.n6360 VSS.n6355 0.000507003
R17987 VSS.n6341 VSS.n6340 0.000507003
R17988 VSS.n6403 VSS.n6344 0.000507003
R17989 VSS.n6399 VSS.n6345 0.000507003
R17990 VSS.n6395 VSS.n6346 0.000507003
R17991 VSS.n11018 VSS.n3835 0.000507003
R17992 VSS.n11042 VSS.n3835 0.000507003
R17993 VSS.n11015 VSS.n11014 0.000507003
R17994 VSS.n11023 VSS.n11022 0.000507003
R17995 VSS.n11026 VSS.n11025 0.000507003
R17996 VSS.n3860 VSS.n3853 0.000507003
R17997 VSS.n10991 VSS.n3855 0.000507003
R17998 VSS.n3857 VSS.n3856 0.000507003
R17999 VSS.n3869 VSS.n3865 0.000507003
R18000 VSS.n10975 VSS.n10974 0.000507003
R18001 VSS.n10978 VSS.n10970 0.000507003
R18002 VSS.n10982 VSS.n10981 0.000507003
R18003 VSS.n10985 VSS.n10984 0.000507003
R18004 VSS.n10913 VSS.n10912 0.000507003
R18005 VSS.n10913 VSS.n3859 0.000507003
R18006 VSS.n10910 VSS.n10909 0.000507003
R18007 VSS.n10951 VSS.n10916 0.000507003
R18008 VSS.n10947 VSS.n10900 0.000507003
R18009 VSS.n7336 VSS.n7293 0.000507003
R18010 VSS.n7333 VSS.n7295 0.000507003
R18011 VSS.n7310 VSS.n7300 0.000507003
R18012 VSS.n7306 VSS.n7301 0.000507003
R18013 VSS.n7287 VSS.n7286 0.000507003
R18014 VSS.n7349 VSS.n7290 0.000507003
R18015 VSS.n7345 VSS.n7291 0.000507003
R18016 VSS.n7341 VSS.n7292 0.000507003
R18017 VSS.n10867 VSS.n3903 0.000507003
R18018 VSS.n10891 VSS.n3903 0.000507003
R18019 VSS.n10864 VSS.n10863 0.000507003
R18020 VSS.n10872 VSS.n10871 0.000507003
R18021 VSS.n10875 VSS.n10874 0.000507003
R18022 VSS.n3973 VSS.n3972 0.000507003
R18023 VSS.n3978 VSS.n3977 0.000507003
R18024 VSS.n3984 VSS.n3983 0.000507003
R18025 VSS.n3990 VSS.n3989 0.000507003
R18026 VSS.n4006 VSS.n4005 0.000507003
R18027 VSS.n4012 VSS.n4011 0.000507003
R18028 VSS.n4022 VSS.n4021 0.000507003
R18029 VSS.n4017 VSS.n4016 0.000507003
R18030 VSS.n4052 VSS.n4051 0.000507003
R18031 VSS.n4083 VSS.n4052 0.000507003
R18032 VSS.n4046 VSS.n4045 0.000507003
R18033 VSS.n4086 VSS.n4085 0.000507003
R18034 VSS.n4036 VSS.n4035 0.000507003
R18035 VSS.n4150 VSS.n4149 0.000507003
R18036 VSS.n4146 VSS.n4145 0.000507003
R18037 VSS.n4449 VSS.n4132 0.000507003
R18038 VSS.n4449 VSS.n4114 0.000507003
R18039 VSS.n4446 VSS.n4445 0.000507003
R18040 VSS.n4399 VSS.n4398 0.000507003
R18041 VSS.n4395 VSS.n4394 0.000507003
R18042 VSS.n4390 VSS.n4389 0.000507003
R18043 VSS.n4372 VSS.n4186 0.000507003
R18044 VSS.n4405 VSS.n4186 0.000507003
R18045 VSS.n4369 VSS.n4366 0.000507003
R18046 VSS.n4379 VSS.n4377 0.000507003
R18047 VSS.n4375 VSS.n4362 0.000507003
R18048 VSS.n4340 VSS.n4254 0.000507003
R18049 VSS.n4337 VSS.n4334 0.000507003
R18050 VSS.n4266 VSS.n4251 0.000507003
R18051 VSS.n4344 VSS.n4251 0.000507003
R18052 VSS.n4256 VSS.n4255 0.000507003
R18053 VSS.n4303 VSS.n4262 0.000507003
R18054 VSS.n4322 VSS.n4306 0.000507003
R18055 VSS.n4318 VSS.n4307 0.000507003
R18056 VSS.n4315 VSS.n4309 0.000507003
R18057 VSS.n4287 VSS.n4286 0.000507003
R18058 VSS.n4291 VSS.n4290 0.000507003
R18059 VSS.n4296 VSS.n4295 0.000507003
R18060 VSS.n4299 VSS.n4298 0.000507003
R18061 VSS.n4248 VSS.n4247 0.000507003
R18062 VSS.n4344 VSS.n4248 0.000507003
R18063 VSS.n4245 VSS.n4244 0.000507003
R18064 VSS.n4348 VSS.n4232 0.000507003
R18065 VSS.n4233 VSS.n4230 0.000507003
R18066 VSS.n4201 VSS.n4200 0.000507003
R18067 VSS.n4212 VSS.n4211 0.000507003
R18068 VSS.n4223 VSS.n4222 0.000507003
R18069 VSS.n4218 VSS.n4217 0.000507003
R18070 VSS.n4214 VSS.n4187 0.000507003
R18071 VSS.n4404 VSS.n4187 0.000507003
R18072 VSS.n4402 VSS.n4401 0.000507003
R18073 VSS.n4177 VSS.n4171 0.000507003
R18074 VSS.n4174 VSS.n4173 0.000507003
R18075 VSS.n4409 VSS.n4164 0.000507003
R18076 VSS.n4165 VSS.n4162 0.000507003
R18077 VSS.n4415 VSS.n4131 0.000507003
R18078 VSS.n4431 VSS.n4418 0.000507003
R18079 VSS.n4428 VSS.n4419 0.000507003
R18080 VSS.n4425 VSS.n4420 0.000507003
R18081 VSS.n4125 VSS.n4124 0.000507003
R18082 VSS.n10780 VSS.n4110 0.000507003
R18083 VSS.n4112 VSS.n4111 0.000507003
R18084 VSS.n10774 VSS.n10773 0.000507003
R18085 VSS.n10762 VSS.n10761 0.000507003
R18086 VSS.n10762 VSS.n4114 0.000507003
R18087 VSS.n10758 VSS.n10757 0.000507003
R18088 VSS.n10768 VSS.n10767 0.000507003
R18089 VSS.n10770 VSS.n4453 0.000507003
R18090 VSS.n1283 VSS.n1282 0.000507003
R18091 VSS.n1277 VSS.n1276 0.000507003
R18092 VSS.n1299 VSS.n1298 0.000507003
R18093 VSS.n1271 VSS.n1270 0.000507003
R18094 VSS.n789 VSS.n788 0.000507003
R18095 VSS.n790 VSS.n789 0.000507003
R18096 VSS.n783 VSS.n782 0.000507003
R18097 VSS.n777 VSS.n776 0.000507003
R18098 VSS.n682 VSS.n681 0.000507003
R18099 VSS.n790 VSS.n682 0.000507003
R18100 VSS.n793 VSS.n792 0.000507003
R18101 VSS.n677 VSS.n676 0.000507003
R18102 VSS.n671 VSS.n670 0.000507003
R18103 VSS.n661 VSS.n660 0.000507003
R18104 VSS.n1261 VSS.n1260 0.000507003
R18105 VSS.n1255 VSS.n1254 0.000507003
R18106 VSS.n1266 VSS.n1265 0.000507003
R18107 VSS.n1292 VSS.n1291 0.000507003
R18108 VSS.n1221 VSS.n1220 0.000507003
R18109 VSS.n1227 VSS.n1226 0.000507003
R18110 VSS.n1335 VSS.n1334 0.000507003
R18111 VSS.n1340 VSS.n1339 0.000507003
R18112 VSS.n1046 VSS.n1045 0.000507003
R18113 VSS.n1047 VSS.n1046 0.000507003
R18114 VSS.n1041 VSS.n1040 0.000507003
R18115 VSS.n1034 VSS.n1033 0.000507003
R18116 VSS.n1028 VSS.n1027 0.000507003
R18117 VSS.n1016 VSS.n1015 0.000507003
R18118 VSS.n1010 VSS.n1009 0.000507003
R18119 VSS.n1050 VSS.n1049 0.000507003
R18120 VSS.n1004 VSS.n1003 0.000507003
R18121 VSS.n1209 VSS.n1208 0.000507003
R18122 VSS.n1203 VSS.n1202 0.000507003
R18123 VSS.n1343 VSS.n1342 0.000507003
R18124 VSS.n1350 VSS.n1349 0.000507003
R18125 VSS.n969 VSS.n968 0.000507003
R18126 VSS.n975 VSS.n974 0.000507003
R18127 VSS.n1085 VSS.n1084 0.000507003
R18128 VSS.n14331 VSS.n14330 0.000507003
R18129 VSS.n14332 VSS.n14331 0.000507003
R18130 VSS.n14325 VSS.n14324 0.000507003
R18131 VSS.n14315 VSS.n14314 0.000507003
R18132 VSS.n14310 VSS.n14309 0.000507003
R18133 VSS.n14223 VSS.n14222 0.000507003
R18134 VSS.n14219 VSS.n14218 0.000507003
R18135 VSS.n14214 VSS.n14213 0.000507003
R18136 VSS.n568 VSS.n567 0.000507003
R18137 VSS.n14229 VSS.n568 0.000507003
R18138 VSS.n565 VSS.n562 0.000507003
R18139 VSS.n549 VSS.n545 0.000507003
R18140 VSS.n14233 VSS.n14232 0.000507003
R18141 VSS.n10691 VSS.n10690 0.000507003
R18142 VSS.n10707 VSS.n10706 0.000507003
R18143 VSS.n10686 VSS.n10685 0.000507003
R18144 VSS.n10680 VSS.n10679 0.000507003
R18145 VSS.n14274 VSS.n14273 0.000507003
R18146 VSS.n14275 VSS.n14274 0.000507003
R18147 VSS.n14268 VSS.n14267 0.000507003
R18148 VSS.n14278 VSS.n14277 0.000507003
R18149 VSS.n14261 VSS.n14260 0.000507003
R18150 VSS.n14275 VSS.n14261 0.000507003
R18151 VSS.n14256 VSS.n14255 0.000507003
R18152 VSS.n532 VSS.n531 0.000507003
R18153 VSS.n526 VSS.n525 0.000507003
R18154 VSS.n516 VSS.n515 0.000507003
R18155 VSS.n10667 VSS.n10666 0.000507003
R18156 VSS.n10661 VSS.n10660 0.000507003
R18157 VSS.n10672 VSS.n10671 0.000507003
R18158 VSS.n10700 VSS.n10699 0.000507003
R18159 VSS.n14201 VSS.n584 0.000507003
R18160 VSS.n14205 VSS.n14204 0.000507003
R18161 VSS.n600 VSS.n599 0.000507003
R18162 VSS.n597 VSS.n596 0.000507003
R18163 VSS.n1147 VSS.n1146 0.000507003
R18164 VSS.n1143 VSS.n1142 0.000507003
R18165 VSS.n1139 VSS.n1138 0.000507003
R18166 VSS.n929 VSS.n910 0.000507003
R18167 VSS.n1151 VSS.n929 0.000507003
R18168 VSS.n1155 VSS.n1154 0.000507003
R18169 VSS.n919 VSS.n914 0.000507003
R18170 VSS.n924 VSS.n918 0.000507003
R18171 VSS.n1135 VSS.n1134 0.000507003
R18172 VSS.n14191 VSS.n14179 0.000507003
R18173 VSS.n14188 VSS.n14187 0.000507003
R18174 VSS.n14197 VSS.n606 0.000507003
R18175 VSS.n14195 VSS.n14178 0.000507003
R18176 VSS.n12447 VSS.n12446 0.000507003
R18177 VSS.n12441 VSS.n12440 0.000507003
R18178 VSS.n12435 VSS.n12434 0.000507003
R18179 VSS.n12391 VSS.n12390 0.000507003
R18180 VSS.n12414 VSS.n2480 0.000507003
R18181 VSS.n12418 VSS.n12417 0.000507003
R18182 VSS.n12411 VSS.n12410 0.000507003
R18183 VSS.n12408 VSS.n12407 0.000507003
R18184 VSS.n13044 VSS.n13043 0.000507003
R18185 VSS.n13045 VSS.n13044 0.000507003
R18186 VSS.n13039 VSS.n13038 0.000507003
R18187 VSS.n13035 VSS.n13034 0.000507003
R18188 VSS.n13046 VSS.n2481 0.000507003
R18189 VSS.n13046 VSS.n13045 0.000507003
R18190 VSS.n2535 VSS.n2534 0.000507003
R18191 VSS.n2546 VSS.n2545 0.000507003
R18192 VSS.n2542 VSS.n2538 0.000507003
R18193 VSS.n2486 VSS.n2482 0.000507003
R18194 VSS.n2476 VSS.n2475 0.000507003
R18195 VSS.n2473 VSS.n2470 0.000507003
R18196 VSS.n13053 VSS.n2461 0.000507003
R18197 VSS.n13057 VSS.n13056 0.000507003
R18198 VSS.n2452 VSS.n2392 0.000507003
R18199 VSS.n2448 VSS.n2393 0.000507003
R18200 VSS.n2444 VSS.n2443 0.000507003
R18201 VSS.n2438 VSS.n2437 0.000507003
R18202 VSS.n13100 VSS.n13099 0.000507003
R18203 VSS.n13101 VSS.n13100 0.000507003
R18204 VSS.n13104 VSS.n13103 0.000507003
R18205 VSS.n2369 VSS.n2368 0.000507003
R18206 VSS.n2391 VSS.n2363 0.000507003
R18207 VSS.n13101 VSS.n2363 0.000507003
R18208 VSS.n2389 VSS.n2375 0.000507003
R18209 VSS.n2386 VSS.n2385 0.000507003
R18210 VSS.n2381 VSS.n2378 0.000507003
R18211 VSS.n13097 VSS.n2372 0.000507003
R18212 VSS.n13085 VSS.n13073 0.000507003
R18213 VSS.n13082 VSS.n13081 0.000507003
R18214 VSS.n13091 VSS.n2457 0.000507003
R18215 VSS.n13089 VSS.n13072 0.000507003
R18216 VSS.n13133 VSS.n1911 0.000507003
R18217 VSS.n13137 VSS.n13136 0.000507003
R18218 VSS.n1920 VSS.n1919 0.000507003
R18219 VSS.n1924 VSS.n1918 0.000507003
R18220 VSS.n2338 VSS.n2337 0.000507003
R18221 VSS.n2334 VSS.n2333 0.000507003
R18222 VSS.n2330 VSS.n2329 0.000507003
R18223 VSS.n2343 VSS.n1929 0.000507003
R18224 VSS.n2343 VSS.n2342 0.000507003
R18225 VSS.n2295 VSS.n2294 0.000507003
R18226 VSS.n2291 VSS.n2290 0.000507003
R18227 VSS.n2287 VSS.n2286 0.000507003
R18228 VSS.n1934 VSS.n1930 0.000507003
R18229 VSS.n13121 VSS.n13120 0.000507003
R18230 VSS.n13117 VSS.n13116 0.000507003
R18231 VSS.n13129 VSS.n13128 0.000507003
R18232 VSS.n13126 VSS.n13125 0.000507003
R18233 VSS.n14157 VSS.n14156 0.000507003
R18234 VSS.n14160 VSS.n14159 0.000507003
R18235 VSS.n14171 VSS.n14170 0.000507003
R18236 VSS.n14166 VSS.n14165 0.000507003
R18237 VSS.n14162 VSS.n569 0.000507003
R18238 VSS.n14228 VSS.n569 0.000507003
R18239 VSS.n14226 VSS.n14225 0.000507003
R18240 VSS.n2415 VSS.n554 0.000507003
R18241 VSS.n14229 VSS.n554 0.000507003
R18242 VSS.n2412 VSS.n2411 0.000507003
R18243 VSS.n2403 VSS.n2402 0.000507003
R18244 VSS.n2418 VSS.n2406 0.000507003
R18245 VSS.n1166 VSS.n881 0.000507003
R18246 VSS.n1166 VSS.n1165 0.000507003
R18247 VSS.n1163 VSS.n1162 0.000507003
R18248 VSS.n907 VSS.n899 0.000507003
R18249 VSS.n904 VSS.n900 0.000507003
R18250 VSS.n943 VSS.n942 0.000507003
R18251 VSS.n947 VSS.n946 0.000507003
R18252 VSS.n953 VSS.n952 0.000507003
R18253 VSS.n886 VSS.n882 0.000507003
R18254 VSS.n1395 VSS.n862 0.000507003
R18255 VSS.n1399 VSS.n1398 0.000507003
R18256 VSS.n871 VSS.n870 0.000507003
R18257 VSS.n875 VSS.n869 0.000507003
R18258 VSS.n1381 VSS.n1373 0.000507003
R18259 VSS.n1385 VSS.n1372 0.000507003
R18260 VSS.n1389 VSS.n1388 0.000507003
R18261 VSS.n1391 VSS.n1171 0.000507003
R18262 VSS.n959 VSS.n958 0.000507003
R18263 VSS.n1111 VSS.n1110 0.000507003
R18264 VSS.n1089 VSS.n1088 0.000507003
R18265 VSS.n1095 VSS.n1094 0.000507003
R18266 VSS.n1104 VSS.n1103 0.000507003
R18267 VSS.n14296 VSS.n14295 0.000507003
R18268 VSS.n14290 VSS.n14289 0.000507003
R18269 VSS.n14335 VSS.n14334 0.000507003
R18270 VSS.n14284 VSS.n14283 0.000507003
R18271 VSS.n1568 VSS.n1567 0.000507003
R18272 VSS.n1569 VSS.n1568 0.000507003
R18273 VSS.n1563 VSS.n1562 0.000507003
R18274 VSS.n1556 VSS.n1555 0.000507003
R18275 VSS.n1550 VSS.n1549 0.000507003
R18276 VSS.n1538 VSS.n1537 0.000507003
R18277 VSS.n1532 VSS.n1531 0.000507003
R18278 VSS.n1572 VSS.n1571 0.000507003
R18279 VSS.n1526 VSS.n1525 0.000507003
R18280 VSS.n13713 VSS.n13712 0.000507003
R18281 VSS.n13858 VSS.n13857 0.000507003
R18282 VSS.n13722 VSS.n13721 0.000507003
R18283 VSS.n13728 VSS.n13727 0.000507003
R18284 VSS.n13710 VSS.n13709 0.000507003
R18285 VSS.n13738 VSS.n13737 0.000507003
R18286 VSS.n13847 VSS.n13846 0.000507003
R18287 VSS.n13718 VSS.n13717 0.000507003
R18288 VSS.n13808 VSS.n13807 0.000507003
R18289 VSS.n13809 VSS.n13808 0.000507003
R18290 VSS.n13803 VSS.n13802 0.000507003
R18291 VSS.n13796 VSS.n13795 0.000507003
R18292 VSS.n13790 VSS.n13789 0.000507003
R18293 VSS.n13778 VSS.n13777 0.000507003
R18294 VSS.n13772 VSS.n13771 0.000507003
R18295 VSS.n13812 VSS.n13811 0.000507003
R18296 VSS.n13766 VSS.n13765 0.000507003
R18297 VSS.n13393 VSS.n13392 0.000507003
R18298 VSS.n13259 VSS.n13258 0.000507003
R18299 VSS.n13265 VSS.n13264 0.000507003
R18300 VSS.n13253 VSS.n13252 0.000507003
R18301 VSS.n13247 VSS.n13246 0.000507003
R18302 VSS.n13275 VSS.n13274 0.000507003
R18303 VSS.n13382 VSS.n13381 0.000507003
R18304 VSS.n13250 VSS.n13249 0.000507003
R18305 VSS.n1490 VSS.n1489 0.000507003
R18306 VSS.n1496 VSS.n1495 0.000507003
R18307 VSS.n1606 VSS.n1605 0.000507003
R18308 VSS.n1611 VSS.n1610 0.000507003
R18309 VSS.n761 VSS.n760 0.000507003
R18310 VSS.n762 VSS.n761 0.000507003
R18311 VSS.n756 VSS.n755 0.000507003
R18312 VSS.n749 VSS.n748 0.000507003
R18313 VSS.n743 VSS.n742 0.000507003
R18314 VSS.n731 VSS.n730 0.000507003
R18315 VSS.n725 VSS.n724 0.000507003
R18316 VSS.n765 VSS.n764 0.000507003
R18317 VSS.n719 VSS.n718 0.000507003
R18318 VSS.n1478 VSS.n1477 0.000507003
R18319 VSS.n1472 VSS.n1471 0.000507003
R18320 VSS.n1614 VSS.n1613 0.000507003
R18321 VSS.n1621 VSS.n1620 0.000507003
R18322 VSS.n14114 VSS.n628 0.000507003
R18323 VSS.n14115 VSS.n14114 0.000507003
R18324 VSS.n14119 VSS.n630 0.000507003
R18325 VSS.n632 VSS.n631 0.000507003
R18326 VSS.n645 VSS.n640 0.000507003
R18327 VSS.n1448 VSS.n1447 0.000507003
R18328 VSS.n1452 VSS.n1451 0.000507003
R18329 VSS.n1457 VSS.n1456 0.000507003
R18330 VSS.n1460 VSS.n1459 0.000507003
R18331 VSS.n1690 VSS.n1684 0.000507003
R18332 VSS.n1694 VSS.n1693 0.000507003
R18333 VSS.n1681 VSS.n1680 0.000507003
R18334 VSS.n1686 VSS.n1461 0.000507003
R18335 VSS.n14098 VSS.n14090 0.000507003
R18336 VSS.n14102 VSS.n14089 0.000507003
R18337 VSS.n14106 VSS.n14105 0.000507003
R18338 VSS.n14108 VSS.n1465 0.000507003
R18339 VSS.n13694 VSS.n13693 0.000507003
R18340 VSS.n13691 VSS.n13673 0.000507003
R18341 VSS.n13687 VSS.n13674 0.000507003
R18342 VSS.n13684 VSS.n13683 0.000507003
R18343 VSS.n13680 VSS.n13676 0.000507003
R18344 VSS.n13680 VSS.n1661 0.000507003
R18345 VSS.n14078 VSS.n14077 0.000507003
R18346 VSS.n14079 VSS.n14078 0.000507003
R18347 VSS.n14075 VSS.n14061 0.000507003
R18348 VSS.n14072 VSS.n14062 0.000507003
R18349 VSS.n14069 VSS.n14066 0.000507003
R18350 VSS.n1653 VSS.n1652 0.000507003
R18351 VSS.n14083 VSS.n1643 0.000507003
R18352 VSS.n1645 VSS.n1644 0.000507003
R18353 VSS.n1667 VSS.n1666 0.000507003
R18354 VSS.n13665 VSS.n13664 0.000507003
R18355 VSS.n13662 VSS.n13661 0.000507003
R18356 VSS.n13701 VSS.n13668 0.000507003
R18357 VSS.n13698 VSS.n13652 0.000507003
R18358 VSS.n13903 VSS.n13204 0.000507003
R18359 VSS.n13907 VSS.n13906 0.000507003
R18360 VSS.n13213 VSS.n13212 0.000507003
R18361 VSS.n13217 VSS.n13211 0.000507003
R18362 VSS.n13642 VSS.n13641 0.000507003
R18363 VSS.n13643 VSS.n13642 0.000507003
R18364 VSS.n13637 VSS.n13636 0.000507003
R18365 VSS.n13633 VSS.n13632 0.000507003
R18366 VSS.n13644 VSS.n13222 0.000507003
R18367 VSS.n13644 VSS.n13643 0.000507003
R18368 VSS.n13534 VSS.n13533 0.000507003
R18369 VSS.n13545 VSS.n13544 0.000507003
R18370 VSS.n13541 VSS.n13537 0.000507003
R18371 VSS.n13227 VSS.n13223 0.000507003
R18372 VSS.n13887 VSS.n13886 0.000507003
R18373 VSS.n13891 VSS.n13890 0.000507003
R18374 VSS.n13896 VSS.n13895 0.000507003
R18375 VSS.n13899 VSS.n13898 0.000507003
R18376 VSS.n830 VSS.n829 0.000507003
R18377 VSS.n833 VSS.n832 0.000507003
R18378 VSS.n1438 VSS.n1437 0.000507003
R18379 VSS.n835 VSS.n813 0.000507003
R18380 VSS.n1410 VSS.n840 0.000507003
R18381 VSS.n1410 VSS.n818 0.000507003
R18382 VSS.n1407 VSS.n1406 0.000507003
R18383 VSS.n859 VSS.n849 0.000507003
R18384 VSS.n855 VSS.n850 0.000507003
R18385 VSS.n1183 VSS.n1176 0.000507003
R18386 VSS.n1187 VSS.n1186 0.000507003
R18387 VSS.n1194 VSS.n1193 0.000507003
R18388 VSS.n1190 VSS.n841 0.000507003
R18389 VSS.n1427 VSS.n1426 0.000507003
R18390 VSS.n1422 VSS.n1421 0.000507003
R18391 VSS.n1416 VSS.n839 0.000507003
R18392 VSS.n1431 VSS.n838 0.000507003
R18393 VSS.n2210 VSS.n2054 0.000507003
R18394 VSS.n2207 VSS.n2055 0.000507003
R18395 VSS.n2203 VSS.n2202 0.000507003
R18396 VSS.n2199 VSS.n2193 0.000507003
R18397 VSS.n2195 VSS.n2194 0.000507003
R18398 VSS.n2194 VSS.n2005 0.000507003
R18399 VSS.n2244 VSS.n1983 0.000507003
R18400 VSS.n2245 VSS.n2244 0.000507003
R18401 VSS.n2249 VSS.n1985 0.000507003
R18402 VSS.n1987 VSS.n1986 0.000507003
R18403 VSS.n2000 VSS.n1995 0.000507003
R18404 VSS.n2042 VSS.n2041 0.000507003
R18405 VSS.n2046 VSS.n2045 0.000507003
R18406 VSS.n2051 VSS.n2050 0.000507003
R18407 VSS.n2053 VSS.n2008 0.000507003
R18408 VSS.n2230 VSS.n2229 0.000507003
R18409 VSS.n2226 VSS.n2225 0.000507003
R18410 VSS.n2236 VSS.n2235 0.000507003
R18411 VSS.n2238 VSS.n2215 0.000507003
R18412 VSS.n2126 VSS.n2103 0.000507003
R18413 VSS.n2123 VSS.n2104 0.000507003
R18414 VSS.n2119 VSS.n2105 0.000507003
R18415 VSS.n2115 VSS.n2107 0.000507003
R18416 VSS.n2113 VSS.n2112 0.000507003
R18417 VSS.n2112 VSS.n2080 0.000507003
R18418 VSS.n2179 VSS.n2058 0.000507003
R18419 VSS.n2180 VSS.n2179 0.000507003
R18420 VSS.n2184 VSS.n2060 0.000507003
R18421 VSS.n2062 VSS.n2061 0.000507003
R18422 VSS.n2075 VSS.n2070 0.000507003
R18423 VSS.n2091 VSS.n2090 0.000507003
R18424 VSS.n2095 VSS.n2094 0.000507003
R18425 VSS.n2100 VSS.n2099 0.000507003
R18426 VSS.n2102 VSS.n2083 0.000507003
R18427 VSS.n2165 VSS.n2164 0.000507003
R18428 VSS.n2161 VSS.n2160 0.000507003
R18429 VSS.n2171 VSS.n2170 0.000507003
R18430 VSS.n2173 VSS.n2131 0.000507003
R18431 VSS.n12649 VSS.n1851 0.000507003
R18432 VSS.n12653 VSS.n12652 0.000507003
R18433 VSS.n12666 VSS.n12665 0.000507003
R18434 VSS.n12662 VSS.n12656 0.000507003
R18435 VSS.n12658 VSS.n12657 0.000507003
R18436 VSS.n12657 VSS.n1849 0.000507003
R18437 VSS.n13189 VSS.n1852 0.000507003
R18438 VSS.n13189 VSS.n13188 0.000507003
R18439 VSS.n13186 VSS.n13185 0.000507003
R18440 VSS.n1878 VSS.n1870 0.000507003
R18441 VSS.n1875 VSS.n1871 0.000507003
R18442 VSS.n2138 VSS.n2137 0.000507003
R18443 VSS.n2148 VSS.n2141 0.000507003
R18444 VSS.n2145 VSS.n2142 0.000507003
R18445 VSS.n1857 VSS.n1853 0.000507003
R18446 VSS.n1846 VSS.n1845 0.000507003
R18447 VSS.n1843 VSS.n1842 0.000507003
R18448 VSS.n13199 VSS.n1833 0.000507003
R18449 VSS.n13196 VSS.n1831 0.000507003
R18450 VSS.n12687 VSS.n1813 0.000507003
R18451 VSS.n12691 VSS.n12690 0.000507003
R18452 VSS.n12683 VSS.n12682 0.000507003
R18453 VSS.n12680 VSS.n12679 0.000507003
R18454 VSS.n13934 VSS.n13933 0.000507003
R18455 VSS.n13935 VSS.n13934 0.000507003
R18456 VSS.n13938 VSS.n13937 0.000507003
R18457 VSS.n1790 VSS.n1789 0.000507003
R18458 VSS.n1812 VSS.n1784 0.000507003
R18459 VSS.n13935 VSS.n1784 0.000507003
R18460 VSS.n1810 VSS.n1796 0.000507003
R18461 VSS.n1807 VSS.n1806 0.000507003
R18462 VSS.n1802 VSS.n1799 0.000507003
R18463 VSS.n13931 VSS.n1793 0.000507003
R18464 VSS.n1828 VSS.n1827 0.000507003
R18465 VSS.n13917 VSS.n1820 0.000507003
R18466 VSS.n13920 VSS.n13919 0.000507003
R18467 VSS.n13925 VSS.n13924 0.000507003
R18468 VSS.n2021 VSS.n2020 0.000507003
R18469 VSS.n2024 VSS.n2023 0.000507003
R18470 VSS.n2032 VSS.n2031 0.000507003
R18471 VSS.n2028 VSS.n1977 0.000507003
R18472 VSS.n2318 VSS.n2317 0.000507003
R18473 VSS.n2319 VSS.n2318 0.000507003
R18474 VSS.n2315 VSS.n2314 0.000507003
R18475 VSS.n2311 VSS.n2310 0.000507003
R18476 VSS.n2306 VSS.n2305 0.000507003
R18477 VSS.n1967 VSS.n1948 0.000507003
R18478 VSS.n2319 VSS.n1967 0.000507003
R18479 VSS.n2322 VSS.n2321 0.000507003
R18480 VSS.n1965 VSS.n1964 0.000507003
R18481 VSS.n1962 VSS.n1959 0.000507003
R18482 VSS.n2268 VSS.n2267 0.000507003
R18483 VSS.n2264 VSS.n2263 0.000507003
R18484 VSS.n2276 VSS.n1980 0.000507003
R18485 VSS.n2274 VSS.n2273 0.000507003
R18486 VSS.n12984 VSS.n2562 0.000507003
R18487 VSS.n12985 VSS.n12984 0.000507003
R18488 VSS.n12989 VSS.n2564 0.000507003
R18489 VSS.n2566 VSS.n2565 0.000507003
R18490 VSS.n2579 VSS.n2574 0.000507003
R18491 VSS.n2649 VSS.n2648 0.000507003
R18492 VSS.n2653 VSS.n2652 0.000507003
R18493 VSS.n2658 VSS.n2657 0.000507003
R18494 VSS.n2660 VSS.n2587 0.000507003
R18495 VSS.n2717 VSS.n2661 0.000507003
R18496 VSS.n2721 VSS.n2720 0.000507003
R18497 VSS.n2713 VSS.n2712 0.000507003
R18498 VSS.n2710 VSS.n2709 0.000507003
R18499 VSS.n12966 VSS.n12965 0.000507003
R18500 VSS.n12970 VSS.n12969 0.000507003
R18501 VSS.n12976 VSS.n12975 0.000507003
R18502 VSS.n12978 VSS.n2665 0.000507003
R18503 VSS.n12948 VSS.n12947 0.000507003
R18504 VSS.n12949 VSS.n12948 0.000507003
R18505 VSS.n12945 VSS.n12931 0.000507003
R18506 VSS.n12942 VSS.n12932 0.000507003
R18507 VSS.n12939 VSS.n12936 0.000507003
R18508 VSS.n2680 VSS.n2679 0.000507003
R18509 VSS.n12953 VSS.n2670 0.000507003
R18510 VSS.n2672 VSS.n2671 0.000507003
R18511 VSS.n2694 VSS.n2693 0.000507003
R18512 VSS.n2811 VSS.n2810 0.000507003
R18513 VSS.n2807 VSS.n2806 0.000507003
R18514 VSS.n2804 VSS.n2792 0.000507003
R18515 VSS.n2801 VSS.n2800 0.000507003
R18516 VSS.n2780 VSS.n2775 0.000507003
R18517 VSS.n2783 VSS.n2782 0.000507003
R18518 VSS.n2819 VSS.n2786 0.000507003
R18519 VSS.n2815 VSS.n2770 0.000507003
R18520 VSS.n12907 VSS.n2743 0.000507003
R18521 VSS.n12908 VSS.n12907 0.000507003
R18522 VSS.n12912 VSS.n2745 0.000507003
R18523 VSS.n2747 VSS.n2746 0.000507003
R18524 VSS.n2760 VSS.n2755 0.000507003
R18525 VSS.n2830 VSS.n2829 0.000507003
R18526 VSS.n2834 VSS.n2833 0.000507003
R18527 VSS.n2839 VSS.n2838 0.000507003
R18528 VSS.n2841 VSS.n2768 0.000507003
R18529 VSS.n2897 VSS.n2842 0.000507003
R18530 VSS.n2901 VSS.n2900 0.000507003
R18531 VSS.n2893 VSS.n2892 0.000507003
R18532 VSS.n2890 VSS.n2889 0.000507003
R18533 VSS.n12889 VSS.n12888 0.000507003
R18534 VSS.n12893 VSS.n12892 0.000507003
R18535 VSS.n12899 VSS.n12898 0.000507003
R18536 VSS.n12901 VSS.n2846 0.000507003
R18537 VSS.n12635 VSS.n12634 0.000507003
R18538 VSS.n12632 VSS.n3057 0.000507003
R18539 VSS.n12628 VSS.n3058 0.000507003
R18540 VSS.n12625 VSS.n12624 0.000507003
R18541 VSS.n12621 VSS.n12617 0.000507003
R18542 VSS.n12621 VSS.n2868 0.000507003
R18543 VSS.n12871 VSS.n12870 0.000507003
R18544 VSS.n12872 VSS.n12871 0.000507003
R18545 VSS.n12868 VSS.n12854 0.000507003
R18546 VSS.n12865 VSS.n12855 0.000507003
R18547 VSS.n12862 VSS.n12859 0.000507003
R18548 VSS.n2860 VSS.n2859 0.000507003
R18549 VSS.n12876 VSS.n2850 0.000507003
R18550 VSS.n2852 VSS.n2851 0.000507003
R18551 VSS.n2874 VSS.n2873 0.000507003
R18552 VSS.n3049 VSS.n3048 0.000507003
R18553 VSS.n3046 VSS.n3045 0.000507003
R18554 VSS.n12642 VSS.n3052 0.000507003
R18555 VSS.n12639 VSS.n3036 0.000507003
R18556 VSS.n3078 VSS.n3018 0.000507003
R18557 VSS.n3082 VSS.n3081 0.000507003
R18558 VSS.n3074 VSS.n3073 0.000507003
R18559 VSS.n3071 VSS.n3070 0.000507003
R18560 VSS.n12729 VSS.n12728 0.000507003
R18561 VSS.n12730 VSS.n12729 0.000507003
R18562 VSS.n12733 VSS.n12732 0.000507003
R18563 VSS.n2968 VSS.n2967 0.000507003
R18564 VSS.n3017 VSS.n2962 0.000507003
R18565 VSS.n12730 VSS.n2962 0.000507003
R18566 VSS.n3015 VSS.n3001 0.000507003
R18567 VSS.n3012 VSS.n3011 0.000507003
R18568 VSS.n3007 VSS.n3004 0.000507003
R18569 VSS.n12726 VSS.n2971 0.000507003
R18570 VSS.n3033 VSS.n3032 0.000507003
R18571 VSS.n12712 VSS.n3025 0.000507003
R18572 VSS.n12715 VSS.n12714 0.000507003
R18573 VSS.n12720 VSS.n12719 0.000507003
R18574 VSS.n2601 VSS.n2600 0.000507003
R18575 VSS.n2604 VSS.n2603 0.000507003
R18576 VSS.n2639 VSS.n2638 0.000507003
R18577 VSS.n2635 VSS.n2590 0.000507003
R18578 VSS.n13023 VSS.n13022 0.000507003
R18579 VSS.n13024 VSS.n13023 0.000507003
R18580 VSS.n13020 VSS.n13019 0.000507003
R18581 VSS.n13016 VSS.n13015 0.000507003
R18582 VSS.n13011 VSS.n13010 0.000507003
R18583 VSS.n2519 VSS.n2500 0.000507003
R18584 VSS.n13024 VSS.n2519 0.000507003
R18585 VSS.n13027 VSS.n13026 0.000507003
R18586 VSS.n2517 VSS.n2516 0.000507003
R18587 VSS.n2514 VSS.n2511 0.000507003
R18588 VSS.n2623 VSS.n2622 0.000507003
R18589 VSS.n2619 VSS.n2618 0.000507003
R18590 VSS.n2631 VSS.n2608 0.000507003
R18591 VSS.n2629 VSS.n2628 0.000507003
R18592 VSS.n11675 VSS.n11674 0.000507003
R18593 VSS.n11676 VSS.n11675 0.000507003
R18594 VSS.n11679 VSS.n11678 0.000507003
R18595 VSS.n11670 VSS.n11669 0.000507003
R18596 VSS.n11664 VSS.n11663 0.000507003
R18597 VSS.n11652 VSS.n11651 0.000507003
R18598 VSS.n11646 VSS.n11645 0.000507003
R18599 VSS.n11640 VSS.n11639 0.000507003
R18600 VSS.n11578 VSS.n11577 0.000507003
R18601 VSS.n12250 VSS.n12249 0.000507003
R18602 VSS.n12261 VSS.n12260 0.000507003
R18603 VSS.n12240 VSS.n12239 0.000507003
R18604 VSS.n12234 VSS.n12233 0.000507003
R18605 VSS.n12224 VSS.n12223 0.000507003
R18606 VSS.n12220 VSS.n12219 0.000507003
R18607 VSS.n12214 VSS.n12213 0.000507003
R18608 VSS.n12245 VSS.n12244 0.000507003
R18609 VSS.n11744 VSS.n11743 0.000507003
R18610 VSS.n11745 VSS.n11744 0.000507003
R18611 VSS.n11748 VSS.n11747 0.000507003
R18612 VSS.n11739 VSS.n11738 0.000507003
R18613 VSS.n11733 VSS.n11732 0.000507003
R18614 VSS.n11721 VSS.n11720 0.000507003
R18615 VSS.n11715 VSS.n11714 0.000507003
R18616 VSS.n11709 VSS.n11708 0.000507003
R18617 VSS.n11702 VSS.n11701 0.000507003
R18618 VSS.n12143 VSS.n12142 0.000507003
R18619 VSS.n12154 VSS.n12153 0.000507003
R18620 VSS.n12133 VSS.n12132 0.000507003
R18621 VSS.n12127 VSS.n12126 0.000507003
R18622 VSS.n12117 VSS.n12116 0.000507003
R18623 VSS.n12113 VSS.n12112 0.000507003
R18624 VSS.n12107 VSS.n12106 0.000507003
R18625 VSS.n12138 VSS.n12137 0.000507003
R18626 VSS.n12097 VSS.n12096 0.000507003
R18627 VSS.n12098 VSS.n12097 0.000507003
R18628 VSS.n12092 VSS.n12091 0.000507003
R18629 VSS.n12085 VSS.n12084 0.000507003
R18630 VSS.n12079 VSS.n12078 0.000507003
R18631 VSS.n12067 VSS.n12066 0.000507003
R18632 VSS.n12061 VSS.n12060 0.000507003
R18633 VSS.n12101 VSS.n12100 0.000507003
R18634 VSS.n12055 VSS.n12054 0.000507003
R18635 VSS.n11975 VSS.n11974 0.000507003
R18636 VSS.n11986 VSS.n11985 0.000507003
R18637 VSS.n11965 VSS.n11964 0.000507003
R18638 VSS.n11959 VSS.n11958 0.000507003
R18639 VSS.n11949 VSS.n11948 0.000507003
R18640 VSS.n11945 VSS.n11944 0.000507003
R18641 VSS.n11939 VSS.n11938 0.000507003
R18642 VSS.n11970 VSS.n11969 0.000507003
R18643 VSS.n11876 VSS.n11875 0.000507003
R18644 VSS.n11877 VSS.n11876 0.000507003
R18645 VSS.n11880 VSS.n11879 0.000507003
R18646 VSS.n11871 VSS.n11870 0.000507003
R18647 VSS.n11865 VSS.n11864 0.000507003
R18648 VSS.n11853 VSS.n11852 0.000507003
R18649 VSS.n11847 VSS.n11846 0.000507003
R18650 VSS.n11841 VSS.n11840 0.000507003
R18651 VSS.n11834 VSS.n11833 0.000507003
R18652 VSS.n3547 VSS.n3546 0.000507003
R18653 VSS.n3558 VSS.n3557 0.000507003
R18654 VSS.n3537 VSS.n3536 0.000507003
R18655 VSS.n3531 VSS.n3530 0.000507003
R18656 VSS.n3521 VSS.n3520 0.000507003
R18657 VSS.n3517 VSS.n3516 0.000507003
R18658 VSS.n3511 VSS.n3510 0.000507003
R18659 VSS.n3542 VSS.n3541 0.000507003
R18660 VSS.n3501 VSS.n3500 0.000507003
R18661 VSS.n3502 VSS.n3501 0.000507003
R18662 VSS.n3496 VSS.n3495 0.000507003
R18663 VSS.n3489 VSS.n3488 0.000507003
R18664 VSS.n3483 VSS.n3482 0.000507003
R18665 VSS.n3471 VSS.n3470 0.000507003
R18666 VSS.n3465 VSS.n3464 0.000507003
R18667 VSS.n3505 VSS.n3504 0.000507003
R18668 VSS.n3459 VSS.n3458 0.000507003
R18669 VSS.n12599 VSS.n12598 0.000507003
R18670 VSS.n12589 VSS.n12588 0.000507003
R18671 VSS.n3112 VSS.n3111 0.000507003
R18672 VSS.n3106 VSS.n3105 0.000507003
R18673 VSS.n3096 VSS.n3095 0.000507003
R18674 VSS.n3092 VSS.n3091 0.000507003
R18675 VSS.n12608 VSS.n12607 0.000507003
R18676 VSS.n12594 VSS.n12593 0.000507003
R18677 VSS.n3119 VSS.n3118 0.000507003
R18678 VSS.n3169 VSS.n3168 0.000507003
R18679 VSS.n3123 VSS.n3122 0.000507003
R18680 VSS.n3129 VSS.n3128 0.000507003
R18681 VSS.n3261 VSS.n3260 0.000507003
R18682 VSS.n3255 VSS.n3254 0.000507003
R18683 VSS.n3270 VSS.n3269 0.000507003
R18684 VSS.n3252 VSS.n3251 0.000507003
R18685 VSS.n3267 VSS.n3252 0.000507003
R18686 VSS.n3247 VSS.n3246 0.000507003
R18687 VSS.n3240 VSS.n3239 0.000507003
R18688 VSS.n3234 VSS.n3233 0.000507003
R18689 VSS.n3224 VSS.n3223 0.000507003
R18690 VSS.n3150 VSS.n3149 0.000507003
R18691 VSS.n3156 VSS.n3155 0.000507003
R18692 VSS.n3160 VSS.n3159 0.000507003
R18693 VSS.n3138 VSS.n3137 0.000507003
R18694 VSS.n11608 VSS.n11607 0.000507003
R18695 VSS.n11616 VSS.n11615 0.000507003
R18696 VSS.n11634 VSS.n11633 0.000507003
R18697 VSS.n11619 VSS.n11618 0.000507003
R18698 VSS.n11600 VSS.n11599 0.000507003
R18699 VSS.n11594 VSS.n11593 0.000507003
R18700 VSS.n11588 VSS.n11587 0.000507003
R18701 VSS.n11583 VSS.n11582 0.000507003
R18702 VSS.n11629 VSS.n11583 0.000507003
R18703 VSS.n11624 VSS.n11623 0.000507003
R18704 VSS.n12384 VSS.n12383 0.000507003
R18705 VSS.n12453 VSS.n12384 0.000507003
R18706 VSS.n12378 VSS.n12377 0.000507003
R18707 VSS.n12368 VSS.n12367 0.000507003
R18708 VSS.n12456 VSS.n12455 0.000507003
R18709 VSS.n2977 VSS.n2943 0.000507003
R18710 VSS.n2996 VSS.n2980 0.000507003
R18711 VSS.n2992 VSS.n2981 0.000507003
R18712 VSS.n2989 VSS.n2983 0.000507003
R18713 VSS.n12743 VSS.n12742 0.000507003
R18714 VSS.n12748 VSS.n12747 0.000507003
R18715 VSS.n12753 VSS.n12752 0.000507003
R18716 VSS.n12756 VSS.n2944 0.000507003
R18717 VSS.n12772 VSS.n2940 0.000507003
R18718 VSS.n12796 VSS.n2940 0.000507003
R18719 VSS.n12769 VSS.n12768 0.000507003
R18720 VSS.n12777 VSS.n12776 0.000507003
R18721 VSS.n12780 VSS.n12779 0.000507003
R18722 VSS.n13968 VSS.n1759 0.000507003
R18723 VSS.n13987 VSS.n13971 0.000507003
R18724 VSS.n13983 VSS.n13972 0.000507003
R18725 VSS.n13980 VSS.n13974 0.000507003
R18726 VSS.n13952 VSS.n13951 0.000507003
R18727 VSS.n13956 VSS.n13955 0.000507003
R18728 VSS.n13961 VSS.n13960 0.000507003
R18729 VSS.n13964 VSS.n13963 0.000507003
R18730 VSS.n1734 VSS.n1733 0.000507003
R18731 VSS.n14016 VSS.n1734 0.000507003
R18732 VSS.n1731 VSS.n1730 0.000507003
R18733 VSS.n14020 VSS.n1718 0.000507003
R18734 VSS.n1719 VSS.n1716 0.000507003
R18735 VSS.n13555 VSS.n13510 0.000507003
R18736 VSS.n13552 VSS.n13513 0.000507003
R18737 VSS.n13528 VSS.n13518 0.000507003
R18738 VSS.n13524 VSS.n13519 0.000507003
R18739 VSS.n13569 VSS.n13568 0.000507003
R18740 VSS.n13572 VSS.n13561 0.000507003
R18741 VSS.n13576 VSS.n13575 0.000507003
R18742 VSS.n13579 VSS.n13511 0.000507003
R18743 VSS.n13499 VSS.n13498 0.000507003
R18744 VSS.n13603 VSS.n13499 0.000507003
R18745 VSS.n13496 VSS.n13495 0.000507003
R18746 VSS.n13607 VSS.n13483 0.000507003
R18747 VSS.n13484 VSS.n13481 0.000507003
R18748 VSS.n13300 VSS.n13299 0.000507003
R18749 VSS.n13305 VSS.n13304 0.000507003
R18750 VSS.n13311 VSS.n13310 0.000507003
R18751 VSS.n13317 VSS.n13316 0.000507003
R18752 VSS.n13333 VSS.n13332 0.000507003
R18753 VSS.n13339 VSS.n13338 0.000507003
R18754 VSS.n13347 VSS.n13346 0.000507003
R18755 VSS.n13342 VSS.n13341 0.000507003
R18756 VSS.n13449 VSS.n13448 0.000507003
R18757 VSS.n13473 VSS.n13449 0.000507003
R18758 VSS.n13443 VSS.n13442 0.000507003
R18759 VSS.n13433 VSS.n13432 0.000507003
R18760 VSS.n13406 VSS.n13405 0.000507003
R18761 VSS.n11499 VSS.n11498 0.000506803
R18762 VSS.n11500 VSS.n11499 0.000506803
R18763 VSS.n11339 VSS.n11338 0.000505632
R18764 VSS.n11342 VSS.n11341 0.000505632
R18765 VSS.n11197 VSS.n11196 0.000505632
R18766 VSS.n11327 VSS.n11326 0.000505632
R18767 VSS.n11505 VSS.n11504 0.000505632
R18768 VSS.n11510 VSS.n11509 0.000505632
R18769 VSS.n10800 VSS.n10799 0.000505597
R18770 VSS.n10793 VSS.n10792 0.000505597
R18771 VSS.n10645 VSS.n10644 0.000505597
R18772 VSS.n4456 VSS.n4455 0.000505597
R18773 VSS.n10741 VSS.n10740 0.000505597
R18774 VSS.n4103 VSS.n4102 0.000505597
R18775 VSS.n10797 VSS.n10796 0.000505597
R18776 VSS.n10789 VSS.n10788 0.000505597
R18777 VSS.n10642 VSS.n10641 0.000505597
R18778 VSS.n10738 VSS.n10737 0.000505597
R18779 VSS.n10608 VSS.n10607 0.000505094
R18780 VSS.n3373 VSS.n3372 0.000505094
R18781 VSS.n5394 VSS.n5393 0.000505094
R18782 VSS.n5396 VSS.n5394 0.000505094
R18783 VSS.n5396 VSS.n5395 0.000505094
R18784 VSS.n6133 VSS.n6132 0.000505094
R18785 VSS.n6135 VSS.n6133 0.000505094
R18786 VSS.n6117 VSS.n6116 0.000505094
R18787 VSS.n6119 VSS.n6117 0.000505094
R18788 VSS.n6119 VSS.n6118 0.000505094
R18789 VSS.n5951 VSS.n5950 0.000505094
R18790 VSS.n5953 VSS.n5951 0.000505094
R18791 VSS.n5953 VSS.n5952 0.000505094
R18792 VSS.n5935 VSS.n5934 0.000505094
R18793 VSS.n5937 VSS.n5935 0.000505094
R18794 VSS.n5937 VSS.n5936 0.000505094
R18795 VSS.n5770 VSS.n5769 0.000505094
R18796 VSS.n5772 VSS.n5770 0.000505094
R18797 VSS.n5772 VSS.n5771 0.000505094
R18798 VSS.n5754 VSS.n5753 0.000505094
R18799 VSS.n5756 VSS.n5754 0.000505094
R18800 VSS.n5756 VSS.n5755 0.000505094
R18801 VSS.n5590 VSS.n5589 0.000505094
R18802 VSS.n5592 VSS.n5590 0.000505094
R18803 VSS.n5592 VSS.n5591 0.000505094
R18804 VSS.n5574 VSS.n5573 0.000505094
R18805 VSS.n5576 VSS.n5574 0.000505094
R18806 VSS.n5576 VSS.n5575 0.000505094
R18807 VSS.n5410 VSS.n5409 0.000505094
R18808 VSS.n5412 VSS.n5410 0.000505094
R18809 VSS.n5412 VSS.n5411 0.000505094
R18810 VSS.n5230 VSS.n5229 0.000505094
R18811 VSS.n5232 VSS.n5230 0.000505094
R18812 VSS.n5232 VSS.n5231 0.000505094
R18813 VSS.n5214 VSS.n5213 0.000505094
R18814 VSS.n5216 VSS.n5214 0.000505094
R18815 VSS.n5216 VSS.n5215 0.000505094
R18816 VSS.n10117 VSS.n10116 0.000505094
R18817 VSS.n10117 VSS.n10111 0.000505094
R18818 VSS.n10111 VSS.n10110 0.000505094
R18819 VSS.n10162 VSS.n10161 0.000505094
R18820 VSS.n10162 VSS.n10127 0.000505094
R18821 VSS.n10127 VSS.n10126 0.000505094
R18822 VSS.n11160 VSS.n11159 0.000505094
R18823 VSS.n11160 VSS.n11154 0.000505094
R18824 VSS.n11154 VSS.n11153 0.000505094
R18825 VSS.n11176 VSS.n11175 0.000505094
R18826 VSS.n11176 VSS.n11170 0.000505094
R18827 VSS.n11170 VSS.n11169 0.000505094
R18828 VSS.n12296 VSS.n12290 0.000505094
R18829 VSS.n12296 VSS.n12295 0.000505094
R18830 VSS.n12319 VSS.n12318 0.000505094
R18831 VSS.n12323 VSS.n12319 0.000505094
R18832 VSS.n11560 VSS.n11559 0.000505094
R18833 VSS.n12475 VSS.n12474 0.000505094
R18834 VSS.n12476 VSS.n3612 0.000505094
R18835 VSS.n12476 VSS.n12475 0.000505094
R18836 VSS.n12176 VSS.n12175 0.000505094
R18837 VSS.n12180 VSS.n12176 0.000505094
R18838 VSS.n12194 VSS.n12193 0.000505094
R18839 VSS.n12198 VSS.n12194 0.000505094
R18840 VSS.n14494 VSS.n14488 0.000505094
R18841 VSS.n14485 VSS.n14482 0.000505094
R18842 VSS.n14485 VSS.n14484 0.000505094
R18843 VSS.n3318 VSS.n3317 0.000505094
R18844 VSS.n12567 VSS.n12559 0.000505094
R18845 VSS.n3410 VSS.n3409 0.000505094
R18846 VSS.n3414 VSS.n3410 0.000505094
R18847 VSS.n3585 VSS.n3579 0.000505094
R18848 VSS.n3585 VSS.n3584 0.000505094
R18849 VSS.n11895 VSS.n11894 0.000505094
R18850 VSS.n11899 VSS.n11895 0.000505094
R18851 VSS.n12009 VSS.n12008 0.000505094
R18852 VSS.n12012 VSS.n12009 0.000505094
R18853 VSS.n12026 VSS.n12025 0.000505094
R18854 VSS.n12028 VSS.n12026 0.000505094
R18855 VSS.n10621 VSS.n10617 0.000505094
R18856 VSS.n11528 VSS.n11527 0.00050467
R18857 VSS.n1508 VSS.n1507 0.00050467
R18858 VSS.n6148 VSS.n6147 0.00050467
R18859 VSS.n9740 VSS.n9739 0.00050467
R18860 VSS.n8423 VSS.n8422 0.00050467
R18861 VSS.n8337 VSS.n8336 0.00050467
R18862 VSS.n8648 VSS.n8647 0.00050467
R18863 VSS.n7514 VSS.n7513 0.00050467
R18864 VSS.n9723 VSS.n9722 0.00050467
R18865 VSS.n7488 VSS.n7487 0.00050467
R18866 VSS.n3965 VSS.n3964 0.00050467
R18867 VSS.n6096 VSS.n6095 0.00050467
R18868 VSS.n5965 VSS.n5964 0.00050467
R18869 VSS.n5914 VSS.n5913 0.00050467
R18870 VSS.n5784 VSS.n5783 0.00050467
R18871 VSS.n5733 VSS.n5732 0.00050467
R18872 VSS.n5603 VSS.n5602 0.00050467
R18873 VSS.n5553 VSS.n5552 0.00050467
R18874 VSS.n5423 VSS.n5422 0.00050467
R18875 VSS.n5373 VSS.n5372 0.00050467
R18876 VSS.n5243 VSS.n5242 0.00050467
R18877 VSS.n5193 VSS.n5192 0.00050467
R18878 VSS.n10103 VSS.n10102 0.00050467
R18879 VSS.n10141 VSS.n10140 0.00050467
R18880 VSS.n3702 VSS.n3701 0.00050467
R18881 VSS.n11146 VSS.n11145 0.00050467
R18882 VSS.n11521 VSS.n11520 0.00050467
R18883 VSS.n10732 VSS.n10731 0.00050467
R18884 VSS.n10722 VSS.n10721 0.00050467
R18885 VSS.n987 VSS.n986 0.00050467
R18886 VSS.n14373 VSS.n14372 0.00050467
R18887 VSS.n10719 VSS.n10717 0.00050467
R18888 VSS.n504 VSS.n503 0.00050467
R18889 VSS.n10648 VSS.n10647 0.00050467
R18890 VSS.n8427 VSS.n8426 0.00050467
R18891 VSS.n8335 VSS.n8334 0.00050467
R18892 VSS.n8637 VSS.n8636 0.00050467
R18893 VSS.n8328 VSS.n8327 0.00050467
R18894 VSS.n8725 VSS.n8724 0.00050467
R18895 VSS.n7512 VSS.n7511 0.00050467
R18896 VSS.n9712 VSS.n9711 0.00050467
R18897 VSS.n7505 VSS.n7504 0.00050467
R18898 VSS.n9729 VSS.n9728 0.00050467
R18899 VSS.n9745 VSS.n9744 0.00050467
R18900 VSS.n9357 VSS.n7493 0.00050467
R18901 VSS.n7485 VSS.n7484 0.00050467
R18902 VSS.n3963 VSS.n3962 0.00050467
R18903 VSS.n10814 VSS.n10813 0.00050467
R18904 VSS.n10807 VSS.n10806 0.00050467
R18905 VSS.n4031 VSS.n4030 0.00050467
R18906 VSS.n9764 VSS.n9763 0.00050467
R18907 VSS.n9767 VSS.n9766 0.00050467
R18908 VSS.n9752 VSS.n9751 0.00050467
R18909 VSS.n9421 VSS.n7491 0.00050467
R18910 VSS.n9736 VSS.n9735 0.00050467
R18911 VSS.n9056 VSS.n7495 0.00050467
R18912 VSS.n9719 VSS.n9718 0.00050467
R18913 VSS.n9698 VSS.n7507 0.00050467
R18914 VSS.n8718 VSS.n8717 0.00050467
R18915 VSS.n8714 VSS.n8713 0.00050467
R18916 VSS.n8644 VSS.n8643 0.00050467
R18917 VSS.n8623 VSS.n8330 0.00050467
R18918 VSS.n4097 VSS.n4096 0.00050467
R18919 VSS.n4093 VSS.n4092 0.00050467
R18920 VSS.n991 VSS.n990 0.00050467
R18921 VSS.n14352 VSS.n14351 0.00050467
R18922 VSS.n14357 VSS.n14356 0.00050467
R18923 VSS.n1242 VSS.n1241 0.00050467
R18924 VSS.n1071 VSS.n1070 0.00050467
R18925 VSS.n1067 VSS.n1066 0.00050467
R18926 VSS.n1233 VSS.n1232 0.00050467
R18927 VSS.n704 VSS.n703 0.00050467
R18928 VSS.n13746 VSS.n13745 0.00050467
R18929 VSS.n13753 VSS.n13752 0.00050467
R18930 VSS.n13283 VSS.n13282 0.00050467
R18931 VSS.n13291 VSS.n13290 0.00050467
R18932 VSS.n13829 VSS.n13828 0.00050467
R18933 VSS.n13833 VSS.n13832 0.00050467
R18934 VSS.n1589 VSS.n1588 0.00050467
R18935 VSS.n1593 VSS.n1592 0.00050467
R18936 VSS.n12354 VSS.n12353 0.00050467
R18937 VSS.n12330 VSS.n12329 0.00050467
R18938 VSS.n12271 VSS.n12270 0.00050467
R18939 VSS.n12204 VSS.n12203 0.00050467
R18940 VSS.n11804 VSS.n11803 0.00050467
R18941 VSS.n12040 VSS.n12039 0.00050467
R18942 VSS.n11821 VSS.n11820 0.00050467
R18943 VSS.n11927 VSS.n11926 0.00050467
R18944 VSS.n3392 VSS.n3391 0.00050467
R18945 VSS.n3442 VSS.n3441 0.00050467
R18946 VSS.n3338 VSS.n3337 0.00050467
R18947 VSS.n12577 VSS.n12576 0.00050467
R18948 VSS.n3296 VSS.n3295 0.00050467
R18949 VSS.n13413 VSS.n13412 0.00050467
R18950 VSS.n13423 VSS.n13422 0.00050467
R18951 VSS.n13352 VSS.n13351 0.00050467
R18952 VSS.n13368 VSS.n13367 0.00050467
R18953 VSS.n1512 VSS.n1511 0.00050467
R18954 VSS.n460 VSS.n459 0.00050467
R18955 VSS.n466 VSS.n465 0.00050467
R18956 VSS.n695 VSS.n694 0.00050467
R18957 VSS.n689 VSS.n688 0.00050467
R18958 VSS.n1318 VSS.n1317 0.00050467
R18959 VSS.n1321 VSS.n1320 0.00050467
R18960 VSS.n3303 VSS.n3302 0.00050467
R18961 VSS.n3360 VSS.n3359 0.00050467
R18962 VSS.n3335 VSS.n3334 0.00050467
R18963 VSS.n3567 VSS.n3566 0.00050467
R18964 VSS.n3389 VSS.n3388 0.00050467
R18965 VSS.n11996 VSS.n11995 0.00050467
R18966 VSS.n11818 VSS.n11817 0.00050467
R18967 VSS.n12163 VSS.n12162 0.00050467
R18968 VSS.n11801 VSS.n11800 0.00050467
R18969 VSS.n12278 VSS.n12277 0.00050467
R18970 VSS.n12350 VSS.n12349 0.00050467
R18971 VSS.n12358 VSS.n12357 0.00050467
R18972 VSS.n12337 VSS.n12336 0.00050467
R18973 VSS.n11756 VSS.n11755 0.00050467
R18974 VSS.n12036 VSS.n12035 0.00050467
R18975 VSS.n11919 VSS.n11918 0.00050467
R18976 VSS.n3438 VSS.n3437 0.00050467
R18977 VSS.n12573 VSS.n12572 0.00050467
R18978 VSS.n12466 VSS.n12465 0.00050467
R18979 VSS.n11518 VSS.n11517 0.00050467
R18980 VSS.n3711 VSS.n3710 0.00050467
R18981 VSS.n6145 VSS.n6144 0.00050467
R18982 VSS.n10138 VSS.n10137 0.00050467
R18983 VSS.n10149 VSS.n10148 0.00050467
R18984 VSS.n5190 VSS.n5189 0.00050467
R18985 VSS.n5201 VSS.n5200 0.00050467
R18986 VSS.n5370 VSS.n5369 0.00050467
R18987 VSS.n5381 VSS.n5380 0.00050467
R18988 VSS.n5550 VSS.n5549 0.00050467
R18989 VSS.n5561 VSS.n5560 0.00050467
R18990 VSS.n5730 VSS.n5729 0.00050467
R18991 VSS.n5741 VSS.n5740 0.00050467
R18992 VSS.n5911 VSS.n5910 0.00050467
R18993 VSS.n5922 VSS.n5921 0.00050467
R18994 VSS.n6093 VSS.n6092 0.00050467
R18995 VSS.n6104 VSS.n6103 0.00050467
R18996 VSS.n5962 VSS.n5961 0.00050467
R18997 VSS.n5781 VSS.n5780 0.00050467
R18998 VSS.n5600 VSS.n5599 0.00050467
R18999 VSS.n5420 VSS.n5419 0.00050467
R19000 VSS.n5240 VSS.n5239 0.00050467
R19001 VSS.n4569 VSS.n4568 0.00050467
R19002 VSS.n11077 VSS.n11076 0.00050467
R19003 VSS.n11191 VSS.n11190 0.00050467
R19004 VSS.n9357 VSS.n9356 0.000504623
R19005 VSS.n9358 VSS.n9357 0.000504623
R19006 VSS.n8636 VSS.n8341 0.000504623
R19007 VSS.n8636 VSS.n8635 0.000504623
R19008 VSS.n8725 VSS.n8323 0.000504623
R19009 VSS.n8726 VSS.n8725 0.000504623
R19010 VSS.n9711 VSS.n7518 0.000504623
R19011 VSS.n9711 VSS.n9710 0.000504623
R19012 VSS.n9728 VSS.n9727 0.000504623
R19013 VSS.n10814 VSS.n3958 0.000504623
R19014 VSS.n10815 VSS.n10814 0.000504623
R19015 VSS.n6092 VSS.n6091 0.000504623
R19016 VSS.n5910 VSS.n5909 0.000504623
R19017 VSS.n5729 VSS.n5728 0.000504623
R19018 VSS.n5549 VSS.n5548 0.000504623
R19019 VSS.n5369 VSS.n5368 0.000504623
R19020 VSS.n5189 VSS.n5188 0.000504623
R19021 VSS.n10137 VSS.n10136 0.000504623
R19022 VSS.n11078 VSS.n11077 0.000504623
R19023 VSS.n11190 VSS.n11189 0.000504623
R19024 VSS.n12349 VSS.n12348 0.000504623
R19025 VSS.n12268 VSS.n11690 0.000504623
R19026 VSS.n12270 VSS.n12268 0.000504623
R19027 VSS.n12162 VSS.n12161 0.000504623
R19028 VSS.n11995 VSS.n11994 0.000504623
R19029 VSS.n3566 VSS.n3565 0.000504623
R19030 VSS.n3359 VSS.n3358 0.000504623
R19031 VSS.n3293 VSS.n3185 0.000504623
R19032 VSS.n3295 VSS.n3293 0.000504623
R19033 VSS.n10 VSS.n9 0.000504623
R19034 VSS.n14507 VSS.n10 0.000504623
R19035 VSS.n11343 VSS.n11342 0.000504168
R19036 VSS.n11504 VSS.n11503 0.000504168
R19037 VSS.n11326 VSS.n11325 0.000504168
R19038 VSS.n10799 VSS.n10798 0.000504146
R19039 VSS.n4102 VSS.n4101 0.000504146
R19040 VSS.n10796 VSS.n10795 0.000504146
R19041 VSS.n10788 VSS.n10787 0.000504146
R19042 VSS.n10644 VSS.n10643 0.000504146
R19043 VSS.n10742 VSS.n10741 0.000504146
R19044 VSS.n4455 VSS.n4454 0.000504146
R19045 VSS.n10641 VSS.n10640 0.000504146
R19046 VSS.n9024 VSS.n9023 0.000503845
R19047 VSS.n7525 VSS.n7524 0.000503845
R19048 VSS.n8780 VSS.n8243 0.000503845
R19049 VSS.n6742 VSS.n6741 0.000503845
R19050 VSS.n8117 VSS.n8116 0.000503845
R19051 VSS.n8874 VSS.n8873 0.000503845
R19052 VSS.n8818 VSS.n8817 0.000503845
R19053 VSS.n9556 VSS.n9555 0.000503845
R19054 VSS.n8461 VSS.n8460 0.000503845
R19055 VSS.n7425 VSS.n7424 0.000503845
R19056 VSS.n9062 VSS.n9061 0.000503845
R19057 VSS.n9513 VSS.n9512 0.000503845
R19058 VSS.n9835 VSS.n9834 0.000503845
R19059 VSS.n7370 VSS.n7369 0.000503845
R19060 VSS.n9242 VSS.n9241 0.000503845
R19061 VSS.n8949 VSS.n8948 0.000503845
R19062 VSS.n7639 VSS.n7632 0.000503845
R19063 VSS.n7674 VSS.n7667 0.000503845
R19064 VSS.n7140 VSS.n7139 0.000503845
R19065 VSS.n8924 VSS.n8923 0.000503845
R19066 VSS.n6857 VSS.n6856 0.000503845
R19067 VSS.n6924 VSS.n6923 0.000503845
R19068 VSS.n6997 VSS.n6996 0.000503845
R19069 VSS.n7056 VSS.n7055 0.000503845
R19070 VSS.n6424 VSS.n6423 0.000503845
R19071 VSS.n6789 VSS.n6788 0.000503845
R19072 VSS.n5797 VSS.n5796 0.000503845
R19073 VSS.n5616 VSS.n5615 0.000503845
R19074 VSS.n5256 VSS.n5255 0.000503845
R19075 VSS.n3758 VSS.n3757 0.000503845
R19076 VSS.n6079 VSS.n6078 0.000503845
R19077 VSS.n6182 VSS.n6181 0.000503845
R19078 VSS.n11072 VSS.n11071 0.000503845
R19079 VSS.n11029 VSS.n11028 0.000503845
R19080 VSS.n10944 VSS.n10917 0.000503845
R19081 VSS.n10878 VSS.n10877 0.000503845
R19082 VSS.n4055 VSS.n4054 0.000503845
R19083 VSS.n4269 VSS.n4268 0.000503845
R19084 VSS.n4381 VSS.n4380 0.000503845
R19085 VSS.n4450 VSS.n4133 0.000503845
R19086 VSS.n513 VSS.n512 0.000503845
R19087 VSS.n1132 VSS.n1131 0.000503845
R19088 VSS.n13048 VSS.n13047 0.000503845
R19089 VSS.n13095 VSS.n13094 0.000503845
R19090 VSS.n2345 VSS.n2344 0.000503845
R19091 VSS.n2401 VSS.n2400 0.000503845
R19092 VSS.n1168 VSS.n1167 0.000503845
R19093 VSS.n1522 VSS.n1521 0.000503845
R19094 VSS.n13762 VSS.n13761 0.000503845
R19095 VSS.n14112 VSS.n14111 0.000503845
R19096 VSS.n1669 VSS.n1662 0.000503845
R19097 VSS.n13646 VSS.n13645 0.000503845
R19098 VSS.n1412 VSS.n1411 0.000503845
R19099 VSS.n2242 VSS.n2241 0.000503845
R19100 VSS.n2177 VSS.n2176 0.000503845
R19101 VSS.n13191 VSS.n13190 0.000503845
R19102 VSS.n13929 VSS.n13928 0.000503845
R19103 VSS.n1976 VSS.n1973 0.000503845
R19104 VSS.n12982 VSS.n12981 0.000503845
R19105 VSS.n2696 VSS.n2689 0.000503845
R19106 VSS.n12905 VSS.n12904 0.000503845
R19107 VSS.n2876 VSS.n2869 0.000503845
R19108 VSS.n12724 VSS.n12723 0.000503845
R19109 VSS.n2528 VSS.n2525 0.000503845
R19110 VSS.n11575 VSS.n11574 0.000503845
R19111 VSS.n11698 VSS.n11697 0.000503845
R19112 VSS.n12051 VSS.n12050 0.000503845
R19113 VSS.n11830 VSS.n11829 0.000503845
R19114 VSS.n3455 VSS.n3454 0.000503845
R19115 VSS.n12387 VSS.n12386 0.000503845
R19116 VSS.n11629 VSS.n11628 0.000503845
R19117 VSS.n12783 VSS.n12782 0.000503845
R19118 VSS.n1766 VSS.n1765 0.000503845
R19119 VSS.n13585 VSS.n13584 0.000503845
R19120 VSS.n13452 VSS.n13451 0.000503845
R19121 VSS.n10614 VSS.n10613 0.000503113
R19122 VSS.n10610 VSS.n10609 0.000503113
R19123 VSS.n4539 VSS.n4538 0.000503113
R19124 VSS.n6125 VSS.n6124 0.000503113
R19125 VSS.n6121 VSS.n6120 0.000503113
R19126 VSS.n6109 VSS.n6108 0.000503113
R19127 VSS.n5955 VSS.n5954 0.000503113
R19128 VSS.n5943 VSS.n5942 0.000503113
R19129 VSS.n5939 VSS.n5938 0.000503113
R19130 VSS.n5927 VSS.n5926 0.000503113
R19131 VSS.n5774 VSS.n5773 0.000503113
R19132 VSS.n5762 VSS.n5761 0.000503113
R19133 VSS.n5758 VSS.n5757 0.000503113
R19134 VSS.n5746 VSS.n5745 0.000503113
R19135 VSS.n5594 VSS.n5593 0.000503113
R19136 VSS.n5582 VSS.n5581 0.000503113
R19137 VSS.n5578 VSS.n5577 0.000503113
R19138 VSS.n5566 VSS.n5565 0.000503113
R19139 VSS.n5414 VSS.n5413 0.000503113
R19140 VSS.n5402 VSS.n5401 0.000503113
R19141 VSS.n5398 VSS.n5397 0.000503113
R19142 VSS.n5386 VSS.n5385 0.000503113
R19143 VSS.n5234 VSS.n5233 0.000503113
R19144 VSS.n5222 VSS.n5221 0.000503113
R19145 VSS.n5218 VSS.n5217 0.000503113
R19146 VSS.n5206 VSS.n5205 0.000503113
R19147 VSS.n10109 VSS.n10108 0.000503113
R19148 VSS.n10121 VSS.n10120 0.000503113
R19149 VSS.n10125 VSS.n10124 0.000503113
R19150 VSS.n10154 VSS.n10153 0.000503113
R19151 VSS.n11152 VSS.n11151 0.000503113
R19152 VSS.n11164 VSS.n11163 0.000503113
R19153 VSS.n11168 VSS.n11167 0.000503113
R19154 VSS.n11180 VSS.n11179 0.000503113
R19155 VSS.n12473 VSS.n12472 0.000503113
R19156 VSS.n11564 VSS.n11563 0.000503113
R19157 VSS.n11557 VSS.n11556 0.000503113
R19158 VSS.n3310 VSS.n3309 0.000503113
R19159 VSS.n3315 VSS.n3314 0.000503113
R19160 VSS.n12556 VSS.n12555 0.000503113
R19161 VSS.n12569 VSS.n12568 0.000503113
R19162 VSS.n3365 VSS.n3364 0.000503113
R19163 VSS.n3370 VSS.n3369 0.000503113
R19164 VSS.n3402 VSS.n3401 0.000503113
R19165 VSS.n3416 VSS.n3415 0.000503113
R19166 VSS.n3572 VSS.n3571 0.000503113
R19167 VSS.n3582 VSS.n3581 0.000503113
R19168 VSS.n11887 VSS.n11886 0.000503113
R19169 VSS.n11901 VSS.n11900 0.000503113
R19170 VSS.n12001 VSS.n12000 0.000503113
R19171 VSS.n12014 VSS.n12013 0.000503113
R19172 VSS.n12018 VSS.n12017 0.000503113
R19173 VSS.n12030 VSS.n12029 0.000503113
R19174 VSS.n12168 VSS.n12167 0.000503113
R19175 VSS.n12182 VSS.n12181 0.000503113
R19176 VSS.n12186 VSS.n12185 0.000503113
R19177 VSS.n12200 VSS.n12199 0.000503113
R19178 VSS.n12283 VSS.n12282 0.000503113
R19179 VSS.n12293 VSS.n12292 0.000503113
R19180 VSS.n12311 VSS.n12310 0.000503113
R19181 VSS.n12325 VSS.n12324 0.000503113
R19182 VSS.n12470 VSS.n12469 0.000503113
R19183 VSS.n6137 VSS.n6136 0.000503113
R19184 VSS.n10637 VSS.n10636 0.000503113
R19185 VSS.n12024 VSS.n12023 0.000503113
R19186 VSS.n12007 VSS.n12006 0.000503113
R19187 VSS.n11893 VSS.n11892 0.000503113
R19188 VSS.n3578 VSS.n3577 0.000503113
R19189 VSS.n3408 VSS.n3407 0.000503113
R19190 VSS.n3325 VSS.n3324 0.000503113
R19191 VSS.n12563 VSS.n12562 0.000503113
R19192 VSS.n3180 VSS.n3179 0.000503113
R19193 VSS.n12192 VSS.n12191 0.000503113
R19194 VSS.n12174 VSS.n12173 0.000503113
R19195 VSS.n11174 VSS.n11173 0.000503113
R19196 VSS.n11158 VSS.n11157 0.000503113
R19197 VSS.n10160 VSS.n10159 0.000503113
R19198 VSS.n10115 VSS.n10114 0.000503113
R19199 VSS.n5212 VSS.n5211 0.000503113
R19200 VSS.n5228 VSS.n5227 0.000503113
R19201 VSS.n5392 VSS.n5391 0.000503113
R19202 VSS.n5408 VSS.n5407 0.000503113
R19203 VSS.n5572 VSS.n5571 0.000503113
R19204 VSS.n5588 VSS.n5587 0.000503113
R19205 VSS.n5752 VSS.n5751 0.000503113
R19206 VSS.n5768 VSS.n5767 0.000503113
R19207 VSS.n5933 VSS.n5932 0.000503113
R19208 VSS.n5949 VSS.n5948 0.000503113
R19209 VSS.n6115 VSS.n6114 0.000503113
R19210 VSS.n6131 VSS.n6130 0.000503113
R19211 VSS.n3609 VSS.n3608 0.000503113
R19212 VSS.n12317 VSS.n12316 0.000503113
R19213 VSS.n12289 VSS.n12288 0.000503113
R19214 VSS.n11551 VSS.n11550 0.000503113
R19215 VSS.n10620 VSS.n10619 0.000503113
R19216 VSS.n10625 VSS.n10624 0.000503113
R19217 VSS.n13462 VSS.n13461 0.000502702
R19218 VSS.n13597 VSS.n13596 0.000502702
R19219 VSS.n14010 VSS.n14009 0.000502702
R19220 VSS.n12792 VSS.n12791 0.000502702
R19221 VSS.n3111 VSS.n3110 0.000502702
R19222 VSS.n3536 VSS.n3535 0.000502702
R19223 VSS.n11964 VSS.n11963 0.000502702
R19224 VSS.n12132 VSS.n12131 0.000502702
R19225 VSS.n2892 VSS.n2879 0.000502702
R19226 VSS.n2804 VSS.n2803 0.000502702
R19227 VSS.n4072 VSS.n4071 0.000502702
R19228 VSS.n10887 VSS.n10886 0.000502702
R19229 VSS.n10932 VSS.n10931 0.000502702
R19230 VSS.n11038 VSS.n11037 0.000502702
R19231 VSS.n10071 VSS.n10070 0.000502702
R19232 VSS.n5337 VSS.n5336 0.000502702
R19233 VSS.n5517 VSS.n5516 0.000502702
R19234 VSS.n5697 VSS.n5696 0.000502702
R19235 VSS.n6575 VSS.n6560 0.000502702
R19236 VSS.n9648 VSS.n9647 0.000502702
R19237 VSS.n9685 VSS.n9684 0.000502702
R19238 VSS.n8486 VSS.n8485 0.000502702
R19239 VSS.n8660 VSS.n8659 0.000502702
R19240 VSS.n8697 VSS.n8696 0.000502702
R19241 VSS.n8595 VSS.n8594 0.000502702
R19242 VSS.n8601 VSS.n8600 0.000502702
R19243 VSS.n8608 VSS.n8607 0.000502702
R19244 VSS.n8793 VSS.n8792 0.000502702
R19245 VSS.n6195 VSS.n6194 0.000502702
R19246 VSS.n6207 VSS.n6206 0.000502702
R19247 VSS.n9962 VSS.n9961 0.000502702
R19248 VSS.n9971 VSS.n9970 0.000502702
R19249 VSS.n8146 VSS.n8145 0.000502702
R19250 VSS.n8856 VSS.n8855 0.000502702
R19251 VSS.n8864 VSS.n8004 0.000502702
R19252 VSS.n8831 VSS.n8830 0.000502702
R19253 VSS.n7577 VSS.n7574 0.000502702
R19254 VSS.n7587 VSS.n7586 0.000502702
R19255 VSS.n9550 VSS.n9549 0.000502702
R19256 VSS.n8451 VSS.n8450 0.000502702
R19257 VSS.n8436 VSS.n8435 0.000502702
R19258 VSS.n9395 VSS.n9394 0.000502702
R19259 VSS.n9408 VSS.n9407 0.000502702
R19260 VSS.n7452 VSS.n7451 0.000502702
R19261 VSS.n7458 VSS.n7457 0.000502702
R19262 VSS.n7465 VSS.n7464 0.000502702
R19263 VSS.n9089 VSS.n9088 0.000502702
R19264 VSS.n9095 VSS.n9094 0.000502702
R19265 VSS.n9102 VSS.n9101 0.000502702
R19266 VSS.n9011 VSS.n9010 0.000502702
R19267 VSS.n9521 VSS.n9520 0.000502702
R19268 VSS.n9843 VSS.n9842 0.000502702
R19269 VSS.n7161 VSS.n7157 0.000502702
R19270 VSS.n7175 VSS.n7174 0.000502702
R19271 VSS.n9481 VSS.n9468 0.000502702
R19272 VSS.n9485 VSS.n9484 0.000502702
R19273 VSS.n9473 VSS.n9469 0.000502702
R19274 VSS.n9830 VSS.n9829 0.000502702
R19275 VSS.n7315 VSS.n7312 0.000502702
R19276 VSS.n7323 VSS.n7313 0.000502702
R19277 VSS.n7205 VSS.n7189 0.000502702
R19278 VSS.n7203 VSS.n7202 0.000502702
R19279 VSS.n9221 VSS.n9218 0.000502702
R19280 VSS.n9231 VSS.n9230 0.000502702
R19281 VSS.n9236 VSS.n9235 0.000502702
R19282 VSS.n8943 VSS.n8942 0.000502702
R19283 VSS.n7860 VSS.n7857 0.000502702
R19284 VSS.n7907 VSS.n7894 0.000502702
R19285 VSS.n7917 VSS.n7916 0.000502702
R19286 VSS.n7902 VSS.n7895 0.000502702
R19287 VSS.n8953 VSS.n7844 0.000502702
R19288 VSS.n8982 VSS.n8981 0.000502702
R19289 VSS.n8978 VSS.n8977 0.000502702
R19290 VSS.n8976 VSS.n8975 0.000502702
R19291 VSS.n7614 VSS.n7610 0.000502702
R19292 VSS.n8990 VSS.n8989 0.000502702
R19293 VSS.n7623 VSS.n7611 0.000502702
R19294 VSS.n7803 VSS.n7802 0.000502702
R19295 VSS.n7772 VSS.n7771 0.000502702
R19296 VSS.n7768 VSS.n7767 0.000502702
R19297 VSS.n7766 VSS.n7765 0.000502702
R19298 VSS.n7658 VSS.n7646 0.000502702
R19299 VSS.n7780 VSS.n7779 0.000502702
R19300 VSS.n7649 VSS.n7645 0.000502702
R19301 VSS.n7724 VSS.n7723 0.000502702
R19302 VSS.n7113 VSS.n7112 0.000502702
R19303 VSS.n7106 VSS.n7105 0.000502702
R19304 VSS.n9877 VSS.n9876 0.000502702
R19305 VSS.n9879 VSS.n9878 0.000502702
R19306 VSS.n7987 VSS.n7986 0.000502702
R19307 VSS.n7998 VSS.n7997 0.000502702
R19308 VSS.n6623 VSS.n6608 0.000502702
R19309 VSS.n6851 VSS.n6850 0.000502702
R19310 VSS.n6651 VSS.n6645 0.000502702
R19311 VSS.n6807 VSS.n6794 0.000502702
R19312 VSS.n6811 VSS.n6810 0.000502702
R19313 VSS.n6799 VSS.n6795 0.000502702
R19314 VSS.n6892 VSS.n6891 0.000502702
R19315 VSS.n6902 VSS.n6901 0.000502702
R19316 VSS.n6918 VSS.n6917 0.000502702
R19317 VSS.n6607 VSS.n6606 0.000502702
R19318 VSS.n6603 VSS.n6597 0.000502702
R19319 VSS.n6875 VSS.n6862 0.000502702
R19320 VSS.n6879 VSS.n6878 0.000502702
R19321 VSS.n6867 VSS.n6863 0.000502702
R19322 VSS.n6965 VSS.n6964 0.000502702
R19323 VSS.n6975 VSS.n6974 0.000502702
R19324 VSS.n6991 VSS.n6990 0.000502702
R19325 VSS.n6559 VSS.n6558 0.000502702
R19326 VSS.n6549 VSS.n6546 0.000502702
R19327 VSS.n6937 VSS.n6930 0.000502702
R19328 VSS.n6952 VSS.n6951 0.000502702
R19329 VSS.n6942 VSS.n6929 0.000502702
R19330 VSS.n7035 VSS.n6533 0.000502702
R19331 VSS.n7050 VSS.n7049 0.000502702
R19332 VSS.n6509 VSS.n6508 0.000502702
R19333 VSS.n6505 VSS.n6499 0.000502702
R19334 VSS.n7020 VSS.n7016 0.000502702
R19335 VSS.n7032 VSS.n7031 0.000502702
R19336 VSS.n7028 VSS.n7015 0.000502702
R19337 VSS.n7065 VSS.n7064 0.000502702
R19338 VSS.n6369 VSS.n6366 0.000502702
R19339 VSS.n6377 VSS.n6367 0.000502702
R19340 VSS.n6439 VSS.n6438 0.000502702
R19341 VSS.n6441 VSS.n6440 0.000502702
R19342 VSS.n6725 VSS.n6724 0.000502702
R19343 VSS.n6736 VSS.n6735 0.000502702
R19344 VSS.n6671 VSS.n6656 0.000502702
R19345 VSS.n5878 VSS.n5877 0.000502702
R19346 VSS.n6035 VSS.n6034 0.000502702
R19347 VSS.n6028 VSS.n6027 0.000502702
R19348 VSS.n6022 VSS.n6021 0.000502702
R19349 VSS.n6046 VSS.n6045 0.000502702
R19350 VSS.n6004 VSS.n6003 0.000502702
R19351 VSS.n6010 VSS.n6009 0.000502702
R19352 VSS.n5862 VSS.n5861 0.000502702
R19353 VSS.n5852 VSS.n5851 0.000502702
R19354 VSS.n5837 VSS.n5836 0.000502702
R19355 VSS.n5830 VSS.n5829 0.000502702
R19356 VSS.n5824 VSS.n5823 0.000502702
R19357 VSS.n5848 VSS.n5847 0.000502702
R19358 VSS.n5806 VSS.n5805 0.000502702
R19359 VSS.n5812 VSS.n5811 0.000502702
R19360 VSS.n5681 VSS.n5680 0.000502702
R19361 VSS.n5671 VSS.n5670 0.000502702
R19362 VSS.n5656 VSS.n5655 0.000502702
R19363 VSS.n5649 VSS.n5648 0.000502702
R19364 VSS.n5643 VSS.n5642 0.000502702
R19365 VSS.n5667 VSS.n5666 0.000502702
R19366 VSS.n5625 VSS.n5624 0.000502702
R19367 VSS.n5631 VSS.n5630 0.000502702
R19368 VSS.n5501 VSS.n5500 0.000502702
R19369 VSS.n5491 VSS.n5490 0.000502702
R19370 VSS.n5476 VSS.n5475 0.000502702
R19371 VSS.n5469 VSS.n5468 0.000502702
R19372 VSS.n5463 VSS.n5462 0.000502702
R19373 VSS.n5487 VSS.n5486 0.000502702
R19374 VSS.n5445 VSS.n5444 0.000502702
R19375 VSS.n5451 VSS.n5450 0.000502702
R19376 VSS.n5321 VSS.n5320 0.000502702
R19377 VSS.n5311 VSS.n5310 0.000502702
R19378 VSS.n5296 VSS.n5295 0.000502702
R19379 VSS.n5289 VSS.n5288 0.000502702
R19380 VSS.n5283 VSS.n5282 0.000502702
R19381 VSS.n5307 VSS.n5306 0.000502702
R19382 VSS.n5265 VSS.n5264 0.000502702
R19383 VSS.n5271 VSS.n5270 0.000502702
R19384 VSS.n10055 VSS.n10054 0.000502702
R19385 VSS.n10045 VSS.n10044 0.000502702
R19386 VSS.n3786 VSS.n3785 0.000502702
R19387 VSS.n3771 VSS.n3770 0.000502702
R19388 VSS.n4615 VSS.n4614 0.000502702
R19389 VSS.n4621 VSS.n4620 0.000502702
R19390 VSS.n6157 VSS.n6156 0.000502702
R19391 VSS.n11096 VSS.n11095 0.000502702
R19392 VSS.n11140 VSS.n11139 0.000502702
R19393 VSS.n3723 VSS.n3722 0.000502702
R19394 VSS.n3729 VSS.n3728 0.000502702
R19395 VSS.n3745 VSS.n3744 0.000502702
R19396 VSS.n3751 VSS.n3750 0.000502702
R19397 VSS.n11128 VSS.n11127 0.000502702
R19398 VSS.n11111 VSS.n11110 0.000502702
R19399 VSS.n6387 VSS.n6386 0.000502702
R19400 VSS.n6365 VSS.n6364 0.000502702
R19401 VSS.n6355 VSS.n6351 0.000502702
R19402 VSS.n6340 VSS.n6334 0.000502702
R19403 VSS.n6404 VSS.n6403 0.000502702
R19404 VSS.n6345 VSS.n6333 0.000502702
R19405 VSS.n11024 VSS.n11023 0.000502702
R19406 VSS.n10992 VSS.n10991 0.000502702
R19407 VSS.n3856 VSS.n3852 0.000502702
R19408 VSS.n3869 VSS.n3868 0.000502702
R19409 VSS.n10976 VSS.n10975 0.000502702
R19410 VSS.n10978 VSS.n10977 0.000502702
R19411 VSS.n10983 VSS.n10982 0.000502702
R19412 VSS.n10952 VSS.n10951 0.000502702
R19413 VSS.n7333 VSS.n7332 0.000502702
R19414 VSS.n7311 VSS.n7310 0.000502702
R19415 VSS.n7301 VSS.n7297 0.000502702
R19416 VSS.n7286 VSS.n7280 0.000502702
R19417 VSS.n7350 VSS.n7349 0.000502702
R19418 VSS.n7291 VSS.n7279 0.000502702
R19419 VSS.n10873 VSS.n10872 0.000502702
R19420 VSS.n3977 VSS.n3976 0.000502702
R19421 VSS.n3983 VSS.n3982 0.000502702
R19422 VSS.n3989 VSS.n3988 0.000502702
R19423 VSS.n4023 VSS.n4022 0.000502702
R19424 VSS.n4011 VSS.n4010 0.000502702
R19425 VSS.n4005 VSS.n4004 0.000502702
R19426 VSS.n4087 VSS.n4086 0.000502702
R19427 VSS.n4145 VSS.n4138 0.000502702
R19428 VSS.n4370 VSS.n4369 0.000502702
R19429 VSS.n4376 VSS.n4375 0.000502702
R19430 VSS.n4338 VSS.n4337 0.000502702
R19431 VSS.n4323 VSS.n4322 0.000502702
R19432 VSS.n4307 VSS.n4261 0.000502702
R19433 VSS.n4315 VSS.n4314 0.000502702
R19434 VSS.n4288 VSS.n4287 0.000502702
R19435 VSS.n4290 VSS.n4289 0.000502702
R19436 VSS.n4297 VSS.n4296 0.000502702
R19437 VSS.n4349 VSS.n4348 0.000502702
R19438 VSS.n4212 VSS.n4208 0.000502702
R19439 VSS.n4217 VSS.n4209 0.000502702
R19440 VSS.n4178 VSS.n4177 0.000502702
R19441 VSS.n4174 VSS.n4161 0.000502702
R19442 VSS.n4432 VSS.n4431 0.000502702
R19443 VSS.n4428 VSS.n4414 0.000502702
R19444 VSS.n4425 VSS.n4424 0.000502702
R19445 VSS.n4124 VSS.n4108 0.000502702
R19446 VSS.n10781 VSS.n10780 0.000502702
R19447 VSS.n4111 VSS.n4107 0.000502702
R19448 VSS.n10769 VSS.n10768 0.000502702
R19449 VSS.n1254 VSS.n1253 0.000502702
R19450 VSS.n1291 VSS.n1290 0.000502702
R19451 VSS.n1027 VSS.n1026 0.000502702
R19452 VSS.n1033 VSS.n1032 0.000502702
R19453 VSS.n1040 VSS.n1039 0.000502702
R19454 VSS.n14324 VSS.n14323 0.000502702
R19455 VSS.n14309 VSS.n14308 0.000502702
R19456 VSS.n565 VSS.n564 0.000502702
R19457 VSS.n14234 VSS.n14233 0.000502702
R19458 VSS.n10699 VSS.n10698 0.000502702
R19459 VSS.n14196 VSS.n14195 0.000502702
R19460 VSS.n12446 VSS.n12445 0.000502702
R19461 VSS.n12440 VSS.n12439 0.000502702
R19462 VSS.n2534 VSS.n2531 0.000502702
R19463 VSS.n2542 VSS.n2532 0.000502702
R19464 VSS.n2473 VSS.n2472 0.000502702
R19465 VSS.n13058 VSS.n13057 0.000502702
R19466 VSS.n2390 VSS.n2389 0.000502702
R19467 VSS.n2382 VSS.n2381 0.000502702
R19468 VSS.n13090 VSS.n13089 0.000502702
R19469 VSS.n13118 VSS.n13117 0.000502702
R19470 VSS.n13127 VSS.n13126 0.000502702
R19471 VSS.n14160 VSS.n14154 0.000502702
R19472 VSS.n14165 VSS.n14155 0.000502702
R19473 VSS.n2419 VSS.n2418 0.000502702
R19474 VSS.n904 VSS.n898 0.000502702
R19475 VSS.n908 VSS.n907 0.000502702
R19476 VSS.n1162 VSS.n1161 0.000502702
R19477 VSS.n14289 VSS.n14288 0.000502702
R19478 VSS.n1549 VSS.n1548 0.000502702
R19479 VSS.n1562 VSS.n1561 0.000502702
R19480 VSS.n13789 VSS.n13788 0.000502702
R19481 VSS.n13795 VSS.n13794 0.000502702
R19482 VSS.n13802 VSS.n13801 0.000502702
R19483 VSS.n742 VSS.n741 0.000502702
R19484 VSS.n748 VSS.n747 0.000502702
R19485 VSS.n755 VSS.n754 0.000502702
R19486 VSS.n645 VSS.n644 0.000502702
R19487 VSS.n14120 VSS.n14119 0.000502702
R19488 VSS.n14076 VSS.n14075 0.000502702
R19489 VSS.n14072 VSS.n14071 0.000502702
R19490 VSS.n14070 VSS.n14069 0.000502702
R19491 VSS.n1644 VSS.n1640 0.000502702
R19492 VSS.n14084 VSS.n14083 0.000502702
R19493 VSS.n1653 VSS.n1641 0.000502702
R19494 VSS.n13702 VSS.n13701 0.000502702
R19495 VSS.n13533 VSS.n13530 0.000502702
R19496 VSS.n13541 VSS.n13531 0.000502702
R19497 VSS.n13890 VSS.n13889 0.000502702
R19498 VSS.n13888 VSS.n13887 0.000502702
R19499 VSS.n850 VSS.n847 0.000502702
R19500 VSS.n860 VSS.n859 0.000502702
R19501 VSS.n1406 VSS.n1405 0.000502702
R19502 VSS.n2250 VSS.n2249 0.000502702
R19503 VSS.n2000 VSS.n1999 0.000502702
R19504 VSS.n2052 VSS.n2051 0.000502702
R19505 VSS.n2045 VSS.n2044 0.000502702
R19506 VSS.n2043 VSS.n2042 0.000502702
R19507 VSS.n2237 VSS.n2236 0.000502702
R19508 VSS.n2185 VSS.n2184 0.000502702
R19509 VSS.n2061 VSS.n2057 0.000502702
R19510 VSS.n2075 VSS.n2074 0.000502702
R19511 VSS.n2101 VSS.n2100 0.000502702
R19512 VSS.n2094 VSS.n2093 0.000502702
R19513 VSS.n2092 VSS.n2091 0.000502702
R19514 VSS.n2172 VSS.n2171 0.000502702
R19515 VSS.n13185 VSS.n13184 0.000502702
R19516 VSS.n1879 VSS.n1878 0.000502702
R19517 VSS.n1875 VSS.n1869 0.000502702
R19518 VSS.n2137 VSS.n2133 0.000502702
R19519 VSS.n2149 VSS.n2148 0.000502702
R19520 VSS.n2145 VSS.n2132 0.000502702
R19521 VSS.n13200 VSS.n13199 0.000502702
R19522 VSS.n1811 VSS.n1810 0.000502702
R19523 VSS.n1803 VSS.n1802 0.000502702
R19524 VSS.n1829 VSS.n1828 0.000502702
R19525 VSS.n13917 VSS.n13916 0.000502702
R19526 VSS.n1962 VSS.n1961 0.000502702
R19527 VSS.n2323 VSS.n2322 0.000502702
R19528 VSS.n2267 VSS.n2266 0.000502702
R19529 VSS.n2712 VSS.n2699 0.000502702
R19530 VSS.n12990 VSS.n12989 0.000502702
R19531 VSS.n2579 VSS.n2578 0.000502702
R19532 VSS.n2659 VSS.n2658 0.000502702
R19533 VSS.n2652 VSS.n2651 0.000502702
R19534 VSS.n2650 VSS.n2649 0.000502702
R19535 VSS.n12967 VSS.n12966 0.000502702
R19536 VSS.n12977 VSS.n12976 0.000502702
R19537 VSS.n12946 VSS.n12945 0.000502702
R19538 VSS.n12942 VSS.n12941 0.000502702
R19539 VSS.n12940 VSS.n12939 0.000502702
R19540 VSS.n2671 VSS.n2667 0.000502702
R19541 VSS.n12954 VSS.n12953 0.000502702
R19542 VSS.n2680 VSS.n2668 0.000502702
R19543 VSS.n2780 VSS.n2779 0.000502702
R19544 VSS.n2820 VSS.n2819 0.000502702
R19545 VSS.n12913 VSS.n12912 0.000502702
R19546 VSS.n2746 VSS.n2742 0.000502702
R19547 VSS.n2760 VSS.n2759 0.000502702
R19548 VSS.n2840 VSS.n2839 0.000502702
R19549 VSS.n2833 VSS.n2832 0.000502702
R19550 VSS.n2831 VSS.n2830 0.000502702
R19551 VSS.n12890 VSS.n12889 0.000502702
R19552 VSS.n12900 VSS.n12899 0.000502702
R19553 VSS.n12869 VSS.n12868 0.000502702
R19554 VSS.n12865 VSS.n12864 0.000502702
R19555 VSS.n12863 VSS.n12862 0.000502702
R19556 VSS.n2860 VSS.n2848 0.000502702
R19557 VSS.n12877 VSS.n12876 0.000502702
R19558 VSS.n2851 VSS.n2847 0.000502702
R19559 VSS.n12643 VSS.n12642 0.000502702
R19560 VSS.n3016 VSS.n3015 0.000502702
R19561 VSS.n3008 VSS.n3007 0.000502702
R19562 VSS.n3034 VSS.n3033 0.000502702
R19563 VSS.n12712 VSS.n12711 0.000502702
R19564 VSS.n2514 VSS.n2513 0.000502702
R19565 VSS.n13028 VSS.n13027 0.000502702
R19566 VSS.n2622 VSS.n2621 0.000502702
R19567 VSS.n12239 VSS.n12238 0.000502702
R19568 VSS.n11680 VSS.n11679 0.000502702
R19569 VSS.n11669 VSS.n11668 0.000502702
R19570 VSS.n11663 VSS.n11662 0.000502702
R19571 VSS.n11639 VSS.n11638 0.000502702
R19572 VSS.n11645 VSS.n11644 0.000502702
R19573 VSS.n11651 VSS.n11650 0.000502702
R19574 VSS.n12223 VSS.n12222 0.000502702
R19575 VSS.n12213 VSS.n12212 0.000502702
R19576 VSS.n11749 VSS.n11748 0.000502702
R19577 VSS.n11738 VSS.n11737 0.000502702
R19578 VSS.n11732 VSS.n11731 0.000502702
R19579 VSS.n11708 VSS.n11707 0.000502702
R19580 VSS.n11714 VSS.n11713 0.000502702
R19581 VSS.n11720 VSS.n11719 0.000502702
R19582 VSS.n12116 VSS.n12115 0.000502702
R19583 VSS.n12106 VSS.n12105 0.000502702
R19584 VSS.n12091 VSS.n12090 0.000502702
R19585 VSS.n12084 VSS.n12083 0.000502702
R19586 VSS.n12078 VSS.n12077 0.000502702
R19587 VSS.n12102 VSS.n12101 0.000502702
R19588 VSS.n12060 VSS.n12059 0.000502702
R19589 VSS.n12066 VSS.n12065 0.000502702
R19590 VSS.n11948 VSS.n11947 0.000502702
R19591 VSS.n11938 VSS.n11937 0.000502702
R19592 VSS.n11881 VSS.n11880 0.000502702
R19593 VSS.n11870 VSS.n11869 0.000502702
R19594 VSS.n11864 VSS.n11863 0.000502702
R19595 VSS.n11840 VSS.n11839 0.000502702
R19596 VSS.n11846 VSS.n11845 0.000502702
R19597 VSS.n11852 VSS.n11851 0.000502702
R19598 VSS.n3520 VSS.n3519 0.000502702
R19599 VSS.n3510 VSS.n3509 0.000502702
R19600 VSS.n3495 VSS.n3494 0.000502702
R19601 VSS.n3488 VSS.n3487 0.000502702
R19602 VSS.n3482 VSS.n3481 0.000502702
R19603 VSS.n3506 VSS.n3505 0.000502702
R19604 VSS.n3464 VSS.n3463 0.000502702
R19605 VSS.n3470 VSS.n3469 0.000502702
R19606 VSS.n3095 VSS.n3094 0.000502702
R19607 VSS.n12609 VSS.n12608 0.000502702
R19608 VSS.n3155 VSS.n3154 0.000502702
R19609 VSS.n3149 VSS.n3148 0.000502702
R19610 VSS.n12377 VSS.n12376 0.000502702
R19611 VSS.n12457 VSS.n12456 0.000502702
R19612 VSS.n3286 VSS.n3285 0.000502702
R19613 VSS.n3276 VSS.n3275 0.000502702
R19614 VSS.n12822 VSS.n12821 0.000502702
R19615 VSS.n2997 VSS.n2996 0.000502702
R19616 VSS.n2981 VSS.n2975 0.000502702
R19617 VSS.n2989 VSS.n2988 0.000502702
R19618 VSS.n12742 VSS.n12736 0.000502702
R19619 VSS.n12749 VSS.n12748 0.000502702
R19620 VSS.n12752 VSS.n12751 0.000502702
R19621 VSS.n12778 VSS.n12777 0.000502702
R19622 VSS.n13988 VSS.n13987 0.000502702
R19623 VSS.n13972 VSS.n1758 0.000502702
R19624 VSS.n13980 VSS.n13979 0.000502702
R19625 VSS.n13953 VSS.n13952 0.000502702
R19626 VSS.n13955 VSS.n13954 0.000502702
R19627 VSS.n13962 VSS.n13961 0.000502702
R19628 VSS.n14021 VSS.n14020 0.000502702
R19629 VSS.n13552 VSS.n13551 0.000502702
R19630 VSS.n13529 VSS.n13528 0.000502702
R19631 VSS.n13519 VSS.n13515 0.000502702
R19632 VSS.n13570 VSS.n13569 0.000502702
R19633 VSS.n13572 VSS.n13571 0.000502702
R19634 VSS.n13575 VSS.n13574 0.000502702
R19635 VSS.n13608 VSS.n13607 0.000502702
R19636 VSS.n13304 VSS.n13303 0.000502702
R19637 VSS.n13310 VSS.n13309 0.000502702
R19638 VSS.n13316 VSS.n13315 0.000502702
R19639 VSS.n13348 VSS.n13347 0.000502702
R19640 VSS.n13338 VSS.n13337 0.000502702
R19641 VSS.n13332 VSS.n13331 0.000502702
R19642 VSS.n13432 VSS.n13431 0.000502702
R19643 VSS.n13477 VSS.n13476 0.000502702
R19644 VSS.n13590 VSS.n13507 0.000502702
R19645 VSS.n1745 VSS.n1742 0.000502702
R19646 VSS.n12801 VSS.n12800 0.000502702
R19647 VSS.n4060 VSS.n4059 0.000502702
R19648 VSS.n10896 VSS.n10895 0.000502702
R19649 VSS.n10941 VSS.n10940 0.000502702
R19650 VSS.n11047 VSS.n11046 0.000502702
R19651 VSS.n9123 VSS.n9122 0.000502702
R19652 VSS.n9654 VSS.n9653 0.000502702
R19653 VSS.n8561 VSS.n8560 0.000502702
R19654 VSS.n8388 VSS.n8387 0.000502702
R19655 VSS.n9638 VSS.n9637 0.000502702
R19656 VSS.n8666 VSS.n8665 0.000502702
R19657 VSS.n8753 VSS.n8752 0.000502702
R19658 VSS.n8773 VSS.n8772 0.000502702
R19659 VSS.n6749 VSS.n6746 0.000502702
R19660 VSS.n8102 VSS.n8099 0.000502702
R19661 VSS.n8106 VSS.n8097 0.000502702
R19662 VSS.n8881 VSS.n8878 0.000502702
R19663 VSS.n9578 VSS.n7550 0.000502702
R19664 VSS.n9401 VSS.n9400 0.000502702
R19665 VSS.n7414 VSS.n7413 0.000502702
R19666 VSS.n3950 VSS.n3949 0.000502702
R19667 VSS.n9450 VSS.n9449 0.000502702
R19668 VSS.n8997 VSS.n8993 0.000502702
R19669 VSS.n9497 VSS.n9490 0.000502702
R19670 VSS.n7253 VSS.n7252 0.000502702
R19671 VSS.n7379 VSS.n7378 0.000502702
R19672 VSS.n9261 VSS.n9260 0.000502702
R19673 VSS.n7870 VSS.n7869 0.000502702
R19674 VSS.n7078 VSS.n7069 0.000502702
R19675 VSS.n9886 VSS.n9885 0.000502702
R19676 VSS.n7989 VSS.n7976 0.000502702
R19677 VSS.n8937 VSS.n8936 0.000502702
R19678 VSS.n6655 VSS.n6654 0.000502702
R19679 VSS.n6894 VSS.n6893 0.000502702
R19680 VSS.n6967 VSS.n6966 0.000502702
R19681 VSS.n6305 VSS.n6296 0.000502702
R19682 VSS.n6448 VSS.n6447 0.000502702
R19683 VSS.n6729 VSS.n6719 0.000502702
R19684 VSS.n5858 VSS.n5857 0.000502702
R19685 VSS.n5677 VSS.n5676 0.000502702
R19686 VSS.n5497 VSS.n5496 0.000502702
R19687 VSS.n5317 VSS.n5316 0.000502702
R19688 VSS.n10051 VSS.n10050 0.000502702
R19689 VSS.n4588 VSS.n4587 0.000502702
R19690 VSS.n4630 VSS.n4629 0.000502702
R19691 VSS.n6051 VSS.n6050 0.000502702
R19692 VSS.n11084 VSS.n11083 0.000502702
R19693 VSS.n4445 VSS.n4444 0.000502702
R19694 VSS.n4372 VSS.n4371 0.000502702
R19695 VSS.n4259 VSS.n4256 0.000502702
R19696 VSS.n4410 VSS.n4409 0.000502702
R19697 VSS.n776 VSS.n775 0.000502702
R19698 VSS.n1260 VSS.n1259 0.000502702
R19699 VSS.n1351 VSS.n1350 0.000502702
R19700 VSS.n1084 VSS.n1083 0.000502702
R19701 VSS.n14330 VSS.n14329 0.000502702
R19702 VSS.n14279 VSS.n14278 0.000502702
R19703 VSS.n1139 VSS.n1136 0.000502702
R19704 VSS.n12434 VSS.n12433 0.000502702
R19705 VSS.n2330 VSS.n2327 0.000502702
R19706 VSS.n1379 VSS.n1372 0.000502702
R19707 VSS.n1555 VSS.n1554 0.000502702
R19708 VSS.n13737 VSS.n13736 0.000502702
R19709 VSS.n13274 VSS.n13273 0.000502702
R19710 VSS.n1622 VSS.n1621 0.000502702
R19711 VSS.n631 VSS.n627 0.000502702
R19712 VSS.n14096 VSS.n14089 0.000502702
R19713 VSS.n13212 VSS.n13203 0.000502702
R19714 VSS.n13897 VSS.n13896 0.000502702
R19715 VSS.n1431 VSS.n1430 0.000502702
R19716 VSS.n1986 VSS.n1982 0.000502702
R19717 VSS.n12682 VSS.n12669 0.000502702
R19718 VSS.n13919 VSS.n1816 0.000502702
R19719 VSS.n1964 VSS.n1947 0.000502702
R19720 VSS.n2565 VSS.n2561 0.000502702
R19721 VSS.n12969 VSS.n12968 0.000502702
R19722 VSS.n2782 VSS.n2769 0.000502702
R19723 VSS.n12892 VSS.n12891 0.000502702
R19724 VSS.n3073 VSS.n3060 0.000502702
R19725 VSS.n12714 VSS.n3021 0.000502702
R19726 VSS.n2516 VSS.n2499 0.000502702
R19727 VSS.n12219 VSS.n12218 0.000502702
R19728 VSS.n12112 VSS.n12111 0.000502702
R19729 VSS.n11944 VSS.n11943 0.000502702
R19730 VSS.n3516 VSS.n3515 0.000502702
R19731 VSS.n3091 VSS.n3090 0.000502702
R19732 VSS.n3122 VSS.n3121 0.000502702
R19733 VSS.n3271 VSS.n3270 0.000502702
R19734 VSS.n3159 VSS.n3158 0.000502702
R19735 VSS.n11635 VSS.n11634 0.000502702
R19736 VSS.n12383 VSS.n12382 0.000502702
R19737 VSS.n12817 VSS.n12816 0.000502702
R19738 VSS.n13468 VSS.n13467 0.000502702
R19739 VSS.n13599 VSS.n13598 0.000502702
R19740 VSS.n14012 VSS.n14011 0.000502702
R19741 VSS.n2933 VSS.n2929 0.000502702
R19742 VSS.n4078 VSS.n4077 0.000502702
R19743 VSS.n3896 VSS.n3892 0.000502702
R19744 VSS.n10928 VSS.n10924 0.000502702
R19745 VSS.n3828 VSS.n3824 0.000502702
R19746 VSS.n9676 VSS.n9675 0.000502702
R19747 VSS.n9670 VSS.n9669 0.000502702
R19748 VSS.n9694 VSS.n9693 0.000502702
R19749 VSS.n9135 VSS.n9134 0.000502702
R19750 VSS.n9129 VSS.n9128 0.000502702
R19751 VSS.n9141 VSS.n9140 0.000502702
R19752 VSS.n9042 VSS.n9041 0.000502702
R19753 VSS.n9036 VSS.n9035 0.000502702
R19754 VSS.n8355 VSS.n8354 0.000502702
R19755 VSS.n8361 VSS.n8360 0.000502702
R19756 VSS.n8480 VSS.n8479 0.000502702
R19757 VSS.n8474 VSS.n8473 0.000502702
R19758 VSS.n8508 VSS.n8507 0.000502702
R19759 VSS.n8500 VSS.n8491 0.000502702
R19760 VSS.n8496 VSS.n8495 0.000502702
R19761 VSS.n8371 VSS.n8369 0.000502702
R19762 VSS.n8379 VSS.n8365 0.000502702
R19763 VSS.n8407 VSS.n8406 0.000502702
R19764 VSS.n8399 VSS.n8390 0.000502702
R19765 VSS.n8395 VSS.n8394 0.000502702
R19766 VSS.n8688 VSS.n8687 0.000502702
R19767 VSS.n8682 VSS.n8681 0.000502702
R19768 VSS.n8706 VSS.n8705 0.000502702
R19769 VSS.n9632 VSS.n9631 0.000502702
R19770 VSS.n9626 VSS.n9625 0.000502702
R19771 VSS.n9614 VSS.n9613 0.000502702
R19772 VSS.n7543 VSS.n7542 0.000502702
R19773 VSS.n7537 VSS.n7536 0.000502702
R19774 VSS.n8309 VSS.n8308 0.000502702
R19775 VSS.n8315 VSS.n8314 0.000502702
R19776 VSS.n8736 VSS.n8735 0.000502702
R19777 VSS.n8583 VSS.n8582 0.000502702
R19778 VSS.n8577 VSS.n8576 0.000502702
R19779 VSS.n8619 VSS.n8618 0.000502702
R19780 VSS.n8297 VSS.n8296 0.000502702
R19781 VSS.n8291 VSS.n8290 0.000502702
R19782 VSS.n8252 VSS.n8246 0.000502702
R19783 VSS.n8260 VSS.n8259 0.000502702
R19784 VSS.n8238 VSS.n8237 0.000502702
R19785 VSS.n8235 VSS.n8223 0.000502702
R19786 VSS.n8230 VSS.n8229 0.000502702
R19787 VSS.n8197 VSS.n8193 0.000502702
R19788 VSS.n8205 VSS.n8204 0.000502702
R19789 VSS.n6201 VSS.n6200 0.000502702
R19790 VSS.n9982 VSS.n9981 0.000502702
R19791 VSS.n6221 VSS.n6212 0.000502702
R19792 VSS.n6226 VSS.n6225 0.000502702
R19793 VSS.n6758 VSS.n6757 0.000502702
R19794 VSS.n6753 VSS.n6717 0.000502702
R19795 VSS.n6766 VSS.n6765 0.000502702
R19796 VSS.n6701 VSS.n6691 0.000502702
R19797 VSS.n6706 VSS.n6705 0.000502702
R19798 VSS.n9964 VSS.n9963 0.000502702
R19799 VSS.n8156 VSS.n8155 0.000502702
R19800 VSS.n8031 VSS.n8015 0.000502702
R19801 VSS.n8029 VSS.n8027 0.000502702
R19802 VSS.n8111 VSS.n8110 0.000502702
R19803 VSS.n8089 VSS.n8088 0.000502702
R19804 VSS.n8086 VSS.n8085 0.000502702
R19805 VSS.n8081 VSS.n8076 0.000502702
R19806 VSS.n8132 VSS.n8129 0.000502702
R19807 VSS.n8138 VSS.n8133 0.000502702
R19808 VSS.n8073 VSS.n8072 0.000502702
R19809 VSS.n8063 VSS.n8050 0.000502702
R19810 VSS.n8061 VSS.n8055 0.000502702
R19811 VSS.n8890 VSS.n8889 0.000502702
R19812 VSS.n8885 VSS.n7974 0.000502702
R19813 VSS.n8898 VSS.n8897 0.000502702
R19814 VSS.n7958 VSS.n7947 0.000502702
R19815 VSS.n7963 VSS.n7962 0.000502702
R19816 VSS.n8862 VSS.n8850 0.000502702
R19817 VSS.n8812 VSS.n8811 0.000502702
R19818 VSS.n8809 VSS.n8808 0.000502702
R19819 VSS.n8803 VSS.n8796 0.000502702
R19820 VSS.n8165 VSS.n8161 0.000502702
R19821 VSS.n8173 VSS.n8172 0.000502702
R19822 VSS.n8267 VSS.n8265 0.000502702
R19823 VSS.n8275 VSS.n8261 0.000502702
R19824 VSS.n8284 VSS.n8283 0.000502702
R19825 VSS.n9564 VSS.n9563 0.000502702
R19826 VSS.n9571 VSS.n9570 0.000502702
R19827 VSS.n9573 VSS.n9572 0.000502702
R19828 VSS.n9586 VSS.n9585 0.000502702
R19829 VSS.n9595 VSS.n9594 0.000502702
R19830 VSS.n8531 VSS.n8530 0.000502702
R19831 VSS.n8537 VSS.n8536 0.000502702
R19832 VSS.n8543 VSS.n8542 0.000502702
R19833 VSS.n8457 VSS.n8456 0.000502702
R19834 VSS.n9383 VSS.n9382 0.000502702
R19835 VSS.n9377 VSS.n9376 0.000502702
R19836 VSS.n9419 VSS.n9418 0.000502702
R19837 VSS.n9791 VSS.n9790 0.000502702
R19838 VSS.n7398 VSS.n7397 0.000502702
R19839 VSS.n7404 VSS.n7403 0.000502702
R19840 VSS.n7386 VSS.n7385 0.000502702
R19841 VSS.n9778 VSS.n9777 0.000502702
R19842 VSS.n7440 VSS.n7439 0.000502702
R19843 VSS.n7434 VSS.n7433 0.000502702
R19844 VSS.n7476 VSS.n7475 0.000502702
R19845 VSS.n10838 VSS.n10837 0.000502702
R19846 VSS.n3934 VSS.n3933 0.000502702
R19847 VSS.n3940 VSS.n3939 0.000502702
R19848 VSS.n3922 VSS.n3921 0.000502702
R19849 VSS.n10825 VSS.n10824 0.000502702
R19850 VSS.n9343 VSS.n9342 0.000502702
R19851 VSS.n9349 VSS.n9348 0.000502702
R19852 VSS.n9433 VSS.n9432 0.000502702
R19853 VSS.n9077 VSS.n9076 0.000502702
R19854 VSS.n9071 VSS.n9070 0.000502702
R19855 VSS.n9113 VSS.n9112 0.000502702
R19856 VSS.n9331 VSS.n9330 0.000502702
R19857 VSS.n9325 VSS.n9324 0.000502702
R19858 VSS.n9279 VSS.n9278 0.000502702
R19859 VSS.n9281 VSS.n9280 0.000502702
R19860 VSS.n9288 VSS.n9287 0.000502702
R19861 VSS.n9311 VSS.n9294 0.000502702
R19862 VSS.n9306 VSS.n9305 0.000502702
R19863 VSS.n9304 VSS.n9303 0.000502702
R19864 VSS.n9499 VSS.n9498 0.000502702
R19865 VSS.n9508 VSS.n9507 0.000502702
R19866 VSS.n7224 VSS.n7216 0.000502702
R19867 VSS.n7239 VSS.n7238 0.000502702
R19868 VSS.n7228 VSS.n7217 0.000502702
R19869 VSS.n9822 VSS.n9821 0.000502702
R19870 VSS.n9820 VSS.n9819 0.000502702
R19871 VSS.n7255 VSS.n7211 0.000502702
R19872 VSS.n7251 VSS.n7250 0.000502702
R19873 VSS.n7365 VSS.n7364 0.000502702
R19874 VSS.n7362 VSS.n7361 0.000502702
R19875 VSS.n7357 VSS.n7352 0.000502702
R19876 VSS.n7328 VSS.n7327 0.000502702
R19877 VSS.n9177 VSS.n9174 0.000502702
R19878 VSS.n9179 VSS.n9159 0.000502702
R19879 VSS.n9269 VSS.n9268 0.000502702
R19880 VSS.n9199 VSS.n9198 0.000502702
R19881 VSS.n9197 VSS.n9190 0.000502702
R19882 VSS.n9208 VSS.n9207 0.000502702
R19883 VSS.n9257 VSS.n9254 0.000502702
R19884 VSS.n9253 VSS.n9252 0.000502702
R19885 VSS.n7846 VSS.n7808 0.000502702
R19886 VSS.n8962 VSS.n8961 0.000502702
R19887 VSS.n7821 VSS.n7809 0.000502702
R19888 VSS.n7841 VSS.n7838 0.000502702
R19889 VSS.n7837 VSS.n7836 0.000502702
R19890 VSS.n7737 VSS.n7729 0.000502702
R19891 VSS.n7752 VSS.n7751 0.000502702
R19892 VSS.n7741 VSS.n7730 0.000502702
R19893 VSS.n7795 VSS.n7794 0.000502702
R19894 VSS.n7793 VSS.n7792 0.000502702
R19895 VSS.n7695 VSS.n7694 0.000502702
R19896 VSS.n7681 VSS.n7677 0.000502702
R19897 VSS.n7687 VSS.n7686 0.000502702
R19898 VSS.n7716 VSS.n7715 0.000502702
R19899 VSS.n7714 VSS.n7713 0.000502702
R19900 VSS.n9897 VSS.n9896 0.000502702
R19901 VSS.n7083 VSS.n7082 0.000502702
R19902 VSS.n7135 VSS.n7134 0.000502702
R19903 VSS.n7131 VSS.n7128 0.000502702
R19904 VSS.n7127 VSS.n7126 0.000502702
R19905 VSS.n7110 VSS.n7107 0.000502702
R19906 VSS.n7927 VSS.n7926 0.000502702
R19907 VSS.n7931 VSS.n7928 0.000502702
R19908 VSS.n7936 VSS.n7935 0.000502702
R19909 VSS.n8918 VSS.n8917 0.000502702
R19910 VSS.n8915 VSS.n8914 0.000502702
R19911 VSS.n8909 VSS.n8902 0.000502702
R19912 VSS.n7875 VSS.n7871 0.000502702
R19913 VSS.n7884 VSS.n7883 0.000502702
R19914 VSS.n6912 VSS.n6911 0.000502702
R19915 VSS.n6621 VSS.n6618 0.000502702
R19916 VSS.n6985 VSS.n6984 0.000502702
R19917 VSS.n6573 VSS.n6570 0.000502702
R19918 VSS.n6535 VSS.n6510 0.000502702
R19919 VSS.n7044 VSS.n7043 0.000502702
R19920 VSS.n6523 VSS.n6511 0.000502702
R19921 VSS.n7013 VSS.n7012 0.000502702
R19922 VSS.n7006 VSS.n7001 0.000502702
R19923 VSS.n6293 VSS.n6292 0.000502702
R19924 VSS.n6474 VSS.n6473 0.000502702
R19925 VSS.n6472 VSS.n6471 0.000502702
R19926 VSS.n6285 VSS.n6270 0.000502702
R19927 VSS.n6283 VSS.n6280 0.000502702
R19928 VSS.n6459 VSS.n6458 0.000502702
R19929 VSS.n6310 VSS.n6309 0.000502702
R19930 VSS.n6419 VSS.n6418 0.000502702
R19931 VSS.n6416 VSS.n6415 0.000502702
R19932 VSS.n6411 VSS.n6406 0.000502702
R19933 VSS.n6382 VSS.n6381 0.000502702
R19934 VSS.n6825 VSS.n6824 0.000502702
R19935 VSS.n6827 VSS.n6826 0.000502702
R19936 VSS.n6834 VSS.n6833 0.000502702
R19937 VSS.n6783 VSS.n6782 0.000502702
R19938 VSS.n6780 VSS.n6779 0.000502702
R19939 VSS.n6775 VSS.n6770 0.000502702
R19940 VSS.n6669 VSS.n6666 0.000502702
R19941 VSS.n6845 VSS.n6844 0.000502702
R19942 VSS.n5901 VSS.n5900 0.000502702
R19943 VSS.n5872 VSS.n5871 0.000502702
R19944 VSS.n5720 VSS.n5719 0.000502702
R19945 VSS.n5691 VSS.n5690 0.000502702
R19946 VSS.n5540 VSS.n5539 0.000502702
R19947 VSS.n5511 VSS.n5510 0.000502702
R19948 VSS.n5360 VSS.n5359 0.000502702
R19949 VSS.n5331 VSS.n5330 0.000502702
R19950 VSS.n10094 VSS.n10093 0.000502702
R19951 VSS.n10065 VSS.n10064 0.000502702
R19952 VSS.n4582 VSS.n4581 0.000502702
R19953 VSS.n4594 VSS.n4593 0.000502702
R19954 VSS.n3812 VSS.n3811 0.000502702
R19955 VSS.n3804 VSS.n3803 0.000502702
R19956 VSS.n3798 VSS.n3797 0.000502702
R19957 VSS.n3777 VSS.n3776 0.000502702
R19958 VSS.n6057 VSS.n6056 0.000502702
R19959 VSS.n6065 VSS.n6064 0.000502702
R19960 VSS.n6083 VSS.n6082 0.000502702
R19961 VSS.n5984 VSS.n5983 0.000502702
R19962 VSS.n5978 VSS.n5977 0.000502702
R19963 VSS.n6178 VSS.n6177 0.000502702
R19964 VSS.n6172 VSS.n6171 0.000502702
R19965 VSS.n11102 VSS.n11101 0.000502702
R19966 VSS.n11068 VSS.n11067 0.000502702
R19967 VSS.n11062 VSS.n11061 0.000502702
R19968 VSS.n11018 VSS.n11017 0.000502702
R19969 VSS.n11016 VSS.n11015 0.000502702
R19970 VSS.n10912 VSS.n10899 0.000502702
R19971 VSS.n10910 VSS.n10904 0.000502702
R19972 VSS.n10867 VSS.n10866 0.000502702
R19973 VSS.n10865 VSS.n10864 0.000502702
R19974 VSS.n4051 VSS.n4050 0.000502702
R19975 VSS.n4045 VSS.n4044 0.000502702
R19976 VSS.n4151 VSS.n4150 0.000502702
R19977 VSS.n4400 VSS.n4399 0.000502702
R19978 VSS.n4395 VSS.n4392 0.000502702
R19979 VSS.n4391 VSS.n4390 0.000502702
R19980 VSS.n4340 VSS.n4339 0.000502702
R19981 VSS.n4247 VSS.n4229 0.000502702
R19982 VSS.n4245 VSS.n4242 0.000502702
R19983 VSS.n4224 VSS.n4223 0.000502702
R19984 VSS.n10761 VSS.n10760 0.000502702
R19985 VSS.n10759 VSS.n10758 0.000502702
R19986 VSS.n1282 VSS.n1281 0.000502702
R19987 VSS.n1276 VSS.n1275 0.000502702
R19988 VSS.n1300 VSS.n1299 0.000502702
R19989 VSS.n788 VSS.n787 0.000502702
R19990 VSS.n782 VSS.n781 0.000502702
R19991 VSS.n794 VSS.n793 0.000502702
R19992 VSS.n676 VSS.n675 0.000502702
R19993 VSS.n670 VSS.n669 0.000502702
R19994 VSS.n1220 VSS.n1219 0.000502702
R19995 VSS.n1226 VSS.n1225 0.000502702
R19996 VSS.n1334 VSS.n1333 0.000502702
R19997 VSS.n1015 VSS.n1014 0.000502702
R19998 VSS.n1009 VSS.n1008 0.000502702
R19999 VSS.n1051 VSS.n1050 0.000502702
R20000 VSS.n1208 VSS.n1207 0.000502702
R20001 VSS.n1202 VSS.n1201 0.000502702
R20002 VSS.n968 VSS.n967 0.000502702
R20003 VSS.n974 VSS.n973 0.000502702
R20004 VSS.n14224 VSS.n14223 0.000502702
R20005 VSS.n14219 VSS.n14216 0.000502702
R20006 VSS.n14215 VSS.n14214 0.000502702
R20007 VSS.n567 VSS.n544 0.000502702
R20008 VSS.n10708 VSS.n10707 0.000502702
R20009 VSS.n10685 VSS.n10684 0.000502702
R20010 VSS.n10679 VSS.n10678 0.000502702
R20011 VSS.n14273 VSS.n14272 0.000502702
R20012 VSS.n14267 VSS.n14266 0.000502702
R20013 VSS.n14255 VSS.n14254 0.000502702
R20014 VSS.n531 VSS.n530 0.000502702
R20015 VSS.n525 VSS.n524 0.000502702
R20016 VSS.n10666 VSS.n10665 0.000502702
R20017 VSS.n10660 VSS.n10659 0.000502702
R20018 VSS.n14206 VSS.n14205 0.000502702
R20019 VSS.n599 VSS.n583 0.000502702
R20020 VSS.n597 VSS.n595 0.000502702
R20021 VSS.n1148 VSS.n1147 0.000502702
R20022 VSS.n1143 VSS.n935 0.000502702
R20023 VSS.n1156 VSS.n1155 0.000502702
R20024 VSS.n919 VSS.n909 0.000502702
R20025 VSS.n924 VSS.n923 0.000502702
R20026 VSS.n14182 VSS.n14179 0.000502702
R20027 VSS.n14188 VSS.n14183 0.000502702
R20028 VSS.n12419 VSS.n12418 0.000502702
R20029 VSS.n12410 VSS.n12397 0.000502702
R20030 VSS.n12408 VSS.n12402 0.000502702
R20031 VSS.n13043 VSS.n13042 0.000502702
R20032 VSS.n13040 VSS.n13039 0.000502702
R20033 VSS.n13035 VSS.n13030 0.000502702
R20034 VSS.n2547 VSS.n2546 0.000502702
R20035 VSS.n2475 VSS.n2460 0.000502702
R20036 VSS.n2448 VSS.n2447 0.000502702
R20037 VSS.n2445 VSS.n2444 0.000502702
R20038 VSS.n2437 VSS.n2430 0.000502702
R20039 VSS.n13099 VSS.n2350 0.000502702
R20040 VSS.n13105 VSS.n13104 0.000502702
R20041 VSS.n2368 VSS.n2351 0.000502702
R20042 VSS.n2386 VSS.n2383 0.000502702
R20043 VSS.n13076 VSS.n13073 0.000502702
R20044 VSS.n13082 VSS.n13077 0.000502702
R20045 VSS.n13138 VSS.n13137 0.000502702
R20046 VSS.n1919 VSS.n1910 0.000502702
R20047 VSS.n1924 VSS.n1923 0.000502702
R20048 VSS.n2339 VSS.n2338 0.000502702
R20049 VSS.n2334 VSS.n1945 0.000502702
R20050 VSS.n2296 VSS.n2295 0.000502702
R20051 VSS.n2291 VSS.n2280 0.000502702
R20052 VSS.n2287 VSS.n2284 0.000502702
R20053 VSS.n13120 VSS.n13119 0.000502702
R20054 VSS.n14172 VSS.n14171 0.000502702
R20055 VSS.n2415 VSS.n2397 0.000502702
R20056 VSS.n2412 VSS.n2409 0.000502702
R20057 VSS.n942 VSS.n941 0.000502702
R20058 VSS.n946 VSS.n937 0.000502702
R20059 VSS.n954 VSS.n953 0.000502702
R20060 VSS.n1400 VSS.n1399 0.000502702
R20061 VSS.n870 VSS.n861 0.000502702
R20062 VSS.n875 VSS.n874 0.000502702
R20063 VSS.n1381 VSS.n1380 0.000502702
R20064 VSS.n1390 VSS.n1389 0.000502702
R20065 VSS.n1112 VSS.n1111 0.000502702
R20066 VSS.n1088 VSS.n1087 0.000502702
R20067 VSS.n1094 VSS.n1093 0.000502702
R20068 VSS.n14295 VSS.n14294 0.000502702
R20069 VSS.n14336 VSS.n14335 0.000502702
R20070 VSS.n1537 VSS.n1536 0.000502702
R20071 VSS.n1531 VSS.n1530 0.000502702
R20072 VSS.n1573 VSS.n1572 0.000502702
R20073 VSS.n13859 VSS.n13858 0.000502702
R20074 VSS.n13721 VSS.n13720 0.000502702
R20075 VSS.n13727 VSS.n13726 0.000502702
R20076 VSS.n13709 VSS.n13708 0.000502702
R20077 VSS.n13846 VSS.n13845 0.000502702
R20078 VSS.n13777 VSS.n13776 0.000502702
R20079 VSS.n13771 VSS.n13770 0.000502702
R20080 VSS.n13813 VSS.n13812 0.000502702
R20081 VSS.n13394 VSS.n13393 0.000502702
R20082 VSS.n13258 VSS.n13257 0.000502702
R20083 VSS.n13264 VSS.n13263 0.000502702
R20084 VSS.n13246 VSS.n13245 0.000502702
R20085 VSS.n13381 VSS.n13380 0.000502702
R20086 VSS.n1489 VSS.n1488 0.000502702
R20087 VSS.n1495 VSS.n1494 0.000502702
R20088 VSS.n1605 VSS.n1604 0.000502702
R20089 VSS.n730 VSS.n729 0.000502702
R20090 VSS.n724 VSS.n723 0.000502702
R20091 VSS.n766 VSS.n765 0.000502702
R20092 VSS.n1477 VSS.n1476 0.000502702
R20093 VSS.n1471 VSS.n1470 0.000502702
R20094 VSS.n1449 VSS.n1448 0.000502702
R20095 VSS.n1451 VSS.n1450 0.000502702
R20096 VSS.n1458 VSS.n1457 0.000502702
R20097 VSS.n1684 VSS.n1672 0.000502702
R20098 VSS.n1695 VSS.n1694 0.000502702
R20099 VSS.n1680 VSS.n1673 0.000502702
R20100 VSS.n14098 VSS.n14097 0.000502702
R20101 VSS.n14107 VSS.n14106 0.000502702
R20102 VSS.n13673 VSS.n13672 0.000502702
R20103 VSS.n13687 VSS.n13686 0.000502702
R20104 VSS.n13685 VSS.n13684 0.000502702
R20105 VSS.n13664 VSS.n13651 0.000502702
R20106 VSS.n13662 VSS.n13656 0.000502702
R20107 VSS.n13908 VSS.n13907 0.000502702
R20108 VSS.n13217 VSS.n13216 0.000502702
R20109 VSS.n13641 VSS.n13640 0.000502702
R20110 VSS.n13638 VSS.n13637 0.000502702
R20111 VSS.n13633 VSS.n13628 0.000502702
R20112 VSS.n13546 VSS.n13545 0.000502702
R20113 VSS.n830 VSS.n827 0.000502702
R20114 VSS.n832 VSS.n812 0.000502702
R20115 VSS.n1439 VSS.n1438 0.000502702
R20116 VSS.n1178 VSS.n1176 0.000502702
R20117 VSS.n1186 VSS.n1172 0.000502702
R20118 VSS.n1195 VSS.n1194 0.000502702
R20119 VSS.n1427 VSS.n1424 0.000502702
R20120 VSS.n1423 VSS.n1422 0.000502702
R20121 VSS.n2207 VSS.n2206 0.000502702
R20122 VSS.n2204 VSS.n2203 0.000502702
R20123 VSS.n2193 VSS.n2189 0.000502702
R20124 VSS.n2229 VSS.n2228 0.000502702
R20125 VSS.n2227 VSS.n2226 0.000502702
R20126 VSS.n2123 VSS.n2122 0.000502702
R20127 VSS.n2109 VSS.n2105 0.000502702
R20128 VSS.n2115 VSS.n2114 0.000502702
R20129 VSS.n2164 VSS.n2163 0.000502702
R20130 VSS.n2162 VSS.n2161 0.000502702
R20131 VSS.n12652 VSS.n12645 0.000502702
R20132 VSS.n12667 VSS.n12666 0.000502702
R20133 VSS.n12656 VSS.n12646 0.000502702
R20134 VSS.n1845 VSS.n1830 0.000502702
R20135 VSS.n1843 VSS.n1840 0.000502702
R20136 VSS.n12692 VSS.n12691 0.000502702
R20137 VSS.n12680 VSS.n12674 0.000502702
R20138 VSS.n13933 VSS.n1771 0.000502702
R20139 VSS.n13939 VSS.n13938 0.000502702
R20140 VSS.n1789 VSS.n1772 0.000502702
R20141 VSS.n1807 VSS.n1804 0.000502702
R20142 VSS.n2021 VSS.n2015 0.000502702
R20143 VSS.n2023 VSS.n2010 0.000502702
R20144 VSS.n2033 VSS.n2032 0.000502702
R20145 VSS.n2316 VSS.n2315 0.000502702
R20146 VSS.n2311 VSS.n2308 0.000502702
R20147 VSS.n2307 VSS.n2306 0.000502702
R20148 VSS.n2265 VSS.n2264 0.000502702
R20149 VSS.n2275 VSS.n2274 0.000502702
R20150 VSS.n2722 VSS.n2721 0.000502702
R20151 VSS.n2710 VSS.n2704 0.000502702
R20152 VSS.n2806 VSS.n2789 0.000502702
R20153 VSS.n2802 VSS.n2801 0.000502702
R20154 VSS.n2902 VSS.n2901 0.000502702
R20155 VSS.n2890 VSS.n2884 0.000502702
R20156 VSS.n3057 VSS.n3056 0.000502702
R20157 VSS.n12628 VSS.n12627 0.000502702
R20158 VSS.n12626 VSS.n12625 0.000502702
R20159 VSS.n3048 VSS.n3035 0.000502702
R20160 VSS.n3046 VSS.n3040 0.000502702
R20161 VSS.n3083 VSS.n3082 0.000502702
R20162 VSS.n3071 VSS.n3065 0.000502702
R20163 VSS.n12728 VSS.n2949 0.000502702
R20164 VSS.n12734 VSS.n12733 0.000502702
R20165 VSS.n2967 VSS.n2950 0.000502702
R20166 VSS.n3012 VSS.n3009 0.000502702
R20167 VSS.n2601 VSS.n2595 0.000502702
R20168 VSS.n2603 VSS.n2589 0.000502702
R20169 VSS.n2640 VSS.n2639 0.000502702
R20170 VSS.n13021 VSS.n13020 0.000502702
R20171 VSS.n13016 VSS.n13013 0.000502702
R20172 VSS.n13012 VSS.n13011 0.000502702
R20173 VSS.n2620 VSS.n2619 0.000502702
R20174 VSS.n2630 VSS.n2629 0.000502702
R20175 VSS.n12262 VSS.n12261 0.000502702
R20176 VSS.n12233 VSS.n12232 0.000502702
R20177 VSS.n12155 VSS.n12154 0.000502702
R20178 VSS.n12126 VSS.n12125 0.000502702
R20179 VSS.n11987 VSS.n11986 0.000502702
R20180 VSS.n11958 VSS.n11957 0.000502702
R20181 VSS.n3559 VSS.n3558 0.000502702
R20182 VSS.n3530 VSS.n3529 0.000502702
R20183 VSS.n12588 VSS.n12587 0.000502702
R20184 VSS.n3105 VSS.n3104 0.000502702
R20185 VSS.n3170 VSS.n3169 0.000502702
R20186 VSS.n3128 VSS.n3127 0.000502702
R20187 VSS.n3260 VSS.n3259 0.000502702
R20188 VSS.n3254 VSS.n3253 0.000502702
R20189 VSS.n3246 VSS.n3245 0.000502702
R20190 VSS.n3239 VSS.n3238 0.000502702
R20191 VSS.n3233 VSS.n3232 0.000502702
R20192 VSS.n11607 VSS.n11606 0.000502702
R20193 VSS.n11615 VSS.n11614 0.000502702
R20194 VSS.n11599 VSS.n11598 0.000502702
R20195 VSS.n11593 VSS.n11592 0.000502702
R20196 VSS.n11587 VSS.n11586 0.000502702
R20197 VSS.n12772 VSS.n12771 0.000502702
R20198 VSS.n12770 VSS.n12769 0.000502702
R20199 VSS.n1733 VSS.n1715 0.000502702
R20200 VSS.n1731 VSS.n1728 0.000502702
R20201 VSS.n13498 VSS.n13480 0.000502702
R20202 VSS.n13496 VSS.n13493 0.000502702
R20203 VSS.n13448 VSS.n13447 0.000502702
R20204 VSS.n13442 VSS.n13441 0.000502702
R20205 VSS.n12465 VSS.n12464 0.000502311
R20206 VSS.n6149 VSS.n6148 0.000502311
R20207 VSS.n5966 VSS.n5965 0.000502311
R20208 VSS.n5785 VSS.n5784 0.000502311
R20209 VSS.n4092 VSS.n4091 0.000502311
R20210 VSS.n1243 VSS.n1242 0.000502311
R20211 VSS.n13754 VSS.n13753 0.000502311
R20212 VSS.n13834 VSS.n13833 0.000502311
R20213 VSS.n1594 VSS.n1593 0.000502311
R20214 VSS.n3196 VSS.n3195 0.000502311
R20215 VSS.n13424 VSS.n13423 0.000502311
R20216 VSS.n1513 VSS.n1512 0.000502311
R20217 VSS.n8428 VSS.n8427 0.000502311
R20218 VSS.n8624 VSS.n8623 0.000502311
R20219 VSS.n8713 VSS.n8712 0.000502311
R20220 VSS.n9699 VSS.n9698 0.000502311
R20221 VSS.n9057 VSS.n9056 0.000502311
R20222 VSS.n7484 VSS.n7483 0.000502311
R20223 VSS.n4030 VSS.n4029 0.000502311
R20224 VSS.n9768 VSS.n9767 0.000502311
R20225 VSS.n9422 VSS.n9421 0.000502311
R20226 VSS.n5604 VSS.n5603 0.000502311
R20227 VSS.n5424 VSS.n5423 0.000502311
R20228 VSS.n5244 VSS.n5243 0.000502311
R20229 VSS.n10102 VSS.n10101 0.000502311
R20230 VSS.n11145 VSS.n11144 0.000502311
R20231 VSS.n11520 VSS.n11519 0.000502311
R20232 VSS.n10647 VSS.n10646 0.000502311
R20233 VSS.n10717 VSS.n10716 0.000502311
R20234 VSS.n992 VSS.n991 0.000502311
R20235 VSS.n14358 VSS.n14357 0.000502311
R20236 VSS.n14372 VSS.n14371 0.000502311
R20237 VSS.n1072 VSS.n1071 0.000502311
R20238 VSS.n1322 VSS.n1321 0.000502311
R20239 VSS.n465 VSS.n464 0.000502311
R20240 VSS.n13292 VSS.n13291 0.000502311
R20241 VSS.n13369 VSS.n13368 0.000502311
R20242 VSS.n12338 VSS.n12337 0.000502311
R20243 VSS.n12205 VSS.n12204 0.000502311
R20244 VSS.n12041 VSS.n12040 0.000502311
R20245 VSS.n11928 VSS.n11927 0.000502311
R20246 VSS.n3443 VSS.n3442 0.000502311
R20247 VSS.n12578 VSS.n12577 0.000502311
R20248 VSS.n3211 VSS.n3210 0.000502311
R20249 VSS.n10636 VSS.n10635 0.000501541
R20250 VSS.n12025 VSS.n12024 0.000501541
R20251 VSS.n12019 VSS.n12018 0.000501541
R20252 VSS.n12008 VSS.n12007 0.000501541
R20253 VSS.n12002 VSS.n12001 0.000501541
R20254 VSS.n11894 VSS.n11893 0.000501541
R20255 VSS.n11888 VSS.n11887 0.000501541
R20256 VSS.n3579 VSS.n3578 0.000501541
R20257 VSS.n3573 VSS.n3572 0.000501541
R20258 VSS.n3409 VSS.n3408 0.000501541
R20259 VSS.n3403 VSS.n3402 0.000501541
R20260 VSS.n3326 VSS.n3325 0.000501541
R20261 VSS.n3366 VSS.n3365 0.000501541
R20262 VSS.n12564 VSS.n12563 0.000501541
R20263 VSS.n12557 VSS.n12556 0.000501541
R20264 VSS.n3181 VSS.n3180 0.000501541
R20265 VSS.n3311 VSS.n3310 0.000501541
R20266 VSS.n14482 VSS.n14481 0.000501541
R20267 VSS.n14473 VSS.n14467 0.000501541
R20268 VSS.n14500 VSS.n14499 0.000501541
R20269 VSS.n12193 VSS.n12192 0.000501541
R20270 VSS.n12187 VSS.n12186 0.000501541
R20271 VSS.n12175 VSS.n12174 0.000501541
R20272 VSS.n12169 VSS.n12168 0.000501541
R20273 VSS.n11175 VSS.n11174 0.000501541
R20274 VSS.n11179 VSS.n11178 0.000501541
R20275 VSS.n11159 VSS.n11158 0.000501541
R20276 VSS.n11163 VSS.n11162 0.000501541
R20277 VSS.n10161 VSS.n10160 0.000501541
R20278 VSS.n10155 VSS.n10154 0.000501541
R20279 VSS.n10116 VSS.n10115 0.000501541
R20280 VSS.n10120 VSS.n10119 0.000501541
R20281 VSS.n5213 VSS.n5212 0.000501541
R20282 VSS.n5207 VSS.n5206 0.000501541
R20283 VSS.n5229 VSS.n5228 0.000501541
R20284 VSS.n5223 VSS.n5222 0.000501541
R20285 VSS.n5393 VSS.n5392 0.000501541
R20286 VSS.n5387 VSS.n5386 0.000501541
R20287 VSS.n5409 VSS.n5408 0.000501541
R20288 VSS.n5403 VSS.n5402 0.000501541
R20289 VSS.n5573 VSS.n5572 0.000501541
R20290 VSS.n5567 VSS.n5566 0.000501541
R20291 VSS.n5589 VSS.n5588 0.000501541
R20292 VSS.n5583 VSS.n5582 0.000501541
R20293 VSS.n5753 VSS.n5752 0.000501541
R20294 VSS.n5747 VSS.n5746 0.000501541
R20295 VSS.n5769 VSS.n5768 0.000501541
R20296 VSS.n5763 VSS.n5762 0.000501541
R20297 VSS.n5934 VSS.n5933 0.000501541
R20298 VSS.n5928 VSS.n5927 0.000501541
R20299 VSS.n5950 VSS.n5949 0.000501541
R20300 VSS.n5944 VSS.n5943 0.000501541
R20301 VSS.n6116 VSS.n6115 0.000501541
R20302 VSS.n6110 VSS.n6109 0.000501541
R20303 VSS.n6132 VSS.n6131 0.000501541
R20304 VSS.n6126 VSS.n6125 0.000501541
R20305 VSS.n3610 VSS.n3609 0.000501541
R20306 VSS.n12318 VSS.n12317 0.000501541
R20307 VSS.n12312 VSS.n12311 0.000501541
R20308 VSS.n12290 VSS.n12289 0.000501541
R20309 VSS.n12284 VSS.n12283 0.000501541
R20310 VSS.n11552 VSS.n11551 0.000501541
R20311 VSS.n11563 VSS.n11562 0.000501541
R20312 VSS.n10626 VSS.n10625 0.000501541
R20313 VSS.n10615 VSS.n10614 0.000501541
R20314 VSS.n10621 VSS.n10620 0.000501541
R20315 VSS.n10609 VSS.n10608 0.000501541
R20316 VSS.n4541 VSS.n4539 0.000501541
R20317 VSS.n3372 VSS.n3370 0.000501541
R20318 VSS.n5397 VSS.n5396 0.000501541
R20319 VSS.n6136 VSS.n6135 0.000501541
R20320 VSS.n6120 VSS.n6119 0.000501541
R20321 VSS.n5954 VSS.n5953 0.000501541
R20322 VSS.n5938 VSS.n5937 0.000501541
R20323 VSS.n5773 VSS.n5772 0.000501541
R20324 VSS.n5757 VSS.n5756 0.000501541
R20325 VSS.n5593 VSS.n5592 0.000501541
R20326 VSS.n5577 VSS.n5576 0.000501541
R20327 VSS.n5413 VSS.n5412 0.000501541
R20328 VSS.n5233 VSS.n5232 0.000501541
R20329 VSS.n5217 VSS.n5216 0.000501541
R20330 VSS.n10111 VSS.n10109 0.000501541
R20331 VSS.n10127 VSS.n10125 0.000501541
R20332 VSS.n11154 VSS.n11152 0.000501541
R20333 VSS.n11170 VSS.n11168 0.000501541
R20334 VSS.n12295 VSS.n12293 0.000501541
R20335 VSS.n12324 VSS.n12323 0.000501541
R20336 VSS.n11559 VSS.n11557 0.000501541
R20337 VSS.n12474 VSS.n12473 0.000501541
R20338 VSS.n12476 VSS.n12470 0.000501541
R20339 VSS.n12181 VSS.n12180 0.000501541
R20340 VSS.n12199 VSS.n12198 0.000501541
R20341 VSS.n14495 VSS.n14494 0.000501541
R20342 VSS.n3317 VSS.n3315 0.000501541
R20343 VSS.n12568 VSS.n12567 0.000501541
R20344 VSS.n3415 VSS.n3414 0.000501541
R20345 VSS.n3584 VSS.n3582 0.000501541
R20346 VSS.n11900 VSS.n11899 0.000501541
R20347 VSS.n12013 VSS.n12012 0.000501541
R20348 VSS.n12029 VSS.n12028 0.000501541
R20349 VSS.n1 VSS.n0 0.000500621
R20350 VSS.n3205 VSS.n3204 0.000500621
R20351 VSS.n3201 VSS.n3200 0.000500621
R20352 VSS.n27 VSS.n26 0.000500621
R20353 VSS.n25 VSS.n24 0.000500621
R20354 VSS.n3198 VSS.n23 0.000500621
R20355 VSS.n3352 VSS.n3351 0.000500621
R20356 VSS.n3348 VSS.n3347 0.000500621
R20357 VSS.n3345 VSS.n3344 0.000500621
R20358 VSS.n11915 VSS.n11914 0.000500621
R20359 VSS.n11911 VSS.n11910 0.000500621
R20360 VSS.n11908 VSS.n11907 0.000500621
R20361 VSS.n11771 VSS.n11770 0.000500621
R20362 VSS.n11767 VSS.n11766 0.000500621
R20363 VSS.n11764 VSS.n11763 0.000500621
R20364 VSS.n3620 VSS.n3619 0.000500621
R20365 VSS.n316 VSS.n315 0.000500621
R20366 VSS.n322 VSS.n316 0.000500621
R20367 VSS.n322 VSS.n321 0.000500621
R20368 VSS.n14402 VSS.n14401 0.000500621
R20369 VSS.n14398 VSS.n14395 0.000500621
R20370 VSS.n296 VSS.n295 0.000500621
R20371 VSS.n294 VSS.n293 0.000500621
R20372 VSS.n300 VSS.n294 0.000500621
R20373 VSS.n300 VSS.n299 0.000500621
R20374 VSS.n4533 VSS.n4532 0.000500621
R20375 VSS.n4530 VSS.n4529 0.000500621
R20376 VSS.n4460 VSS.n4459 0.000500621
R20377 VSS.n4466 VSS.n4460 0.000500621
R20378 VSS.n4466 VSS.n4465 0.000500621
R20379 VSS.n4463 VSS.n4462 0.000500621
R20380 VSS.n4472 VSS.n4470 0.000500621
R20381 VSS.n4477 VSS.n4470 0.000500621
R20382 VSS.n4477 VSS.n4476 0.000500621
R20383 VSS.n4474 VSS.n4473 0.000500621
R20384 VSS.n4484 VSS.n4483 0.000500621
R20385 VSS.n4497 VSS.n4496 0.000500621
R20386 VSS.n4493 VSS.n4492 0.000500621
R20387 VSS.n4499 VSS.n4493 0.000500621
R20388 VSS.n4499 VSS.n4498 0.000500621
R20389 VSS.n4511 VSS.n4510 0.000500621
R20390 VSS.n4507 VSS.n4506 0.000500621
R20391 VSS.n4513 VSS.n4507 0.000500621
R20392 VSS.n4513 VSS.n4512 0.000500621
R20393 VSS.n4520 VSS.n4519 0.000500621
R20394 VSS.n4524 VSS.n4523 0.000500621
R20395 VSS.n1055 VSS.n1054 0.000500621
R20396 VSS.n1061 VSS.n1060 0.000500621
R20397 VSS.n1058 VSS.n1057 0.000500621
R20398 VSS.n13817 VSS.n13816 0.000500621
R20399 VSS.n13823 VSS.n13822 0.000500621
R20400 VSS.n13820 VSS.n13819 0.000500621
R20401 VSS.n13360 VSS.n13359 0.000500621
R20402 VSS.n13357 VSS.n13356 0.000500621
R20403 VSS.n13354 VSS.n13353 0.000500621
R20404 VSS.n13418 VSS.n487 0.000500621
R20405 VSS.n376 VSS.n374 0.000500621
R20406 VSS.n381 VSS.n374 0.000500621
R20407 VSS.n381 VSS.n380 0.000500621
R20408 VSS.n14388 VSS.n14385 0.000500621
R20409 VSS.n14385 VSS.n383 0.000500621
R20410 VSS.n14388 VSS.n14387 0.000500621
R20411 VSS.n378 VSS.n377 0.000500621
R20412 VSS.n238 VSS.n237 0.000500621
R20413 VSS.n235 VSS.n231 0.000500621
R20414 VSS.n120 VSS.n115 0.000500621
R20415 VSS.n119 VSS.n114 0.000500621
R20416 VSS.n120 VSS.n119 0.000500621
R20417 VSS.n32 VSS.n31 0.000500621
R20418 VSS.n30 VSS.n29 0.000500621
R20419 VSS.n36 VSS.n29 0.000500621
R20420 VSS.n36 VSS.n35 0.000500621
R20421 VSS.n175 VSS.n174 0.000500621
R20422 VSS.n173 VSS.n172 0.000500621
R20423 VSS.n179 VSS.n172 0.000500621
R20424 VSS.n179 VSS.n178 0.000500621
R20425 VSS.n14451 VSS.n14449 0.000500621
R20426 VSS.n14449 VSS.n14448 0.000500621
R20427 VSS.n14451 VSS.n14450 0.000500621
R20428 VSS.n331 VSS.n327 0.000500621
R20429 VSS.n331 VSS.n330 0.000500621
R20430 VSS.n327 VSS.n326 0.000500621
R20431 VSS.n202 VSS.n201 0.000500621
R20432 VSS.n208 VSS.n202 0.000500621
R20433 VSS.n208 VSS.n207 0.000500621
R20434 VSS.n218 VSS.n213 0.000500621
R20435 VSS.n218 VSS.n217 0.000500621
R20436 VSS.n213 VSS.n212 0.000500621
R20437 VSS.n313 VSS.n312 0.000500621
R20438 VSS.n14438 VSS.n313 0.000500621
R20439 VSS.n14439 VSS.n14438 0.000500621
R20440 VSS.n385 VSS.n384 0.000500621
R20441 VSS.n391 VSS.n385 0.000500621
R20442 VSS.n391 VSS.n390 0.000500621
R20443 VSS.n395 VSS.n394 0.000500621
R20444 VSS.n401 VSS.n395 0.000500621
R20445 VSS.n401 VSS.n400 0.000500621
R20446 VSS.n1577 VSS.n1576 0.000500621
R20447 VSS.n1583 VSS.n1582 0.000500621
R20448 VSS.n1580 VSS.n1579 0.000500621
R20449 VSS.n454 VSS.n453 0.000500621
R20450 VSS.n471 VSS.n470 0.000500621
R20451 VSS.n452 VSS.n451 0.000500621
R20452 VSS.n1311 VSS.n1310 0.000500621
R20453 VSS.n1308 VSS.n1307 0.000500621
R20454 VSS.n1305 VSS.n1304 0.000500621
R20455 VSS.n435 VSS.n434 0.000500621
R20456 VSS.n441 VSS.n435 0.000500621
R20457 VSS.n441 VSS.n440 0.000500621
R20458 VSS.n431 VSS.n426 0.000500621
R20459 VSS.n431 VSS.n430 0.000500621
R20460 VSS.n426 VSS.n425 0.000500621
R20461 VSS.n14431 VSS.n14429 0.000500621
R20462 VSS.n14429 VSS.n14428 0.000500621
R20463 VSS.n14432 VSS.n14431 0.000500621
R20464 VSS.n14411 VSS.n14409 0.000500621
R20465 VSS.n14412 VSS.n14405 0.000500621
R20466 VSS.n14412 VSS.n14411 0.000500621
R20467 VSS.n222 VSS.n221 0.000500621
R20468 VSS.n228 VSS.n222 0.000500621
R20469 VSS.n228 VSS.n227 0.000500621
R20470 VSS.n86 VSS.n81 0.000500621
R20471 VSS.n87 VSS.n86 0.000500621
R20472 VSS.n56 VSS.n53 0.000500621
R20473 VSS.n59 VSS.n58 0.000500621
R20474 VSS.n257 VSS.n251 0.000500621
R20475 VSS.n257 VSS.n256 0.000500621
R20476 VSS.n247 VSS.n241 0.000500621
R20477 VSS.n247 VSS.n246 0.000500621
R20478 VSS.n14422 VSS.n14416 0.000500621
R20479 VSS.n14422 VSS.n14421 0.000500621
R20480 VSS.n14421 VSS.n14420 0.000500621
R20481 VSS.n411 VSS.n406 0.000500621
R20482 VSS.n411 VSS.n410 0.000500621
R20483 VSS.n406 VSS.n405 0.000500621
R20484 VSS.n421 VSS.n416 0.000500621
R20485 VSS.n421 VSS.n420 0.000500621
R20486 VSS.n416 VSS.n415 0.000500621
R20487 VSS.n14347 VSS.n14346 0.000500621
R20488 VSS.n14344 VSS.n14343 0.000500621
R20489 VSS.n14341 VSS.n14340 0.000500621
R20490 VSS.n14378 VSS.n14377 0.000500621
R20491 VSS.n498 VSS.n497 0.000500621
R20492 VSS.n343 VSS.n338 0.000500621
R20493 VSS.n337 VSS.n336 0.000500621
R20494 VSS.n343 VSS.n337 0.000500621
R20495 VSS.n342 VSS.n341 0.000500621
R20496 VSS.n270 VSS.n265 0.000500621
R20497 VSS.n264 VSS.n263 0.000500621
R20498 VSS.n270 VSS.n264 0.000500621
R20499 VSS.n269 VSS.n268 0.000500621
R20500 VSS.n158 VSS.n153 0.000500621
R20501 VSS.n152 VSS.n151 0.000500621
R20502 VSS.n158 VSS.n152 0.000500621
R20503 VSS.n157 VSS.n156 0.000500621
R20504 VSS.n97 VSS.n92 0.000500621
R20505 VSS.n91 VSS.n90 0.000500621
R20506 VSS.n97 VSS.n91 0.000500621
R20507 VSS.n96 VSS.n95 0.000500621
R20508 VSS.n11546 VSS.n11545 0.000500621
R20509 VSS.n11542 VSS.n11541 0.000500621
R20510 VSS.n11539 VSS.n11538 0.000500621
R20511 VSS.n75 VSS.n70 0.000500621
R20512 VSS.n71 VSS.n69 0.000500621
R20513 VSS.n11795 VSS.n11794 0.000500621
R20514 VSS.n11792 VSS.n11784 0.000500621
R20515 VSS.n11790 VSS.n11789 0.000500621
R20516 VSS.n103 VSS.n102 0.000500621
R20517 VSS.n108 VSS.n107 0.000500621
R20518 VSS.n3430 VSS.n3429 0.000500621
R20519 VSS.n3426 VSS.n3425 0.000500621
R20520 VSS.n3423 VSS.n3422 0.000500621
R20521 VSS.n133 VSS.n128 0.000500621
R20522 VSS.n134 VSS.n133 0.000500621
R20523 VSS.n144 VSS.n139 0.000500621
R20524 VSS.n143 VSS.n142 0.000500621
R20525 VSS.n144 VSS.n143 0.000500621
R20526 VSS.n318 VSS.n317 0.00050031
R20527 VSS.n14415 VSS.n261 0.00050031
R20528 VSS.n14397 VSS.n14396 0.00050031
R20529 VSS.n14400 VSS.n279 0.00050031
R20530 VSS.n404 VSS.n334 0.00050031
R20531 VSS.n389 VSS.n352 0.00050031
R20532 VSS.n1056 VSS.n444 0.00050031
R20533 VSS.n13818 VSS.n491 0.00050031
R20534 VSS.n13355 VSS.n483 0.00050031
R20535 VSS.n14391 VSS.n14390 0.00050031
R20536 VSS.n14386 VSS.n368 0.00050031
R20537 VSS.n255 VSS.n149 0.00050031
R20538 VSS.n233 VSS.n232 0.00050031
R20539 VSS.n234 VSS.n167 0.00050031
R20540 VSS.n123 VSS.n122 0.00050031
R20541 VSS.n14453 VSS.n14452 0.00050031
R20542 VSS.n199 VSS.n198 0.00050031
R20543 VSS.n329 VSS.n328 0.00050031
R20544 VSS.n314 VSS.n304 0.00050031
R20545 VSS.n325 VSS.n308 0.00050031
R20546 VSS.n206 VSS.n196 0.00050031
R20547 VSS.n204 VSS.n203 0.00050031
R20548 VSS.n215 VSS.n214 0.00050031
R20549 VSS.n14441 VSS.n14440 0.00050031
R20550 VSS.n388 VSS.n387 0.00050031
R20551 VSS.n399 VSS.n364 0.00050031
R20552 VSS.n397 VSS.n396 0.00050031
R20553 VSS.n1578 VSS.n479 0.00050031
R20554 VSS.n1306 VSS.n477 0.00050031
R20555 VSS.n473 VSS.n472 0.00050031
R20556 VSS.n437 VSS.n436 0.00050031
R20557 VSS.n428 VSS.n427 0.00050031
R20558 VSS.n424 VSS.n362 0.00050031
R20559 VSS.n439 VSS.n358 0.00050031
R20560 VSS.n14426 VSS.n14425 0.00050031
R20561 VSS.n14407 VSS.n14406 0.00050031
R20562 VSS.n14410 VSS.n289 0.00050031
R20563 VSS.n14430 VSS.n285 0.00050031
R20564 VSS.n224 VSS.n223 0.00050031
R20565 VSS.n226 VSS.n186 0.00050031
R20566 VSS.n211 VSS.n190 0.00050031
R20567 VSS.n80 VSS.n79 0.00050031
R20568 VSS.n62 VSS.n61 0.00050031
R20569 VSS.n254 VSS.n253 0.00050031
R20570 VSS.n243 VSS.n242 0.00050031
R20571 VSS.n14419 VSS.n14418 0.00050031
R20572 VSS.n409 VSS.n408 0.00050031
R20573 VSS.n418 VSS.n417 0.00050031
R20574 VSS.n14342 VSS.n500 0.00050031
R20575 VSS.n414 VSS.n347 0.00050031
R20576 VSS.n320 VSS.n274 0.00050031
R20577 VSS.n245 VSS.n164 0.00050031
R20578 VSS.n83 VSS.n82 0.00050031
R20579 VSS.n68 VSS.n67 0.00050031
R20580 VSS.n74 VSS.n73 0.00050031
R20581 VSS.n55 VSS.n54 0.00050031
R20582 VSS.n110 VSS.n109 0.00050031
R20583 VSS.n105 VSS.n104 0.00050031
R20584 VSS.n117 VSS.n116 0.00050031
R20585 VSS.n136 VSS.n135 0.00050031
R20586 VSS.n131 VSS.n130 0.00050031
R20587 VSS.n141 VSS.n49 0.00050031
R20588 VSS.n146 VSS.n145 0.00050031
R20589 VSS.n8514 VSS.n8513 0.000500172
R20590 VSS.n8512 VSS.n8511 0.000500172
R20591 VSS.n9986 VSS.n9985 0.000500172
R20592 VSS.n6211 VSS.n6210 0.000500172
R20593 VSS.n8123 VSS.n8122 0.000500172
R20594 VSS.n9949 VSS.n9948 0.000500172
R20595 VSS.n6241 VSS.n6240 0.000500172
R20596 VSS.n6240 VSS.n6237 0.000500172
R20597 VSS.n9943 VSS.n6238 0.000500172
R20598 VSS.n9944 VSS.n9943 0.000500172
R20599 VSS.n6238 VSS.n6236 0.000500172
R20600 VSS.n9944 VSS.n6236 0.000500172
R20601 VSS.n8835 VSS.n8834 0.000500172
R20602 VSS.n8160 VSS.n8159 0.000500172
R20603 VSS.n8846 VSS.n8011 0.000500172
R20604 VSS.n8846 VSS.n8845 0.000500172
R20605 VSS.n8011 VSS.n8009 0.000500172
R20606 VSS.n8845 VSS.n8009 0.000500172
R20607 VSS.n8840 VSS.n8839 0.000500172
R20608 VSS.n8844 VSS.n8839 0.000500172
R20609 VSS.n9542 VSS.n9541 0.000500172
R20610 VSS.n9541 VSS.n9540 0.000500172
R20611 VSS.n9544 VSS.n7589 0.000500172
R20612 VSS.n9544 VSS.n9543 0.000500172
R20613 VSS.n7591 VSS.n7589 0.000500172
R20614 VSS.n9543 VSS.n7591 0.000500172
R20615 VSS.n9606 VSS.n9604 0.000500172
R20616 VSS.n9606 VSS.n9605 0.000500172
R20617 VSS.n9608 VSS.n9599 0.000500172
R20618 VSS.n8764 VSS.n8762 0.000500172
R20619 VSS.n8764 VSS.n8763 0.000500172
R20620 VSS.n8761 VSS.n8757 0.000500172
R20621 VSS.n8521 VSS.n8519 0.000500172
R20622 VSS.n8521 VSS.n8520 0.000500172
R20623 VSS.n8518 VSS.n8410 0.000500172
R20624 VSS.n8432 VSS.n8414 0.000500172
R20625 VSS.n8431 VSS.n8430 0.000500172
R20626 VSS.n8416 VSS.n8415 0.000500172
R20627 VSS.n8633 VSS.n8632 0.000500172
R20628 VSS.n8627 VSS.n8626 0.000500172
R20629 VSS.n8622 VSS.n8621 0.000500172
R20630 VSS.n8730 VSS.n8729 0.000500172
R20631 VSS.n8710 VSS.n8709 0.000500172
R20632 VSS.n8652 VSS.n8651 0.000500172
R20633 VSS.n9708 VSS.n9707 0.000500172
R20634 VSS.n9702 VSS.n9701 0.000500172
R20635 VSS.n9697 VSS.n9696 0.000500172
R20636 VSS.n7499 VSS.n7498 0.000500172
R20637 VSS.n9117 VSS.n9116 0.000500172
R20638 VSS.n9055 VSS.n9054 0.000500172
R20639 VSS.n9362 VSS.n9361 0.000500172
R20640 VSS.n3969 VSS.n3968 0.000500172
R20641 VSS.n4027 VSS.n4026 0.000500172
R20642 VSS.n10819 VSS.n10818 0.000500172
R20643 VSS.n9770 VSS.n9769 0.000500172
R20644 VSS.n9772 VSS.n9771 0.000500172
R20645 VSS.n9424 VSS.n9423 0.000500172
R20646 VSS.n9426 VSS.n9425 0.000500172
R20647 VSS.n9804 VSS.n9802 0.000500172
R20648 VSS.n9804 VSS.n9803 0.000500172
R20649 VSS.n9801 VSS.n9795 0.000500172
R20650 VSS.n9461 VSS.n9459 0.000500172
R20651 VSS.n9461 VSS.n9460 0.000500172
R20652 VSS.n9458 VSS.n9454 0.000500172
R20653 VSS.n9152 VSS.n9150 0.000500172
R20654 VSS.n9152 VSS.n9151 0.000500172
R20655 VSS.n9149 VSS.n9145 0.000500172
R20656 VSS.n9861 VSS.n9860 0.000500172
R20657 VSS.n9860 VSS.n9859 0.000500172
R20658 VSS.n9862 VSS.n7147 0.000500172
R20659 VSS.n7148 VSS.n7147 0.000500172
R20660 VSS.n9863 VSS.n7148 0.000500172
R20661 VSS.n9863 VSS.n9862 0.000500172
R20662 VSS.n9853 VSS.n9850 0.000500172
R20663 VSS.n9853 VSS.n9852 0.000500172
R20664 VSS.n9849 VSS.n7154 0.000500172
R20665 VSS.n7154 VSS.n7153 0.000500172
R20666 VSS.n9849 VSS.n9848 0.000500172
R20667 VSS.n9848 VSS.n7153 0.000500172
R20668 VSS.n7606 VSS.n7600 0.000500172
R20669 VSS.n7606 VSS.n7605 0.000500172
R20670 VSS.n7608 VSS.n7601 0.000500172
R20671 VSS.n9527 VSS.n7608 0.000500172
R20672 VSS.n7601 VSS.n7599 0.000500172
R20673 VSS.n9527 VSS.n7599 0.000500172
R20674 VSS.n9530 VSS.n7598 0.000500172
R20675 VSS.n9531 VSS.n7598 0.000500172
R20676 VSS.n9536 VSS.n9535 0.000500172
R20677 VSS.n9535 VSS.n7596 0.000500172
R20678 VSS.n9537 VSS.n7596 0.000500172
R20679 VSS.n9537 VSS.n9536 0.000500172
R20680 VSS.n9908 VSS.n9907 0.000500172
R20681 VSS.n9907 VSS.n9906 0.000500172
R20682 VSS.n6266 VSS.n6265 0.000500172
R20683 VSS.n6267 VSS.n6265 0.000500172
R20684 VSS.n9902 VSS.n6267 0.000500172
R20685 VSS.n9902 VSS.n6266 0.000500172
R20686 VSS.n6264 VSS.n6261 0.000500172
R20687 VSS.n9911 VSS.n6264 0.000500172
R20688 VSS.n6262 VSS.n6260 0.000500172
R20689 VSS.n9916 VSS.n6260 0.000500172
R20690 VSS.n9916 VSS.n9915 0.000500172
R20691 VSS.n9915 VSS.n6262 0.000500172
R20692 VSS.n6259 VSS.n6256 0.000500172
R20693 VSS.n9919 VSS.n6259 0.000500172
R20694 VSS.n6257 VSS.n6255 0.000500172
R20695 VSS.n9924 VSS.n6255 0.000500172
R20696 VSS.n9924 VSS.n9923 0.000500172
R20697 VSS.n9923 VSS.n6257 0.000500172
R20698 VSS.n9929 VSS.n6251 0.000500172
R20699 VSS.n9929 VSS.n9928 0.000500172
R20700 VSS.n9931 VSS.n6252 0.000500172
R20701 VSS.n9932 VSS.n9931 0.000500172
R20702 VSS.n6252 VSS.n6250 0.000500172
R20703 VSS.n9932 VSS.n6250 0.000500172
R20704 VSS.n6247 VSS.n6244 0.000500172
R20705 VSS.n6248 VSS.n6247 0.000500172
R20706 VSS.n9937 VSS.n6245 0.000500172
R20707 VSS.n9938 VSS.n9937 0.000500172
R20708 VSS.n6245 VSS.n6243 0.000500172
R20709 VSS.n9938 VSS.n6243 0.000500172
R20710 VSS.n10038 VSS.n10037 0.000500172
R20711 VSS.n10037 VSS.n10036 0.000500172
R20712 VSS.n10039 VSS.n4633 0.000500172
R20713 VSS.n4634 VSS.n4633 0.000500172
R20714 VSS.n10040 VSS.n4634 0.000500172
R20715 VSS.n10040 VSS.n10039 0.000500172
R20716 VSS.n4641 VSS.n4636 0.000500172
R20717 VSS.n4637 VSS.n4636 0.000500172
R20718 VSS.n10028 VSS.n4640 0.000500172
R20719 VSS.n10028 VSS.n10027 0.000500172
R20720 VSS.n10026 VSS.n4640 0.000500172
R20721 VSS.n10027 VSS.n10026 0.000500172
R20722 VSS.n10023 VSS.n4643 0.000500172
R20723 VSS.n10023 VSS.n10022 0.000500172
R20724 VSS.n10019 VSS.n4645 0.000500172
R20725 VSS.n10019 VSS.n10018 0.000500172
R20726 VSS.n10017 VSS.n4645 0.000500172
R20727 VSS.n10018 VSS.n10017 0.000500172
R20728 VSS.n10014 VSS.n4647 0.000500172
R20729 VSS.n10014 VSS.n10013 0.000500172
R20730 VSS.n10010 VSS.n4649 0.000500172
R20731 VSS.n10010 VSS.n10009 0.000500172
R20732 VSS.n10008 VSS.n4649 0.000500172
R20733 VSS.n10009 VSS.n10008 0.000500172
R20734 VSS.n10005 VSS.n4651 0.000500172
R20735 VSS.n10005 VSS.n10004 0.000500172
R20736 VSS.n10001 VSS.n4653 0.000500172
R20737 VSS.n10001 VSS.n10000 0.000500172
R20738 VSS.n9999 VSS.n4653 0.000500172
R20739 VSS.n10000 VSS.n9999 0.000500172
R20740 VSS.n9996 VSS.n4655 0.000500172
R20741 VSS.n9996 VSS.n9995 0.000500172
R20742 VSS.n9992 VSS.n4657 0.000500172
R20743 VSS.n9992 VSS.n9991 0.000500172
R20744 VSS.n9990 VSS.n4657 0.000500172
R20745 VSS.n9991 VSS.n9990 0.000500172
R20746 VSS.n6150 VSS.n4663 0.000500172
R20747 VSS.n6152 VSS.n6151 0.000500172
R20748 VSS.n6100 VSS.n6099 0.000500172
R20749 VSS.n6089 VSS.n6088 0.000500172
R20750 VSS.n6087 VSS.n5970 0.000500172
R20751 VSS.n6087 VSS.n6086 0.000500172
R20752 VSS.n5967 VSS.n4672 0.000500172
R20753 VSS.n5969 VSS.n5968 0.000500172
R20754 VSS.n5918 VSS.n5917 0.000500172
R20755 VSS.n5907 VSS.n5906 0.000500172
R20756 VSS.n5905 VSS.n5789 0.000500172
R20757 VSS.n5905 VSS.n5904 0.000500172
R20758 VSS.n5786 VSS.n4681 0.000500172
R20759 VSS.n5788 VSS.n5787 0.000500172
R20760 VSS.n5726 VSS.n5725 0.000500172
R20761 VSS.n5724 VSS.n5608 0.000500172
R20762 VSS.n5724 VSS.n5723 0.000500172
R20763 VSS.n5607 VSS.n5606 0.000500172
R20764 VSS.n4691 VSS.n4690 0.000500172
R20765 VSS.n5546 VSS.n5545 0.000500172
R20766 VSS.n5544 VSS.n5428 0.000500172
R20767 VSS.n5544 VSS.n5543 0.000500172
R20768 VSS.n5427 VSS.n5426 0.000500172
R20769 VSS.n4702 VSS.n4701 0.000500172
R20770 VSS.n5366 VSS.n5365 0.000500172
R20771 VSS.n5364 VSS.n5248 0.000500172
R20772 VSS.n5364 VSS.n5363 0.000500172
R20773 VSS.n5247 VSS.n5246 0.000500172
R20774 VSS.n4714 VSS.n4713 0.000500172
R20775 VSS.n5186 VSS.n4574 0.000500172
R20776 VSS.n10099 VSS.n10098 0.000500172
R20777 VSS.n10098 VSS.n10097 0.000500172
R20778 VSS.n10100 VSS.n4572 0.000500172
R20779 VSS.n4571 VSS.n4570 0.000500172
R20780 VSS.n10134 VSS.n10133 0.000500172
R20781 VSS.n11188 VSS.n11187 0.000500172
R20782 VSS.n3713 VSS.n3712 0.000500172
R20783 VSS.n11143 VSS.n3714 0.000500172
R20784 VSS.n11142 VSS.n3716 0.000500172
R20785 VSS.n3783 VSS.n3716 0.000500172
R20786 VSS.n11113 VSS.n3821 0.000500172
R20787 VSS.n11116 VSS.n3821 0.000500172
R20788 VSS.n11117 VSS.n11116 0.000500172
R20789 VSS.n11116 VSS.n11115 0.000500172
R20790 VSS.n11121 VSS.n11120 0.000500172
R20791 VSS.n11120 VSS.n11119 0.000500172
R20792 VSS.n11122 VSS.n3815 0.000500172
R20793 VSS.n3816 VSS.n3815 0.000500172
R20794 VSS.n11123 VSS.n3816 0.000500172
R20795 VSS.n11123 VSS.n11122 0.000500172
R20796 VSS.n3844 VSS.n3843 0.000500172
R20797 VSS.n11005 VSS.n3843 0.000500172
R20798 VSS.n11005 VSS.n11004 0.000500172
R20799 VSS.n11006 VSS.n11005 0.000500172
R20800 VSS.n11002 VSS.n10999 0.000500172
R20801 VSS.n11002 VSS.n11001 0.000500172
R20802 VSS.n3849 VSS.n3848 0.000500172
R20803 VSS.n10998 VSS.n3849 0.000500172
R20804 VSS.n10998 VSS.n10997 0.000500172
R20805 VSS.n10997 VSS.n3848 0.000500172
R20806 VSS.n10954 VSS.n3889 0.000500172
R20807 VSS.n10957 VSS.n3889 0.000500172
R20808 VSS.n10958 VSS.n10957 0.000500172
R20809 VSS.n10957 VSS.n10956 0.000500172
R20810 VSS.n10962 VSS.n10961 0.000500172
R20811 VSS.n10961 VSS.n10960 0.000500172
R20812 VSS.n10963 VSS.n3883 0.000500172
R20813 VSS.n3884 VSS.n3883 0.000500172
R20814 VSS.n10964 VSS.n3884 0.000500172
R20815 VSS.n10964 VSS.n10963 0.000500172
R20816 VSS.n10852 VSS.n10850 0.000500172
R20817 VSS.n10854 VSS.n10850 0.000500172
R20818 VSS.n10854 VSS.n10853 0.000500172
R20819 VSS.n10855 VSS.n10854 0.000500172
R20820 VSS.n10848 VSS.n10846 0.000500172
R20821 VSS.n10848 VSS.n10847 0.000500172
R20822 VSS.n10845 VSS.n10844 0.000500172
R20823 VSS.n10786 VSS.n10785 0.000500172
R20824 VSS.n4105 VSS.n4104 0.000500172
R20825 VSS.n10784 VSS.n4106 0.000500172
R20826 VSS.n4156 VSS.n4155 0.000500172
R20827 VSS.n4441 VSS.n4440 0.000500172
R20828 VSS.n4440 VSS.n4439 0.000500172
R20829 VSS.n4440 VSS.n4156 0.000500172
R20830 VSS.n4358 VSS.n4357 0.000500172
R20831 VSS.n4275 VSS.n4274 0.000500172
R20832 VSS.n4327 VSS.n4260 0.000500172
R20833 VSS.n4329 VSS.n4328 0.000500172
R20834 VSS.n4226 VSS.n4206 0.000500172
R20835 VSS.n4354 VSS.n4353 0.000500172
R20836 VSS.n4353 VSS.n4206 0.000500172
R20837 VSS.n4353 VSS.n4352 0.000500172
R20838 VSS.n4436 VSS.n4435 0.000500172
R20839 VSS.n4413 VSS.n4160 0.000500172
R20840 VSS.n10746 VSS.n10745 0.000500172
R20841 VSS.n10714 VSS.n10713 0.000500172
R20842 VSS.n10652 VSS.n10651 0.000500172
R20843 VSS.n10712 VSS.n10711 0.000500172
R20844 VSS.n14241 VSS.n14240 0.000500172
R20845 VSS.n14239 VSS.n14237 0.000500172
R20846 VSS.n14247 VSS.n14246 0.000500172
R20847 VSS.n14246 VSS.n14245 0.000500172
R20848 VSS.n14249 VSS.n14248 0.000500172
R20849 VSS.n12423 VSS.n12422 0.000500172
R20850 VSS.n12430 VSS.n12429 0.000500172
R20851 VSS.n13067 VSS.n13066 0.000500172
R20852 VSS.n13062 VSS.n13061 0.000500172
R20853 VSS.n13147 VSS.n1903 0.000500172
R20854 VSS.n13147 VSS.n13146 0.000500172
R20855 VSS.n13144 VSS.n1907 0.000500172
R20856 VSS.n1907 VSS.n1906 0.000500172
R20857 VSS.n13143 VSS.n1906 0.000500172
R20858 VSS.n13144 VSS.n13143 0.000500172
R20859 VSS.n2423 VSS.n2422 0.000500172
R20860 VSS.n2428 VSS.n2427 0.000500172
R20861 VSS.n14150 VSS.n609 0.000500172
R20862 VSS.n609 VSS.n607 0.000500172
R20863 VSS.n14151 VSS.n607 0.000500172
R20864 VSS.n14151 VSS.n14150 0.000500172
R20865 VSS.n613 VSS.n612 0.000500172
R20866 VSS.n14149 VSS.n612 0.000500172
R20867 VSS.n14141 VSS.n615 0.000500172
R20868 VSS.n14141 VSS.n14140 0.000500172
R20869 VSS.n14143 VSS.n616 0.000500172
R20870 VSS.n14144 VSS.n14143 0.000500172
R20871 VSS.n616 VSS.n614 0.000500172
R20872 VSS.n14144 VSS.n614 0.000500172
R20873 VSS.n1364 VSS.n1362 0.000500172
R20874 VSS.n1364 VSS.n1363 0.000500172
R20875 VSS.n1361 VSS.n1355 0.000500172
R20876 VSS.n1123 VSS.n1121 0.000500172
R20877 VSS.n1123 VSS.n1122 0.000500172
R20878 VSS.n1120 VSS.n1116 0.000500172
R20879 VSS.n14360 VSS.n14359 0.000500172
R20880 VSS.n14362 VSS.n14361 0.000500172
R20881 VSS.n1074 VSS.n1073 0.000500172
R20882 VSS.n1076 VSS.n1075 0.000500172
R20883 VSS.n1324 VSS.n1323 0.000500172
R20884 VSS.n1326 VSS.n1325 0.000500172
R20885 VSS.n710 VSS.n709 0.000500172
R20886 VSS.n463 VSS.n462 0.000500172
R20887 VSS.n770 VSS.n769 0.000500172
R20888 VSS.n13371 VSS.n13370 0.000500172
R20889 VSS.n13373 VSS.n13372 0.000500172
R20890 VSS.n13836 VSS.n13835 0.000500172
R20891 VSS.n13838 VSS.n13837 0.000500172
R20892 VSS.n1596 VSS.n1595 0.000500172
R20893 VSS.n1598 VSS.n1597 0.000500172
R20894 VSS.n13872 VSS.n13870 0.000500172
R20895 VSS.n13872 VSS.n13871 0.000500172
R20896 VSS.n13869 VSS.n13863 0.000500172
R20897 VSS.n1631 VSS.n1630 0.000500172
R20898 VSS.n1630 VSS.n1629 0.000500172
R20899 VSS.n1632 VSS.n1625 0.000500172
R20900 VSS.n1636 VSS.n1625 0.000500172
R20901 VSS.n1636 VSS.n1635 0.000500172
R20902 VSS.n805 VSS.n803 0.000500172
R20903 VSS.n805 VSS.n804 0.000500172
R20904 VSS.n802 VSS.n798 0.000500172
R20905 VSS.n14041 VSS.n14040 0.000500172
R20906 VSS.n14040 VSS.n14039 0.000500172
R20907 VSS.n1703 VSS.n1702 0.000500172
R20908 VSS.n1704 VSS.n1702 0.000500172
R20909 VSS.n13912 VSS.n1704 0.000500172
R20910 VSS.n13912 VSS.n1703 0.000500172
R20911 VSS.n14052 VSS.n1701 0.000500172
R20912 VSS.n14044 VSS.n1701 0.000500172
R20913 VSS.n1700 VSS.n1699 0.000500172
R20914 VSS.n1699 VSS.n1697 0.000500172
R20915 VSS.n14056 VSS.n1700 0.000500172
R20916 VSS.n14056 VSS.n1697 0.000500172
R20917 VSS.n14045 VSS.n623 0.000500172
R20918 VSS.n14046 VSS.n14045 0.000500172
R20919 VSS.n625 VSS.n624 0.000500172
R20920 VSS.n14126 VSS.n625 0.000500172
R20921 VSS.n624 VSS.n622 0.000500172
R20922 VSS.n14126 VSS.n622 0.000500172
R20923 VSS.n14129 VSS.n621 0.000500172
R20924 VSS.n14130 VSS.n621 0.000500172
R20925 VSS.n14135 VSS.n14134 0.000500172
R20926 VSS.n14134 VSS.n619 0.000500172
R20927 VSS.n14136 VSS.n619 0.000500172
R20928 VSS.n14136 VSS.n14135 0.000500172
R20929 VSS.n12705 VSS.n12704 0.000500172
R20930 VSS.n12704 VSS.n12703 0.000500172
R20931 VSS.n12706 VSS.n12696 0.000500172
R20932 VSS.n12697 VSS.n12696 0.000500172
R20933 VSS.n12707 VSS.n12697 0.000500172
R20934 VSS.n12707 VSS.n12706 0.000500172
R20935 VSS.n13175 VSS.n1885 0.000500172
R20936 VSS.n1887 VSS.n1885 0.000500172
R20937 VSS.n1883 VSS.n1881 0.000500172
R20938 VSS.n1884 VSS.n1883 0.000500172
R20939 VSS.n13179 VSS.n1884 0.000500172
R20940 VSS.n13179 VSS.n1881 0.000500172
R20941 VSS.n1893 VSS.n1888 0.000500172
R20942 VSS.n1889 VSS.n1888 0.000500172
R20943 VSS.n13170 VSS.n1892 0.000500172
R20944 VSS.n13170 VSS.n13169 0.000500172
R20945 VSS.n13168 VSS.n1892 0.000500172
R20946 VSS.n13169 VSS.n13168 0.000500172
R20947 VSS.n13165 VSS.n1895 0.000500172
R20948 VSS.n13165 VSS.n13164 0.000500172
R20949 VSS.n13161 VSS.n1897 0.000500172
R20950 VSS.n13161 VSS.n13160 0.000500172
R20951 VSS.n13159 VSS.n1897 0.000500172
R20952 VSS.n13160 VSS.n13159 0.000500172
R20953 VSS.n13156 VSS.n1899 0.000500172
R20954 VSS.n13156 VSS.n13155 0.000500172
R20955 VSS.n13152 VSS.n1901 0.000500172
R20956 VSS.n13152 VSS.n13151 0.000500172
R20957 VSS.n13150 VSS.n1901 0.000500172
R20958 VSS.n13151 VSS.n13150 0.000500172
R20959 VSS.n12842 VSS.n12841 0.000500172
R20960 VSS.n12841 VSS.n12840 0.000500172
R20961 VSS.n12612 VSS.n2918 0.000500172
R20962 VSS.n12612 VSS.n2919 0.000500172
R20963 VSS.n2918 VSS.n2917 0.000500172
R20964 VSS.n2919 VSS.n2917 0.000500172
R20965 VSS.n12847 VSS.n12846 0.000500172
R20966 VSS.n12846 VSS.n12845 0.000500172
R20967 VSS.n12849 VSS.n2904 0.000500172
R20968 VSS.n12849 VSS.n12848 0.000500172
R20969 VSS.n2906 VSS.n2904 0.000500172
R20970 VSS.n12848 VSS.n2906 0.000500172
R20971 VSS.n2912 VSS.n2738 0.000500172
R20972 VSS.n2912 VSS.n2911 0.000500172
R20973 VSS.n2740 VSS.n2739 0.000500172
R20974 VSS.n12919 VSS.n2740 0.000500172
R20975 VSS.n2739 VSS.n2737 0.000500172
R20976 VSS.n12919 VSS.n2737 0.000500172
R20977 VSS.n12924 VSS.n12923 0.000500172
R20978 VSS.n12923 VSS.n12922 0.000500172
R20979 VSS.n12926 VSS.n2724 0.000500172
R20980 VSS.n12926 VSS.n12925 0.000500172
R20981 VSS.n2726 VSS.n2724 0.000500172
R20982 VSS.n12925 VSS.n2726 0.000500172
R20983 VSS.n2732 VSS.n2557 0.000500172
R20984 VSS.n2732 VSS.n2731 0.000500172
R20985 VSS.n2559 VSS.n2558 0.000500172
R20986 VSS.n12996 VSS.n2559 0.000500172
R20987 VSS.n2558 VSS.n2556 0.000500172
R20988 VSS.n12996 VSS.n2556 0.000500172
R20989 VSS.n12425 VSS.n2553 0.000500172
R20990 VSS.n2554 VSS.n2553 0.000500172
R20991 VSS.n2552 VSS.n2551 0.000500172
R20992 VSS.n2551 VSS.n2549 0.000500172
R20993 VSS.n13001 VSS.n2552 0.000500172
R20994 VSS.n13001 VSS.n2549 0.000500172
R20995 VSS.n12364 VSS.n12363 0.000500172
R20996 VSS.n12462 VSS.n12461 0.000500172
R20997 VSS.n12347 VSS.n12346 0.000500172
R20998 VSS.n12343 VSS.n12342 0.000500172
R20999 VSS.n12342 VSS.n12341 0.000500172
R21000 VSS.n12339 VSS.n11684 0.000500172
R21001 VSS.n11683 VSS.n11682 0.000500172
R21002 VSS.n12267 VSS.n12266 0.000500172
R21003 VSS.n12265 VSS.n12264 0.000500172
R21004 VSS.n12265 VSS.n12208 0.000500172
R21005 VSS.n12206 VSS.n11753 0.000500172
R21006 VSS.n11752 VSS.n11751 0.000500172
R21007 VSS.n12160 VSS.n12159 0.000500172
R21008 VSS.n12158 VSS.n12157 0.000500172
R21009 VSS.n12158 VSS.n12044 0.000500172
R21010 VSS.n12042 VSS.n11782 0.000500172
R21011 VSS.n11781 VSS.n11780 0.000500172
R21012 VSS.n11992 VSS.n11991 0.000500172
R21013 VSS.n11990 VSS.n11989 0.000500172
R21014 VSS.n11990 VSS.n11933 0.000500172
R21015 VSS.n11931 VSS.n11930 0.000500172
R21016 VSS.n11884 VSS.n11883 0.000500172
R21017 VSS.n3564 VSS.n3563 0.000500172
R21018 VSS.n3562 VSS.n3561 0.000500172
R21019 VSS.n3562 VSS.n3448 0.000500172
R21020 VSS.n3446 VSS.n3445 0.000500172
R21021 VSS.n3399 VSS.n3398 0.000500172
R21022 VSS.n3357 VSS.n3116 0.000500172
R21023 VSS.n12585 VSS.n12584 0.000500172
R21024 VSS.n12584 VSS.n12583 0.000500172
R21025 VSS.n12581 VSS.n12580 0.000500172
R21026 VSS.n3173 VSS.n3172 0.000500172
R21027 VSS.n3291 VSS.n3290 0.000500172
R21028 VSS.n12812 VSS.n12811 0.000500172
R21029 VSS.n3191 VSS.n3190 0.000500172
R21030 VSS.n3214 VSS.n3213 0.000500172
R21031 VSS.n3289 VSS.n3188 0.000500172
R21032 VSS.n3289 VSS.n3288 0.000500172
R21033 VSS.n12824 VSS.n2926 0.000500172
R21034 VSS.n12827 VSS.n2926 0.000500172
R21035 VSS.n12828 VSS.n12827 0.000500172
R21036 VSS.n12827 VSS.n12826 0.000500172
R21037 VSS.n12831 VSS.n2925 0.000500172
R21038 VSS.n12830 VSS.n2925 0.000500172
R21039 VSS.n12837 VSS.n2924 0.000500172
R21040 VSS.n12837 VSS.n12836 0.000500172
R21041 VSS.n12836 VSS.n12835 0.000500172
R21042 VSS.n12835 VSS.n2924 0.000500172
R21043 VSS.n1750 VSS.n1749 0.000500172
R21044 VSS.n14001 VSS.n1749 0.000500172
R21045 VSS.n14001 VSS.n14000 0.000500172
R21046 VSS.n14002 VSS.n14001 0.000500172
R21047 VSS.n13998 VSS.n13995 0.000500172
R21048 VSS.n13998 VSS.n13997 0.000500172
R21049 VSS.n1755 VSS.n1754 0.000500172
R21050 VSS.n13994 VSS.n1755 0.000500172
R21051 VSS.n13994 VSS.n13993 0.000500172
R21052 VSS.n13993 VSS.n1754 0.000500172
R21053 VSS.n14023 VSS.n1711 0.000500172
R21054 VSS.n14026 VSS.n1711 0.000500172
R21055 VSS.n14027 VSS.n14026 0.000500172
R21056 VSS.n14026 VSS.n14025 0.000500172
R21057 VSS.n14030 VSS.n1710 0.000500172
R21058 VSS.n14029 VSS.n1710 0.000500172
R21059 VSS.n14036 VSS.n1709 0.000500172
R21060 VSS.n14036 VSS.n14035 0.000500172
R21061 VSS.n14035 VSS.n14034 0.000500172
R21062 VSS.n14034 VSS.n1709 0.000500172
R21063 VSS.n13613 VSS.n13400 0.000500172
R21064 VSS.n13613 VSS.n13612 0.000500172
R21065 VSS.n13612 VSS.n13402 0.000500172
R21066 VSS.n13612 VSS.n13611 0.000500172
R21067 VSS.n13621 VSS.n13619 0.000500172
R21068 VSS.n13621 VSS.n13620 0.000500172
R21069 VSS.n13618 VSS.n13398 0.000500172
R21070 VSS.n13617 VSS.n13398 0.000500172
R21071 VSS.n13428 VSS.n13427 0.000500172
R21072 VSS.n8515 VSS.n8514 0.000500086
R21073 VSS.n8512 VSS.n8490 0.000500086
R21074 VSS.n9987 VSS.n9986 0.000500086
R21075 VSS.n6211 VSS.n4658 0.000500086
R21076 VSS.n8122 VSS.n6235 0.000500086
R21077 VSS.n9948 VSS.n9947 0.000500086
R21078 VSS.n8836 VSS.n8835 0.000500086
R21079 VSS.n8160 VSS.n8012 0.000500086
R21080 VSS.n4274 VSS.n4205 0.000500086
R21081 VSS.n4357 VSS.n4356 0.000500086
R21082 VSS.n4413 VSS.n4157 0.000500086
R21083 VSS.n4437 VSS.n4436 0.000500086
R21084 VSS.n14242 VSS.n14241 0.000500086
R21085 VSS.n14239 VSS.n14238 0.000500086
R21086 VSS.n12424 VSS.n12423 0.000500086
R21087 VSS.n12429 VSS.n12428 0.000500086
R21088 VSS.n13066 VSS.n13065 0.000500086
R21089 VSS.n13063 VSS.n13062 0.000500086
R21090 VSS.n2424 VSS.n2423 0.000500086
R21091 VSS.n2427 VSS.n2426 0.000500086
R21092 VDD VDD 1546.9
R21093 VDD VDD 1544.17
R21094 VDD VDD.n27 896.29
R21095 VDD VDD.n232 896.29
R21096 VDD.n88 VDD 646.457
R21097 VDD.n296 VDD.n295 469.212
R21098 VDD VDD 468.286
R21099 VDD VDD 468.286
R21100 VDD VDD 464.93
R21101 VDD VDD 464.93
R21102 VDD VDD 463.252
R21103 VDD VDD 463.252
R21104 VDD.n233 VDD 459.156
R21105 VDD VDD 459.027
R21106 VDD VDD 458.216
R21107 VDD VDD 458.216
R21108 VDD.n28 VDD 454.192
R21109 VDD.n295 VDD 436.397
R21110 VDD.n86 VDD 279.115
R21111 VDD.n232 VDD 189.665
R21112 VDD.n89 VDD.n88 147.387
R21113 VDD VDD 146.025
R21114 VDD.n87 VDD.n86 141.239
R21115 VDD.n27 VDD.n26 140.989
R21116 VDD.n295 VDD.n294 120.481
R21117 VDD.n86 VDD.n85 116.73
R21118 VDD.n27 VDD.n18 116.73
R21119 VDD.n232 VDD.n226 116.73
R21120 VDD.n88 VDD.n87 61.4756
R21121 VDD.n26 VDD 48.7616
R21122 VDD.n26 VDD 48.6754
R21123 VDD.n87 VDD 42.0359
R21124 VDD.n41 VDD.n23 34.6358
R21125 VDD.n85 VDD.n10 34.6358
R21126 VDD.n35 VDD.n25 34.6358
R21127 VDD.n40 VDD.n24 34.6358
R21128 VDD.n55 VDD.n20 34.6358
R21129 VDD.n56 VDD.n55 34.6358
R21130 VDD.n57 VDD.n18 34.6358
R21131 VDD.n61 VDD.n18 34.6358
R21132 VDD.n62 VDD.n61 34.6358
R21133 VDD.n62 VDD.n17 34.6358
R21134 VDD.n67 VDD.n66 34.6358
R21135 VDD.n68 VDD.n67 34.6358
R21136 VDD.n72 VDD.n15 34.6358
R21137 VDD.n73 VDD.n72 34.6358
R21138 VDD.n74 VDD.n13 34.6358
R21139 VDD.n85 VDD.n11 34.6358
R21140 VDD.n268 VDD.n226 34.6358
R21141 VDD.n269 VDD.n268 34.6358
R21142 VDD.n240 VDD.n231 34.6358
R21143 VDD.n245 VDD.n230 34.6358
R21144 VDD.n246 VDD.n229 34.6358
R21145 VDD.n264 VDD.n226 34.6358
R21146 VDD.n46 VDD.n45 28.9887
R21147 VDD.n251 VDD.n250 28.9887
R21148 VDD.n139 VDD.t0 27.8779
R21149 VDD.n146 VDD.t2 27.8779
R21150 VDD.n153 VDD.t4 27.8779
R21151 VDD.t4 VDD.n152 27.8777
R21152 VDD.t2 VDD.n145 27.8777
R21153 VDD.t0 VDD.n138 27.8777
R21154 VDD.n41 VDD 27.8593
R21155 VDD.n246 VDD 27.8593
R21156 VDD.n79 VDD.n78 25.977
R21157 VDD.n80 VDD.n79 24.4711
R21158 VDD.n290 VDD.n289 24.4711
R21159 VDD.n89 VDD.n10 23.7181
R21160 VDD.n30 VDD.n28 23.7181
R21161 VDD.n51 VDD.n20 23.7181
R21162 VDD.n78 VDD.n13 23.7181
R21163 VDD.n80 VDD.n11 23.7181
R21164 VDD.n289 VDD.n288 23.7181
R21165 VDD.n235 VDD.n233 23.7181
R21166 VDD.n51 VDD 20.7064
R21167 VDD.n256 VDD 20.7064
R21168 VDD.n31 VDD.n30 18.824
R21169 VDD.n36 VDD.n35 18.824
R21170 VDD.n236 VDD.n235 18.824
R21171 VDD.n241 VDD.n240 18.824
R21172 VDD.n45 VDD.n23 15.4358
R21173 VDD.n250 VDD.n229 15.4358
R21174 VDD.n31 VDD.n25 13.9299
R21175 VDD.n36 VDD.n24 13.9299
R21176 VDD.n66 VDD.n17 13.9299
R21177 VDD.n68 VDD.n15 13.9299
R21178 VDD.n236 VDD.n231 13.9299
R21179 VDD.n241 VDD.n230 13.9299
R21180 VDD.n294 VDD.n224 12.8005
R21181 VDD.n202 VDD.n201 10.416
R21182 VDD.n47 VDD.n46 9.78874
R21183 VDD.n57 VDD.n56 9.78874
R21184 VDD.n252 VDD.n251 9.78874
R21185 VDD.n47 VDD.n21 8.28285
R21186 VDD.n252 VDD.n227 8.28285
R21187 VDD VDD.n40 6.77697
R21188 VDD VDD.n50 6.77697
R21189 VDD VDD.n245 6.77697
R21190 VDD VDD.n255 6.77697
R21191 VDD.n74 VDD.n73 5.64756
R21192 VDD.n50 VDD.n21 5.64756
R21193 VDD.n255 VDD.n227 5.64756
R21194 VDD VDD.n28 4.68175
R21195 VDD VDD.n233 4.68175
R21196 VDD.n32 VDD.n31 4.6505
R21197 VDD.n45 VDD.n44 4.6505
R21198 VDD.n48 VDD.n47 4.6505
R21199 VDD.n52 VDD.n51 4.6505
R21200 VDD.n64 VDD.n17 4.6505
R21201 VDD.n78 VDD.n77 4.6505
R21202 VDD.n81 VDD.n80 4.6505
R21203 VDD.n85 VDD.n84 4.6505
R21204 VDD.n30 VDD.n29 4.6505
R21205 VDD.n33 VDD.n25 4.6505
R21206 VDD.n35 VDD.n34 4.6505
R21207 VDD.n37 VDD.n36 4.6505
R21208 VDD.n38 VDD.n24 4.6505
R21209 VDD.n40 VDD.n39 4.6505
R21210 VDD.n42 VDD.n41 4.6505
R21211 VDD.n43 VDD.n23 4.6505
R21212 VDD.n46 VDD.n22 4.6505
R21213 VDD.n50 VDD.n49 4.6505
R21214 VDD.n53 VDD.n20 4.6505
R21215 VDD.n55 VDD.n54 4.6505
R21216 VDD.n56 VDD.n19 4.6505
R21217 VDD.n58 VDD.n57 4.6505
R21218 VDD.n59 VDD.n18 4.6505
R21219 VDD.n61 VDD.n60 4.6505
R21220 VDD.n63 VDD.n62 4.6505
R21221 VDD.n66 VDD.n65 4.6505
R21222 VDD.n67 VDD.n16 4.6505
R21223 VDD.n69 VDD.n68 4.6505
R21224 VDD.n70 VDD.n15 4.6505
R21225 VDD.n72 VDD.n71 4.6505
R21226 VDD.n73 VDD.n14 4.6505
R21227 VDD.n75 VDD.n74 4.6505
R21228 VDD.n76 VDD.n13 4.6505
R21229 VDD.n79 VDD.n12 4.6505
R21230 VDD.n82 VDD.n11 4.6505
R21231 VDD.n83 VDD.n10 4.6505
R21232 VDD.n90 VDD.n89 4.6505
R21233 VDD.n235 VDD.n234 4.6505
R21234 VDD.n237 VDD.n236 4.6505
R21235 VDD.n238 VDD.n231 4.6505
R21236 VDD.n240 VDD.n239 4.6505
R21237 VDD.n242 VDD.n241 4.6505
R21238 VDD.n243 VDD.n230 4.6505
R21239 VDD.n245 VDD.n244 4.6505
R21240 VDD.n247 VDD.n246 4.6505
R21241 VDD.n248 VDD.n229 4.6505
R21242 VDD.n250 VDD.n249 4.6505
R21243 VDD.n251 VDD.n228 4.6505
R21244 VDD.n253 VDD.n252 4.6505
R21245 VDD.n255 VDD.n254 4.6505
R21246 VDD.n257 VDD.n256 4.6505
R21247 VDD.n259 VDD.n258 4.6505
R21248 VDD.n261 VDD.n260 4.6505
R21249 VDD.n263 VDD.n262 4.6505
R21250 VDD.n265 VDD.n264 4.6505
R21251 VDD.n266 VDD.n226 4.6505
R21252 VDD.n268 VDD.n267 4.6505
R21253 VDD.n270 VDD.n269 4.6505
R21254 VDD.n272 VDD.n271 4.6505
R21255 VDD.n274 VDD.n273 4.6505
R21256 VDD.n276 VDD.n275 4.6505
R21257 VDD.n278 VDD.n277 4.6505
R21258 VDD.n280 VDD.n279 4.6505
R21259 VDD.n282 VDD.n281 4.6505
R21260 VDD.n284 VDD.n283 4.6505
R21261 VDD.n286 VDD.n285 4.6505
R21262 VDD.n288 VDD.n287 4.6505
R21263 VDD.n289 VDD.n225 4.6505
R21264 VDD.n291 VDD.n290 4.6505
R21265 VDD.n292 VDD.n224 4.6505
R21266 VDD.n294 VDD.n293 4.6505
R21267 VDD.n9 VDD 4.39723
R21268 VDD.n111 VDD 4.05613
R21269 VDD.n21 VDD 3.55008
R21270 VDD.n227 VDD 3.55008
R21271 VDD.n217 VDD.n98 3.4105
R21272 VDD.n220 VDD.n98 3.4105
R21273 VDD.n216 VDD.n99 3.4105
R21274 VDD.n97 VDD.n8 3.4105
R21275 VDD.n9 VDD.n8 3.4105
R21276 VDD.n9 VDD.n5 3.4105
R21277 VDD.n97 VDD.n5 3.4105
R21278 VDD.n97 VDD.n96 3.4105
R21279 VDD.n96 VDD.n9 3.4105
R21280 VDD.n219 VDD.n217 3.4105
R21281 VDD.n221 VDD.n220 3.4105
R21282 VDD.n220 VDD.n219 3.4105
R21283 VDD.n136 VDD 2.29217
R21284 VDD.n155 VDD 2.29217
R21285 VDD.n103 VDD.n102 1.7055
R21286 VDD.n207 VDD.n203 1.7055
R21287 VDD.n137 VDD.n133 1.57342
R21288 VDD.n140 VDD.n133 1.57342
R21289 VDD.n144 VDD.n130 1.57342
R21290 VDD.n147 VDD.n130 1.57342
R21291 VDD.n151 VDD.n127 1.57342
R21292 VDD.n154 VDD.n127 1.57342
R21293 VDD VDD.n223 1.4367
R21294 VDD.n125 VDD.n124 1.38439
R21295 VDD.n91 VDD 1.34425
R21296 VDD.n132 VDD 0.828181
R21297 VDD.n129 VDD 0.828181
R21298 VDD.n126 VDD 0.828181
R21299 VDD.n132 VDD 0.827501
R21300 VDD.n129 VDD 0.827501
R21301 VDD.n126 VDD 0.827501
R21302 VDD.n198 VDD.n188 0.579775
R21303 VDD.n155 VDD.n124 0.5505
R21304 VDD VDD.n131 0.3755
R21305 VDD VDD.n128 0.3755
R21306 VDD.n178 VDD.n177 0.355402
R21307 VDD.n134 VDD 0.234474
R21308 VDD.n133 VDD.n132 0.232147
R21309 VDD.n130 VDD.n129 0.232147
R21310 VDD.n127 VDD.n126 0.232147
R21311 VDD.n135 VDD.n134 0.222956
R21312 VDD VDD.n296 0.207531
R21313 VDD.n142 VDD.n131 0.167065
R21314 VDD.n149 VDD.n128 0.167065
R21315 VDD.n92 VDD.n91 0.149442
R21316 VDD.n223 VDD.n0 0.14944
R21317 VDD.n94 VDD.n93 0.148938
R21318 VDD.n222 VDD.n1 0.148938
R21319 VDD.n296 VDD 0.129576
R21320 VDD.n33 VDD.n32 0.120292
R21321 VDD.n38 VDD.n37 0.120292
R21322 VDD.n43 VDD.n42 0.120292
R21323 VDD.n44 VDD.n43 0.120292
R21324 VDD.n48 VDD.n22 0.120292
R21325 VDD.n53 VDD.n52 0.120292
R21326 VDD.n54 VDD.n53 0.120292
R21327 VDD.n54 VDD.n19 0.120292
R21328 VDD.n58 VDD.n19 0.120292
R21329 VDD.n64 VDD.n63 0.120292
R21330 VDD.n65 VDD.n64 0.120292
R21331 VDD.n65 VDD.n16 0.120292
R21332 VDD.n69 VDD.n16 0.120292
R21333 VDD.n70 VDD.n69 0.120292
R21334 VDD.n71 VDD.n70 0.120292
R21335 VDD.n71 VDD.n14 0.120292
R21336 VDD.n75 VDD.n14 0.120292
R21337 VDD.n76 VDD.n75 0.120292
R21338 VDD.n77 VDD.n12 0.120292
R21339 VDD.n81 VDD.n12 0.120292
R21340 VDD.n84 VDD.n82 0.120292
R21341 VDD.n238 VDD.n237 0.120292
R21342 VDD.n243 VDD.n242 0.120292
R21343 VDD.n248 VDD.n247 0.120292
R21344 VDD.n249 VDD.n248 0.120292
R21345 VDD.n253 VDD.n228 0.120292
R21346 VDD.n259 VDD.n257 0.120292
R21347 VDD.n261 VDD.n259 0.120292
R21348 VDD.n263 VDD.n261 0.120292
R21349 VDD.n265 VDD.n263 0.120292
R21350 VDD.n272 VDD.n270 0.120292
R21351 VDD.n274 VDD.n272 0.120292
R21352 VDD.n276 VDD.n274 0.120292
R21353 VDD.n278 VDD.n276 0.120292
R21354 VDD.n280 VDD.n278 0.120292
R21355 VDD.n282 VDD.n280 0.120292
R21356 VDD.n284 VDD.n282 0.120292
R21357 VDD.n286 VDD.n284 0.120292
R21358 VDD.n287 VDD.n286 0.120292
R21359 VDD.n292 VDD.n291 0.120292
R21360 VDD.n217 VDD.n216 0.119058
R21361 VDD.n220 VDD.n97 0.119058
R21362 VDD.n131 VDD 0.117487
R21363 VDD.n128 VDD 0.117487
R21364 VDD.n135 VDD 0.117222
R21365 VDD.n156 VDD 0.105191
R21366 VDD.t1 VDD 0.104171
R21367 VDD.n291 VDD 0.0994583
R21368 VDD.n32 VDD 0.0981562
R21369 VDD.n37 VDD 0.0981562
R21370 VDD.n237 VDD 0.0981562
R21371 VDD.n242 VDD 0.0981562
R21372 VDD.n42 VDD 0.0968542
R21373 VDD.n52 VDD 0.0968542
R21374 VDD.n247 VDD 0.0968542
R21375 VDD.n257 VDD 0.0968542
R21376 VDD.n141 VDD.n140 0.0914585
R21377 VDD.n144 VDD.n143 0.0914585
R21378 VDD.n148 VDD.n147 0.0914585
R21379 VDD.n151 VDD.n150 0.0914585
R21380 VDD.n153 VDD.n125 0.0888625
R21381 VDD.n157 VDD.n156 0.0878059
R21382 VDD.t5 VDD 0.0806706
R21383 VDD.t3 VDD 0.0806706
R21384 VDD.t1 VDD 0.0806706
R21385 VDD.t5 VDD 0.0805539
R21386 VDD.t3 VDD 0.0805539
R21387 VDD.t1 VDD 0.0805539
R21388 VDD.n167 VDD.n157 0.0799118
R21389 VDD.n92 VDD.n8 0.075973
R21390 VDD.n98 VDD.n0 0.0752244
R21391 VDD.n186 VDD.n185 0.0617864
R21392 VDD.n194 VDD.n193 0.0617864
R21393 VDD.n211 VDD.n210 0.0617766
R21394 VDD.n210 VDD.n202 0.0617745
R21395 VDD.n175 VDD.n118 0.0612843
R21396 VDD.n171 VDD.n122 0.0612843
R21397 VDD.n115 VDD.n114 0.0612843
R21398 VDD.n123 VDD.n116 0.0612843
R21399 VDD.n170 VDD.n169 0.0612843
R21400 VDD.n184 VDD.n113 0.0612843
R21401 VDD.n183 VDD.n181 0.0612843
R21402 VDD.n192 VDD.n190 0.0612843
R21403 VDD.n196 VDD.n105 0.0612843
R21404 VDD.n195 VDD.n104 0.0612843
R21405 VDD.n29 VDD 0.0603958
R21406 VDD VDD.n33 0.0603958
R21407 VDD.n34 VDD 0.0603958
R21408 VDD VDD.n38 0.0603958
R21409 VDD.n39 VDD 0.0603958
R21410 VDD VDD.n22 0.0603958
R21411 VDD VDD.n48 0.0603958
R21412 VDD.n49 VDD 0.0603958
R21413 VDD VDD.n58 0.0603958
R21414 VDD.n59 VDD 0.0603958
R21415 VDD.n60 VDD 0.0603958
R21416 VDD.n63 VDD 0.0603958
R21417 VDD.n77 VDD 0.0603958
R21418 VDD.n82 VDD 0.0603958
R21419 VDD VDD.n83 0.0603958
R21420 VDD.n90 VDD 0.0603958
R21421 VDD.n234 VDD 0.0603958
R21422 VDD VDD.n238 0.0603958
R21423 VDD.n239 VDD 0.0603958
R21424 VDD VDD.n243 0.0603958
R21425 VDD.n244 VDD 0.0603958
R21426 VDD VDD.n228 0.0603958
R21427 VDD VDD.n253 0.0603958
R21428 VDD.n254 VDD 0.0603958
R21429 VDD VDD.n265 0.0603958
R21430 VDD.n266 VDD 0.0603958
R21431 VDD.n267 VDD 0.0603958
R21432 VDD.n270 VDD 0.0603958
R21433 VDD VDD.n225 0.0603958
R21434 VDD VDD.n292 0.0603958
R21435 VDD.n293 VDD 0.0603958
R21436 VDD.n95 VDD.n5 0.0585072
R21437 VDD.n221 VDD.n3 0.0573205
R21438 VDD.n165 VDD.n160 0.0497515
R21439 VDD.n137 VDD.n136 0.049413
R21440 VDD.n155 VDD.n154 0.049413
R21441 VDD.n205 VDD.n203 0.0484911
R21442 VDD.n164 VDD 0.0482381
R21443 VDD.n204 VDD.n103 0.047933
R21444 VDD.n138 VDD.n134 0.0466957
R21445 VDD.n139 VDD.n131 0.0466957
R21446 VDD.n145 VDD.n131 0.0466957
R21447 VDD.n146 VDD.n128 0.0466957
R21448 VDD.n152 VDD.n128 0.0466957
R21449 VDD.n161 VDD 0.0430763
R21450 VDD.n162 VDD 0.0430763
R21451 VDD.n165 VDD.n164 0.0424716
R21452 VDD.n156 VDD.n155 0.0394617
R21453 VDD.n164 VDD.n163 0.0390868
R21454 VDD VDD.n59 0.0382604
R21455 VDD VDD.n266 0.0382604
R21456 VDD.n168 VDD.n124 0.0357941
R21457 VDD.n84 VDD 0.03175
R21458 VDD VDD.n90 0.03175
R21459 VDD.n293 VDD 0.03175
R21460 VDD.n296 VDD 0.03175
R21461 VDD.n166 VDD.n165 0.0294373
R21462 VDD.n157 VDD.n125 0.0287781
R21463 VDD.n44 VDD 0.0278438
R21464 VDD.n60 VDD 0.0278438
R21465 VDD VDD.n76 0.0278438
R21466 VDD.n249 VDD 0.0278438
R21467 VDD.n267 VDD 0.0278438
R21468 VDD.n287 VDD 0.0278438
R21469 VDD.n136 VDD.n135 0.0270767
R21470 VDD.n161 VDD.t1 0.024
R21471 VDD.n162 VDD.t3 0.024
R21472 VDD.t3 VDD.n161 0.024
R21473 VDD.n163 VDD.t5 0.024
R21474 VDD.t5 VDD.n162 0.024
R21475 VDD.n39 VDD 0.0239375
R21476 VDD.n49 VDD 0.0239375
R21477 VDD VDD.n81 0.0239375
R21478 VDD.n244 VDD 0.0239375
R21479 VDD.n254 VDD 0.0239375
R21480 VDD.n119 VDD.n117 0.0238632
R21481 VDD.n174 VDD.n173 0.0233549
R21482 VDD.n172 VDD.n121 0.0233549
R21483 VDD.n158 VDD.n120 0.0233549
R21484 VDD.n112 VDD.n109 0.0233549
R21485 VDD.n182 VDD.n110 0.0233549
R21486 VDD.n189 VDD.n108 0.0233549
R21487 VDD.n197 VDD.n106 0.0233549
R21488 VDD.n29 VDD 0.0226354
R21489 VDD.n34 VDD 0.0226354
R21490 VDD.n83 VDD 0.0226354
R21491 VDD.n234 VDD 0.0226354
R21492 VDD.n239 VDD 0.0226354
R21493 VDD.n209 VDD.n203 0.0222634
R21494 VDD.n211 VDD.n103 0.0222634
R21495 VDD.n225 VDD 0.0213333
R21496 VDD.n143 VDD 0.0209545
R21497 VDD.n150 VDD 0.0209545
R21498 VDD.n207 VDD.n206 0.0185446
R21499 VDD.n141 VDD 0.0150455
R21500 VDD.n148 VDD 0.0150455
R21501 VDD.n198 VDD.n107 0.0146
R21502 VDD.n188 VDD.n111 0.0146
R21503 VDD.n160 VDD.n159 0.0137706
R21504 VDD.n213 VDD.n99 0.0101288
R21505 VDD.n102 VDD.n99 0.00994196
R21506 VDD.n212 VDD.n102 0.00918401
R21507 VDD.n208 VDD.n207 0.00868304
R21508 VDD.n163 VDD.n160 0.0073069
R21509 VDD VDD 0.00640909
R21510 VDD VDD 0.00640909
R21511 VDD.n217 VDD.n2 0.00633075
R21512 VDD.n220 VDD.n4 0.0052
R21513 VDD.n9 VDD.n6 0.0052
R21514 VDD.n97 VDD.n6 0.0050825
R21515 VDD.n138 VDD.n137 0.00321739
R21516 VDD.n140 VDD.n139 0.00321739
R21517 VDD.n145 VDD.n144 0.00321739
R21518 VDD.n147 VDD.n146 0.00321739
R21519 VDD.n152 VDD.n151 0.00321739
R21520 VDD.n154 VDD.n153 0.00321739
R21521 VDD.n8 VDD.n7 0.00298917
R21522 VDD.n218 VDD.n98 0.00298831
R21523 VDD.n143 VDD.n142 0.00239442
R21524 VDD.n150 VDD.n149 0.00239442
R21525 VDD.n219 VDD.n218 0.00202897
R21526 VDD.n7 VDD.n5 0.00201061
R21527 VDD.n96 VDD.n95 0.00152605
R21528 VDD.n95 VDD.n6 0.00151551
R21529 VDD.n187 VDD.n186 0.00125069
R21530 VDD.n193 VDD.n191 0.00125069
R21531 VDD.n215 VDD.n212 0.0011527
R21532 VDD.n176 VDD.n117 0.00109775
R21533 VDD.n209 VDD.n204 0.00105804
R21534 VDD.n4 VDD.n3 0.00102396
R21535 VDD.n214 VDD.n100 0.00101664
R21536 VDD.n216 VDD.n100 0.00101664
R21537 VDD.n214 VDD.n213 0.00101293
R21538 VDD.n221 VDD.n2 0.00101239
R21539 VDD.n213 VDD.n101 0.00101167
R21540 VDD.n4 VDD.n2 0.00101141
R21541 VDD.n218 VDD.n4 0.00100941
R21542 VDD.n7 VDD.n6 0.00100876
R21543 VDD.n174 VDD.n117 0.00100765
R21544 VDD.n93 VDD.n92 0.00100479
R21545 VDD.n212 VDD.n211 0.00100265
R21546 VDD.n1 VDD.n0 0.00100208
R21547 VDD.n186 VDD.n113 0.00100206
R21548 VDD.n193 VDD.n192 0.00100206
R21549 VDD.n219 VDD.n3 0.0010004
R21550 VDD.n142 VDD.n141 0.0010003
R21551 VDD.n149 VDD.n148 0.0010003
R21552 VDD.n206 VDD.n100 0.00100002
R21553 VDD.n176 VDD.n175 0.000990196
R21554 VDD.n171 VDD.n118 0.000990196
R21555 VDD.n167 VDD.n122 0.000990196
R21556 VDD.n185 VDD.n114 0.000990196
R21557 VDD.n178 VDD.n115 0.000990196
R21558 VDD.n177 VDD.n116 0.000990196
R21559 VDD.n170 VDD.n123 0.000990196
R21560 VDD.n169 VDD.n168 0.000990196
R21561 VDD.n184 VDD.n183 0.000990196
R21562 VDD.n181 VDD.n180 0.000990196
R21563 VDD.n196 VDD.n190 0.000990196
R21564 VDD.n200 VDD.n105 0.000990196
R21565 VDD.n195 VDD.n194 0.000990196
R21566 VDD.n201 VDD.n104 0.000990196
R21567 VDD.n208 VDD.n101 0.000709821
R21568 VDD.n173 VDD.n172 0.000684314
R21569 VDD.n166 VDD.n121 0.000684314
R21570 VDD.n120 VDD.n119 0.000684314
R21571 VDD.n159 VDD.n158 0.000684314
R21572 VDD.n187 VDD.n112 0.000684314
R21573 VDD.n182 VDD.n109 0.000684314
R21574 VDD.n179 VDD.n110 0.000684314
R21575 VDD.n191 VDD.n108 0.000684314
R21576 VDD.n197 VDD.n189 0.000684314
R21577 VDD.n199 VDD.n106 0.000684314
R21578 VDD.n216 VDD.n215 0.000517546
R21579 VDD.n215 VDD.n214 0.000517546
R21580 VDD.n216 VDD.n101 0.000517191
R21581 VDD.n173 VDD.n119 0.000516685
R21582 VDD.n158 VDD.n121 0.000516685
R21583 VDD.n172 VDD.n120 0.000516685
R21584 VDD.n166 VDD.n159 0.000516685
R21585 VDD.n199 VDD.n198 0.000516685
R21586 VDD.n198 VDD.n108 0.000516685
R21587 VDD.n188 VDD.n110 0.000516685
R21588 VDD.n182 VDD.n111 0.000516685
R21589 VDD.n179 VDD.n111 0.000516685
R21590 VDD.n188 VDD.n109 0.000516685
R21591 VDD.n188 VDD.n187 0.000516685
R21592 VDD.n112 VDD.n111 0.000516685
R21593 VDD.n189 VDD.n107 0.000516685
R21594 VDD.n198 VDD.n197 0.000516685
R21595 VDD.n191 VDD.n107 0.000516685
R21596 VDD.n107 VDD.n106 0.000516685
R21597 VDD.n204 VDD.n101 0.000512596
R21598 VDD.n219 VDD.n1 0.000505632
R21599 VDD.n96 VDD.n94 0.000505632
R21600 VDD.n93 VDD.n5 0.000505632
R21601 VDD.n222 VDD.n221 0.000505632
R21602 VDD.n173 VDD.n118 0.000505597
R21603 VDD.n122 VDD.n121 0.000505597
R21604 VDD.n175 VDD.n174 0.000505597
R21605 VDD.n172 VDD.n171 0.000505597
R21606 VDD.n167 VDD.n166 0.000505597
R21607 VDD.n183 VDD.n182 0.000505597
R21608 VDD.n181 VDD.n110 0.000505597
R21609 VDD.n180 VDD.n179 0.000505597
R21610 VDD.n184 VDD.n109 0.000505597
R21611 VDD.n113 VDD.n112 0.000505597
R21612 VDD.n197 VDD.n196 0.000505597
R21613 VDD.n200 VDD.n199 0.000505597
R21614 VDD.n192 VDD.n108 0.000505597
R21615 VDD.n190 VDD.n189 0.000505597
R21616 VDD.n106 VDD.n105 0.000505597
R21617 VDD.n94 VDD.n91 0.000504168
R21618 VDD.n223 VDD.n222 0.000504168
R21619 VDD.n123 VDD.n118 0.000504146
R21620 VDD.n169 VDD.n122 0.000504146
R21621 VDD.n175 VDD.n116 0.000504146
R21622 VDD.n171 VDD.n170 0.000504146
R21623 VDD.n168 VDD.n167 0.000504146
R21624 VDD.n177 VDD.n176 0.000504146
R21625 VDD.n183 VDD.n114 0.000504146
R21626 VDD.n180 VDD.n178 0.000504146
R21627 VDD.n181 VDD.n115 0.000504146
R21628 VDD.n185 VDD.n184 0.000504146
R21629 VDD.n196 VDD.n195 0.000504146
R21630 VDD.n201 VDD.n200 0.000504146
R21631 VDD.n194 VDD.n190 0.000504146
R21632 VDD.n105 VDD.n104 0.000504146
R21633 VDD.n209 VDD.n208 0.000503644
R21634 VDD.n206 VDD.n205 0.000502799
R21635 VDD.n205 VDD.n202 0.000502073
R21636 VDD.n210 VDD.n209 0.000502073
R21637 vcm.n386 vcm.t11 27.8779
R21638 vcm.n75 vcm.t54 27.8779
R21639 vcm.n62 vcm.t63 27.8779
R21640 vcm.n106 vcm.t70 27.8779
R21641 vcm.n120 vcm.t79 27.8779
R21642 vcm.n28 vcm.t47 27.8779
R21643 vcm.n910 vcm.t42 27.8779
R21644 vcm.n500 vcm.t37 27.8779
R21645 vcm.n296 vcm.t2 27.8779
R21646 vcm.n372 vcm.t3 27.8779
R21647 vcm.n487 vcm.t36 27.8779
R21648 vcm.n266 vcm.t33 27.8779
R21649 vcm.n186 vcm.t24 27.8779
R21650 vcm.n177 vcm.t16 27.8779
R21651 vcm.n168 vcm.t8 27.8779
R21652 vcm.n242 vcm.t17 27.8779
R21653 vcm.n231 vcm.t9 27.8779
R21654 vcm.n220 vcm.t1 27.8779
R21655 vcm.n340 vcm.t34 27.8779
R21656 vcm.n414 vcm.t27 27.8779
R21657 vcm.n471 vcm.t20 27.8779
R21658 vcm.n537 vcm.t21 27.8779
R21659 vcm.n526 vcm.t13 27.8779
R21660 vcm.n515 vcm.t5 27.8779
R21661 vcm.n714 vcm.t39 27.8779
R21662 vcm.n643 vcm.t30 27.8779
R21663 vcm.n697 vcm.t23 27.8779
R21664 vcm.n621 vcm.t14 27.8779
R21665 vcm.n680 vcm.t7 27.8779
R21666 vcm.n898 vcm.t74 27.8779
R21667 vcm.n737 vcm.t72 27.8779
R21668 vcm.n804 vcm.t73 27.8779
R21669 vcm.n954 vcm.t75 27.8779
R21670 vcm.n1073 vcm.t68 27.8779
R21671 vcm.n1062 vcm.t60 27.8779
R21672 vcm.n1161 vcm.t77 27.8779
R21673 vcm.n1148 vcm.t69 27.8779
R21674 vcm.n1126 vcm.t53 27.8779
R21675 vcm.n768 vcm.t48 27.8779
R21676 vcm.n828 vcm.t41 27.8779
R21677 vcm.n983 vcm.t51 27.8779
R21678 vcm.n1043 vcm.t44 27.8779
R21679 vcm.n39 vcm.t46 27.8779
R21680 vcm.n651 vcm.t38 27.8769
R21681 vcm.n463 vcm.t12 27.8769
R21682 vcm.n479 vcm.t28 27.8769
R21683 vcm.n422 vcm.t35 27.8769
R21684 vcm.n307 vcm.t10 27.8769
R21685 vcm.n329 vcm.t26 27.8769
R21686 vcm.n400 vcm.t19 27.8769
R21687 vcm.n548 vcm.t29 27.8769
R21688 vcm.n705 vcm.t31 27.8769
R21689 vcm.n629 vcm.t22 27.8769
R21690 vcm.n688 vcm.t15 27.8769
R21691 vcm.n607 vcm.t6 27.8769
R21692 vcm.n776 vcm.t56 27.8769
R21693 vcm.n1081 vcm.t76 27.8769
R21694 vcm.n926 vcm.t58 27.8769
R21695 vcm.n934 vcm.t66 27.8769
R21696 vcm.n836 vcm.t49 27.8769
R21697 vcm.n864 vcm.t65 27.8769
R21698 vcm.n991 vcm.t59 27.8769
R21699 vcm.n1002 vcm.t67 27.8769
R21700 vcm.n1051 vcm.t52 27.8769
R21701 vcm.n1115 vcm.t45 27.8769
R21702 vcm.n1137 vcm.t61 27.8769
R21703 vcm.n759 vcm.t40 27.8769
R21704 vcm.n1173 vcm.t78 27.8769
R21705 vcm.n97 vcm.t71 27.8769
R21706 vcm.n85 vcm.t62 27.8769
R21707 vcm.n51 vcm.t55 27.8769
R21708 vcm.n195 vcm.t32 27.8769
R21709 vcm.n253 vcm.t25 27.8769
R21710 vcm.n455 vcm.t4 27.8769
R21711 vcm.n318 vcm.t18 27.8759
R21712 vcm.n784 vcm.t64 27.8759
R21713 vcm.n850 vcm.t57 27.8759
R21714 vcm.n918 vcm.t50 27.8759
R21715 vcm.n972 vcm.t43 27.8759
R21716 vcm.n159 vcm.t0 3.2325
R21717 vcm.n11 vcm 2.29217
R21718 vcm.n906 vcm 2.29217
R21719 vcm.n559 vcm 2.29217
R21720 vcm.n289 vcm 2.29217
R21721 vcm.n362 vcm 2.29217
R21722 vcm.n425 vcm 2.29217
R21723 vcm.n147 vcm 2.29217
R21724 vcm.n264 vcm 2.29217
R21725 vcm.n154 vcm 2.29217
R21726 vcm.n213 vcm 2.29217
R21727 vcm.n281 vcm 2.29217
R21728 vcm.n451 vcm 2.29217
R21729 vcm.n508 vcm 2.29217
R21730 vcm.n597 vcm 2.29217
R21731 vcm.n672 vcm 2.29217
R21732 vcm.n878 vcm 2.29217
R21733 vcm.n1108 vcm 2.29217
R21734 vcm.n747 vcm 2.29217
R21735 vcm.n818 vcm 2.29217
R21736 vcm.n965 vcm 2.29217
R21737 vcm.n1036 vcm 2.29217
R21738 vcm.n17 vcm 2.29217
R21739 vcm.n717 vcm.n716 1.63383
R21740 vcm.n1015 vcm.n953 1.58855
R21741 vcm.n118 vcm.n101 1.57342
R21742 vcm.n93 vcm.n89 1.57342
R21743 vcm.n60 vcm.n55 1.57342
R21744 vcm.n26 vcm.n12 1.57342
R21745 vcm.n916 vcm.n915 1.57342
R21746 vcm.n908 vcm.n907 1.57342
R21747 vcm.n650 vcm.n649 1.57342
R21748 vcm.n546 vcm.n542 1.57342
R21749 vcm.n294 vcm.n290 1.57342
R21750 vcm.n384 vcm.n377 1.57342
R21751 vcm.n370 vcm.n363 1.57342
R21752 vcm.n371 vcm.n370 1.57342
R21753 vcm.n470 vcm.n469 1.57342
R21754 vcm.n488 vcm.n485 1.57342
R21755 vcm.n485 vcm.n484 1.57342
R21756 vcm.n478 vcm.n477 1.57342
R21757 vcm.n421 vcm.n420 1.57342
R21758 vcm.n265 vcm.n262 1.57342
R21759 vcm.n262 vcm.n258 1.57342
R21760 vcm.n184 vcm.n182 1.57342
R21761 vcm.n157 vcm.n155 1.57342
R21762 vcm.n230 vcm.n229 1.57342
R21763 vcm.n240 vcm.n236 1.57342
R21764 vcm.n229 vcm.n225 1.57342
R21765 vcm.n218 vcm.n214 1.57342
R21766 vcm.n219 vcm.n218 1.57342
R21767 vcm.n158 vcm.n157 1.57342
R21768 vcm.n166 vcm.n164 1.57342
R21769 vcm.n167 vcm.n166 1.57342
R21770 vcm.n175 vcm.n173 1.57342
R21771 vcm.n176 vcm.n175 1.57342
R21772 vcm.n241 vcm.n240 1.57342
R21773 vcm.n251 vcm.n247 1.57342
R21774 vcm.n252 vcm.n251 1.57342
R21775 vcm.n185 vcm.n184 1.57342
R21776 vcm.n193 vcm.n191 1.57342
R21777 vcm.n194 vcm.n193 1.57342
R21778 vcm.n327 vcm.n323 1.57342
R21779 vcm.n316 vcm.n312 1.57342
R21780 vcm.n317 vcm.n316 1.57342
R21781 vcm.n328 vcm.n327 1.57342
R21782 vcm.n338 vcm.n334 1.57342
R21783 vcm.n339 vcm.n338 1.57342
R21784 vcm.n420 vcm.n419 1.57342
R21785 vcm.n412 vcm.n405 1.57342
R21786 vcm.n413 vcm.n412 1.57342
R21787 vcm.n477 vcm.n476 1.57342
R21788 vcm.n469 vcm.n468 1.57342
R21789 vcm.n462 vcm.n461 1.57342
R21790 vcm.n461 vcm.n460 1.57342
R21791 vcm.n453 vcm.n452 1.57342
R21792 vcm.n454 vcm.n453 1.57342
R21793 vcm.n525 vcm.n524 1.57342
R21794 vcm.n535 vcm.n531 1.57342
R21795 vcm.n524 vcm.n520 1.57342
R21796 vcm.n513 vcm.n509 1.57342
R21797 vcm.n514 vcm.n513 1.57342
R21798 vcm.n295 vcm.n294 1.57342
R21799 vcm.n305 vcm.n301 1.57342
R21800 vcm.n306 vcm.n305 1.57342
R21801 vcm.n385 vcm.n384 1.57342
R21802 vcm.n398 vcm.n391 1.57342
R21803 vcm.n399 vcm.n398 1.57342
R21804 vcm.n536 vcm.n535 1.57342
R21805 vcm.n547 vcm.n546 1.57342
R21806 vcm.n557 vcm.n553 1.57342
R21807 vcm.n558 vcm.n557 1.57342
R21808 vcm.n704 vcm.n703 1.57342
R21809 vcm.n712 vcm.n710 1.57342
R21810 vcm.n713 vcm.n712 1.57342
R21811 vcm.n649 vcm.n648 1.57342
R21812 vcm.n628 vcm.n627 1.57342
R21813 vcm.n641 vcm.n634 1.57342
R21814 vcm.n642 vcm.n641 1.57342
R21815 vcm.n703 vcm.n702 1.57342
R21816 vcm.n687 vcm.n686 1.57342
R21817 vcm.n695 vcm.n693 1.57342
R21818 vcm.n696 vcm.n695 1.57342
R21819 vcm.n627 vcm.n626 1.57342
R21820 vcm.n605 vcm.n598 1.57342
R21821 vcm.n606 vcm.n605 1.57342
R21822 vcm.n619 vcm.n612 1.57342
R21823 vcm.n620 vcm.n619 1.57342
R21824 vcm.n686 vcm.n685 1.57342
R21825 vcm.n678 vcm.n673 1.57342
R21826 vcm.n679 vcm.n678 1.57342
R21827 vcm.n1080 vcm.n1079 1.57342
R21828 vcm.n932 vcm.n931 1.57342
R21829 vcm.n933 vcm.n932 1.57342
R21830 vcm.n940 vcm.n939 1.57342
R21831 vcm.n941 vcm.n940 1.57342
R21832 vcm.n783 vcm.n782 1.57342
R21833 vcm.n791 vcm.n789 1.57342
R21834 vcm.n792 vcm.n791 1.57342
R21835 vcm.n862 vcm.n855 1.57342
R21836 vcm.n848 vcm.n841 1.57342
R21837 vcm.n835 vcm.n834 1.57342
R21838 vcm.n849 vcm.n848 1.57342
R21839 vcm.n863 vcm.n862 1.57342
R21840 vcm.n876 vcm.n869 1.57342
R21841 vcm.n877 vcm.n876 1.57342
R21842 vcm.n1000 vcm.n996 1.57342
R21843 vcm.n990 vcm.n989 1.57342
R21844 vcm.n1001 vcm.n1000 1.57342
R21845 vcm.n1011 vcm.n1007 1.57342
R21846 vcm.n1012 vcm.n1011 1.57342
R21847 vcm.n1079 vcm.n1078 1.57342
R21848 vcm.n1050 vcm.n1049 1.57342
R21849 vcm.n1060 vcm.n1056 1.57342
R21850 vcm.n1061 vcm.n1060 1.57342
R21851 vcm.n1071 vcm.n1067 1.57342
R21852 vcm.n1072 vcm.n1071 1.57342
R21853 vcm.n1160 vcm.n1157 1.57342
R21854 vcm.n1157 vcm.n1153 1.57342
R21855 vcm.n1135 vcm.n1131 1.57342
R21856 vcm.n1113 vcm.n1109 1.57342
R21857 vcm.n1114 vcm.n1113 1.57342
R21858 vcm.n1124 vcm.n1120 1.57342
R21859 vcm.n1125 vcm.n1124 1.57342
R21860 vcm.n1136 vcm.n1135 1.57342
R21861 vcm.n1146 vcm.n1142 1.57342
R21862 vcm.n1147 vcm.n1146 1.57342
R21863 vcm.n782 vcm.n781 1.57342
R21864 vcm.n775 vcm.n774 1.57342
R21865 vcm.n774 vcm.n773 1.57342
R21866 vcm.n757 vcm.n748 1.57342
R21867 vcm.n758 vcm.n757 1.57342
R21868 vcm.n766 vcm.n764 1.57342
R21869 vcm.n767 vcm.n766 1.57342
R21870 vcm.n834 vcm.n833 1.57342
R21871 vcm.n826 vcm.n819 1.57342
R21872 vcm.n827 vcm.n826 1.57342
R21873 vcm.n909 vcm.n908 1.57342
R21874 vcm.n917 vcm.n916 1.57342
R21875 vcm.n924 vcm.n923 1.57342
R21876 vcm.n925 vcm.n924 1.57342
R21877 vcm.n989 vcm.n988 1.57342
R21878 vcm.n970 vcm.n966 1.57342
R21879 vcm.n971 vcm.n970 1.57342
R21880 vcm.n981 vcm.n977 1.57342
R21881 vcm.n982 vcm.n981 1.57342
R21882 vcm.n1049 vcm.n1048 1.57342
R21883 vcm.n1041 vcm.n1037 1.57342
R21884 vcm.n1042 vcm.n1041 1.57342
R21885 vcm.n47 vcm.n43 1.57342
R21886 vcm.n22 vcm.n18 1.57342
R21887 vcm.n27 vcm.n26 1.57342
R21888 vcm.n49 vcm.n32 1.57342
R21889 vcm.n50 vcm.n49 1.57342
R21890 vcm.n83 vcm.n79 1.57342
R21891 vcm.n84 vcm.n83 1.57342
R21892 vcm.n61 vcm.n60 1.57342
R21893 vcm.n95 vcm.n66 1.57342
R21894 vcm.n96 vcm.n95 1.57342
R21895 vcm.n114 vcm.n110 1.57342
R21896 vcm.n121 vcm.n118 1.57342
R21897 vcm.n1015 vcm.n1014 1.49217
R21898 vcm.n717 vcm.n715 1.44689
R21899 vcm.n944 vcm.n943 1.42133
R21900 vcm.n491 vcm.n490 1.4005
R21901 vcm.n1177 vcm.n1176 1.388
R21902 vcm.n1188 vcm.n1187 1.388
R21903 vcm.n1176 vcm 1.14633
R21904 vcm.n654 vcm 1.14633
R21905 vcm.n490 vcm 1.14633
R21906 vcm.n716 vcm 1.14633
R21907 vcm.n1021 vcm 1.14633
R21908 vcm.n943 vcm 1.14633
R21909 vcm.n794 vcm 1.14633
R21910 vcm.n1014 vcm 1.14633
R21911 vcm.n1158 vcm 1.14633
R21912 vcm vcm.n1188 1.14633
R21913 vcm.n157 vcm.n156 1.1065
R21914 vcm.n166 vcm.n165 1.1065
R21915 vcm.n175 vcm.n174 1.1065
R21916 vcm.n184 vcm.n183 1.1065
R21917 vcm.n193 vcm.n192 1.1065
R21918 vcm.n791 vcm.n790 1.1065
R21919 vcm.n782 vcm.n739 1.1065
R21920 vcm.n774 vcm.n741 1.1065
R21921 vcm.n766 vcm.n765 1.1065
R21922 vcm.n712 vcm.n711 1.101
R21923 vcm.n703 vcm.n664 1.101
R21924 vcm.n695 vcm.n694 1.101
R21925 vcm.n686 vcm.n667 1.101
R21926 vcm.n26 vcm.n13 1.101
R21927 vcm.n49 vcm.n33 1.101
R21928 vcm.n60 vcm.n56 1.101
R21929 vcm.n95 vcm.n67 1.101
R21930 vcm.n118 vcm.n102 1.101
R21931 vcm.n218 vcm.n217 1.1005
R21932 vcm.n240 vcm.n239 1.1005
R21933 vcm.n251 vcm.n250 1.1005
R21934 vcm.n338 vcm.n337 1.1005
R21935 vcm.n262 vcm.n261 1.1005
R21936 vcm.n420 vcm.n351 1.1005
R21937 vcm.n420 vcm.n354 1.1005
R21938 vcm.n412 vcm.n408 1.1005
R21939 vcm.n412 vcm.n411 1.1005
R21940 vcm.n327 vcm.n326 1.1005
R21941 vcm.n513 vcm.n512 1.1005
R21942 vcm.n370 vcm.n366 1.1005
R21943 vcm.n370 vcm.n369 1.1005
R21944 vcm.n294 vcm.n293 1.1005
R21945 vcm.n305 vcm.n304 1.1005
R21946 vcm.n229 vcm.n228 1.1005
R21947 vcm.n384 vcm.n380 1.1005
R21948 vcm.n384 vcm.n383 1.1005
R21949 vcm.n398 vcm.n394 1.1005
R21950 vcm.n398 vcm.n397 1.1005
R21951 vcm.n316 vcm.n315 1.1005
R21952 vcm.n535 vcm.n534 1.1005
R21953 vcm.n557 vcm.n556 1.1005
R21954 vcm.n649 vcm.n580 1.1005
R21955 vcm.n649 vcm.n583 1.1005
R21956 vcm.n641 vcm.n637 1.1005
R21957 vcm.n641 vcm.n640 1.1005
R21958 vcm.n546 vcm.n545 1.1005
R21959 vcm.n627 vcm.n588 1.1005
R21960 vcm.n627 vcm.n591 1.1005
R21961 vcm.n619 vcm.n615 1.1005
R21962 vcm.n619 vcm.n618 1.1005
R21963 vcm.n524 vcm.n523 1.1005
R21964 vcm.n678 vcm.n677 1.1005
R21965 vcm.n605 vcm.n601 1.1005
R21966 vcm.n605 vcm.n604 1.1005
R21967 vcm.n876 vcm.n872 1.1005
R21968 vcm.n876 vcm.n875 1.1005
R21969 vcm.n1011 vcm.n1010 1.1005
R21970 vcm.n1079 vcm.n1025 1.1005
R21971 vcm.n1060 vcm.n1059 1.1005
R21972 vcm.n1124 vcm.n1123 1.1005
R21973 vcm.n1146 vcm.n1145 1.1005
R21974 vcm.n1071 vcm.n1070 1.1005
R21975 vcm.n1000 vcm.n999 1.1005
R21976 vcm.n862 vcm.n858 1.1005
R21977 vcm.n862 vcm.n861 1.1005
R21978 vcm.n834 vcm.n810 1.1005
R21979 vcm.n834 vcm.n813 1.1005
R21980 vcm.n826 vcm.n822 1.1005
R21981 vcm.n826 vcm.n825 1.1005
R21982 vcm.n757 vcm.n756 1.1005
R21983 vcm.n848 vcm.n844 1.1005
R21984 vcm.n848 vcm.n847 1.1005
R21985 vcm.n989 vcm.n959 1.1005
R21986 vcm.n981 vcm.n980 1.1005
R21987 vcm.n1049 vcm.n1031 1.1005
R21988 vcm.n1041 vcm.n1040 1.1005
R21989 vcm.n970 vcm.n969 1.1005
R21990 vcm.n25 vcm.n22 1.1005
R21991 vcm.n22 vcm.n21 1.1005
R21992 vcm.n1113 vcm.n1112 1.1005
R21993 vcm.n26 vcm.n25 1.1005
R21994 vcm.n49 vcm.n48 1.1005
R21995 vcm.n48 vcm.n47 1.1005
R21996 vcm.n47 vcm.n46 1.1005
R21997 vcm.n83 vcm.n82 1.1005
R21998 vcm.n1135 vcm.n1134 1.1005
R21999 vcm.n60 vcm.n59 1.1005
R22000 vcm.n95 vcm.n94 1.1005
R22001 vcm.n94 vcm.n93 1.1005
R22002 vcm.n93 vcm.n92 1.1005
R22003 vcm.n117 vcm.n114 1.1005
R22004 vcm.n114 vcm.n113 1.1005
R22005 vcm.n1157 vcm.n1156 1.1005
R22006 vcm.n118 vcm.n117 1.1005
R22007 vcm.n730 vcm.n729 1.05236
R22008 vcm.n426 vcm.n425 1.013
R22009 vcm.n655 vcm.n654 0.971333
R22010 vcm.n655 vcm.n652 0.9255
R22011 vcm.n426 vcm.n423 0.921888
R22012 vcm.n197 vcm.n196 0.822638
R22013 vcm.n268 vcm.n267 0.821888
R22014 vcm.n729 vcm.n728 0.78775
R22015 vcm.n342 vcm.n341 0.771888
R22016 vcm.n560 vcm.n559 0.7005
R22017 vcm.n795 vcm.n794 0.6755
R22018 vcm.n879 vcm.n878 0.604667
R22019 vcm.n1083 vcm.n1082 0.567167
R22020 vcm.n1163 vcm.n1162 0.563
R22021 vcm.n1178 vcm.n1177 0.539716
R22022 vcm.n656 vcm.n655 0.539716
R22023 vcm.n561 vcm.n560 0.539716
R22024 vcm.n492 vcm.n491 0.539716
R22025 vcm.n427 vcm.n426 0.539716
R22026 vcm.n198 vcm.n197 0.539716
R22027 vcm.n269 vcm.n268 0.539716
R22028 vcm.n343 vcm.n342 0.539716
R22029 vcm.n718 vcm.n717 0.539716
R22030 vcm.n1084 vcm.n1083 0.539716
R22031 vcm.n945 vcm.n944 0.539716
R22032 vcm.n796 vcm.n795 0.539716
R22033 vcm.n880 vcm.n879 0.539716
R22034 vcm.n1016 vcm.n1015 0.539716
R22035 vcm.n1164 vcm.n1163 0.539716
R22036 vcm.n1187 vcm.n1186 0.539716
R22037 vcm.n801 vcm.n800 0.48695
R22038 vcm.n661 vcm.n660 0.475318
R22039 vcm.n497 vcm.n496 0.469208
R22040 vcm.n950 vcm.n949 0.458633
R22041 vcm.n1169 vcm.n1168 0.458162
R22042 vcm.n274 vcm.n273 0.458045
R22043 vcm.n1095 vcm.n1094 0.456753
R22044 vcm.n1183 vcm.n1182 0.456635
R22045 vcm.n203 vcm.n202 0.456635
R22046 vcm.n348 vcm.n347 0.452405
R22047 vcm.n1087 vcm.n1020 0.452052
R22048 vcm.n891 vcm.n890 0.447353
R22049 vcm.n438 vcm.n437 0.43525
R22050 vcm.n572 vcm.n571 0.43196
R22051 vcm vcm.n98 0.3755
R22052 vcm vcm.n86 0.3755
R22053 vcm vcm.n52 0.3755
R22054 vcm vcm.n373 0.3755
R22055 vcm vcm.n480 0.3755
R22056 vcm vcm.n254 0.3755
R22057 vcm vcm.n178 0.3755
R22058 vcm vcm.n232 0.3755
R22059 vcm vcm.n221 0.3755
R22060 vcm vcm.n160 0.3755
R22061 vcm vcm.n169 0.3755
R22062 vcm vcm.n243 0.3755
R22063 vcm vcm.n187 0.3755
R22064 vcm vcm.n308 0.3755
R22065 vcm vcm.n319 0.3755
R22066 vcm vcm.n330 0.3755
R22067 vcm vcm.n415 0.3755
R22068 vcm vcm.n401 0.3755
R22069 vcm vcm.n472 0.3755
R22070 vcm vcm.n464 0.3755
R22071 vcm vcm.n456 0.3755
R22072 vcm vcm.n527 0.3755
R22073 vcm vcm.n516 0.3755
R22074 vcm vcm.n297 0.3755
R22075 vcm vcm.n387 0.3755
R22076 vcm vcm.n538 0.3755
R22077 vcm vcm.n549 0.3755
R22078 vcm vcm.n706 0.3755
R22079 vcm vcm.n644 0.3755
R22080 vcm vcm.n630 0.3755
R22081 vcm vcm.n698 0.3755
R22082 vcm vcm.n689 0.3755
R22083 vcm vcm.n622 0.3755
R22084 vcm vcm.n608 0.3755
R22085 vcm vcm.n681 0.3755
R22086 vcm vcm.n927 0.3755
R22087 vcm vcm.n935 0.3755
R22088 vcm vcm.n785 0.3755
R22089 vcm vcm.n837 0.3755
R22090 vcm vcm.n851 0.3755
R22091 vcm vcm.n865 0.3755
R22092 vcm vcm.n992 0.3755
R22093 vcm vcm.n1003 0.3755
R22094 vcm vcm.n1074 0.3755
R22095 vcm vcm.n1052 0.3755
R22096 vcm vcm.n1063 0.3755
R22097 vcm vcm.n1149 0.3755
R22098 vcm vcm.n1116 0.3755
R22099 vcm vcm.n1127 0.3755
R22100 vcm vcm.n1138 0.3755
R22101 vcm vcm.n777 0.3755
R22102 vcm vcm.n769 0.3755
R22103 vcm vcm.n760 0.3755
R22104 vcm vcm.n829 0.3755
R22105 vcm vcm.n911 0.3755
R22106 vcm vcm.n919 0.3755
R22107 vcm vcm.n984 0.3755
R22108 vcm vcm.n973 0.3755
R22109 vcm vcm.n1044 0.3755
R22110 vcm vcm.n40 0.3755
R22111 vcm vcm.n29 0.3755
R22112 vcm vcm.n76 0.3755
R22113 vcm vcm.n63 0.3755
R22114 vcm vcm.n107 0.3755
R22115 vcm.n8 vcm 0.234474
R22116 vcm.n903 vcm 0.234474
R22117 vcm.n652 vcm 0.234474
R22118 vcm.n286 vcm 0.234474
R22119 vcm.n359 vcm 0.234474
R22120 vcm.n152 vcm 0.234474
R22121 vcm.n210 vcm 0.234474
R22122 vcm.n448 vcm 0.234474
R22123 vcm.n505 vcm 0.234474
R22124 vcm.n594 vcm 0.234474
R22125 vcm.n669 vcm 0.234474
R22126 vcm.n1082 vcm 0.234474
R22127 vcm.n736 vcm 0.234474
R22128 vcm.n1162 vcm 0.234474
R22129 vcm.n1105 vcm 0.234474
R22130 vcm.n744 vcm 0.234474
R22131 vcm.n815 vcm 0.234474
R22132 vcm.n962 vcm 0.234474
R22133 vcm.n1033 vcm 0.234474
R22134 vcm.n14 vcm 0.234474
R22135 vcm.n664 vcm 0.187646
R22136 vcm.n667 vcm 0.187646
R22137 vcm.n13 vcm 0.187646
R22138 vcm.n56 vcm 0.187646
R22139 vcm.n102 vcm 0.187646
R22140 vcm.n711 vcm 0.186894
R22141 vcm.n694 vcm 0.186894
R22142 vcm.n33 vcm 0.186894
R22143 vcm.n67 vcm 0.186894
R22144 vcm.n156 vcm 0.185131
R22145 vcm.n165 vcm 0.185131
R22146 vcm.n183 vcm 0.185131
R22147 vcm.n790 vcm 0.185131
R22148 vcm.n739 vcm 0.185131
R22149 vcm.n741 vcm 0.185131
R22150 vcm.n174 vcm 0.185131
R22151 vcm.n192 vcm 0.185131
R22152 vcm.n765 vcm 0.185131
R22153 vcm.n98 vcm 0.117487
R22154 vcm.n86 vcm 0.117487
R22155 vcm.n52 vcm 0.117487
R22156 vcm.n373 vcm 0.117487
R22157 vcm.n480 vcm 0.117487
R22158 vcm.n254 vcm 0.117487
R22159 vcm.n178 vcm 0.117487
R22160 vcm.n232 vcm 0.117487
R22161 vcm.n221 vcm 0.117487
R22162 vcm.n160 vcm 0.117487
R22163 vcm.n169 vcm 0.117487
R22164 vcm.n243 vcm 0.117487
R22165 vcm.n187 vcm 0.117487
R22166 vcm.n308 vcm 0.117487
R22167 vcm.n319 vcm 0.117487
R22168 vcm.n330 vcm 0.117487
R22169 vcm.n415 vcm 0.117487
R22170 vcm.n401 vcm 0.117487
R22171 vcm.n472 vcm 0.117487
R22172 vcm.n464 vcm 0.117487
R22173 vcm.n456 vcm 0.117487
R22174 vcm.n527 vcm 0.117487
R22175 vcm.n516 vcm 0.117487
R22176 vcm.n297 vcm 0.117487
R22177 vcm.n387 vcm 0.117487
R22178 vcm.n538 vcm 0.117487
R22179 vcm.n549 vcm 0.117487
R22180 vcm.n706 vcm 0.117487
R22181 vcm.n644 vcm 0.117487
R22182 vcm.n630 vcm 0.117487
R22183 vcm.n698 vcm 0.117487
R22184 vcm.n689 vcm 0.117487
R22185 vcm.n622 vcm 0.117487
R22186 vcm.n608 vcm 0.117487
R22187 vcm.n681 vcm 0.117487
R22188 vcm.n927 vcm 0.117487
R22189 vcm.n935 vcm 0.117487
R22190 vcm.n785 vcm 0.117487
R22191 vcm.n837 vcm 0.117487
R22192 vcm.n851 vcm 0.117487
R22193 vcm.n865 vcm 0.117487
R22194 vcm.n992 vcm 0.117487
R22195 vcm.n1003 vcm 0.117487
R22196 vcm.n1074 vcm 0.117487
R22197 vcm.n1052 vcm 0.117487
R22198 vcm.n1063 vcm 0.117487
R22199 vcm.n1149 vcm 0.117487
R22200 vcm.n1116 vcm 0.117487
R22201 vcm.n1127 vcm 0.117487
R22202 vcm.n1138 vcm 0.117487
R22203 vcm.n777 vcm 0.117487
R22204 vcm.n769 vcm 0.117487
R22205 vcm.n760 vcm 0.117487
R22206 vcm.n829 vcm 0.117487
R22207 vcm.n911 vcm 0.117487
R22208 vcm.n919 vcm 0.117487
R22209 vcm.n984 vcm 0.117487
R22210 vcm.n973 vcm 0.117487
R22211 vcm.n1044 vcm 0.117487
R22212 vcm.n40 vcm 0.117487
R22213 vcm.n29 vcm 0.117487
R22214 vcm.n76 vcm 0.117487
R22215 vcm.n63 vcm 0.117487
R22216 vcm.n107 vcm 0.117487
R22217 vcm.n10 vcm 0.117222
R22218 vcm.n905 vcm 0.117222
R22219 vcm.n288 vcm 0.117222
R22220 vcm.n361 vcm 0.117222
R22221 vcm.n153 vcm 0.117222
R22222 vcm.n212 vcm 0.117222
R22223 vcm.n450 vcm 0.117222
R22224 vcm.n507 vcm 0.117222
R22225 vcm.n596 vcm 0.117222
R22226 vcm.n671 vcm 0.117222
R22227 vcm.n1107 vcm 0.117222
R22228 vcm.n746 vcm 0.117222
R22229 vcm.n817 vcm 0.117222
R22230 vcm.n964 vcm 0.117222
R22231 vcm.n1035 vcm 0.117222
R22232 vcm.n16 vcm 0.117222
R22233 vcm.n498 vcm 0.105191
R22234 vcm.n424 vcm 0.105191
R22235 vcm.n146 vcm 0.105191
R22236 vcm.n263 vcm 0.105191
R22237 vcm.n280 vcm 0.105191
R22238 vcm.n802 vcm 0.105191
R22239 vcm.n260 vcm 0.0970784
R22240 vcm.n336 vcm 0.0970784
R22241 vcm.n353 vcm 0.0970784
R22242 vcm.n410 vcm 0.0970784
R22243 vcm.n407 vcm 0.0970784
R22244 vcm.n511 vcm 0.0970784
R22245 vcm.n396 vcm 0.0970784
R22246 vcm.n393 vcm 0.0970784
R22247 vcm.n555 vcm 0.0970784
R22248 vcm.n582 vcm 0.0970784
R22249 vcm.n639 vcm 0.0970784
R22250 vcm.n636 vcm 0.0970784
R22251 vcm.n590 vcm 0.0970784
R22252 vcm.n617 vcm 0.0970784
R22253 vcm.n614 vcm 0.0970784
R22254 vcm.n600 vcm 0.0970784
R22255 vcm.n1069 vcm 0.0970784
R22256 vcm.n998 vcm 0.0970784
R22257 vcm.n857 vcm 0.0970784
R22258 vcm.n824 vcm 0.0970784
R22259 vcm.n821 vcm 0.0970784
R22260 vcm.n843 vcm 0.0970784
R22261 vcm.n958 vcm 0.0970784
R22262 vcm.n979 vcm 0.0970784
R22263 vcm.n1030 vcm 0.0970784
R22264 vcm.n35 vcm 0.0965779
R22265 vcm.n69 vcm 0.0965779
R22266 vcm.n325 vcm 0.0965766
R22267 vcm.n350 vcm 0.0965766
R22268 vcm.n544 vcm 0.0965766
R22269 vcm.n603 vcm 0.0965766
R22270 vcm.n522 vcm 0.0965766
R22271 vcm.n379 vcm 0.0965766
R22272 vcm.n533 vcm 0.0965766
R22273 vcm.n579 vcm 0.0965766
R22274 vcm.n587 vcm 0.0965766
R22275 vcm.n1144 vcm 0.0965766
R22276 vcm.n860 vcm 0.0965766
R22277 vcm.n968 vcm 0.0965766
R22278 vcm.n1133 vcm 0.0965766
R22279 vcm.n1058 vcm 0.0965766
R22280 vcm.n1122 vcm 0.0965766
R22281 vcm.n216 vcm 0.0958266
R22282 vcm.n227 vcm 0.0958266
R22283 vcm.n314 vcm 0.0958266
R22284 vcm.n249 vcm 0.0958266
R22285 vcm.n365 vcm 0.0958266
R22286 vcm.n368 vcm 0.0958266
R22287 vcm.n303 vcm 0.0958266
R22288 vcm.n874 vcm 0.0958266
R22289 vcm.n1009 vcm 0.0958266
R22290 vcm.n1155 vcm 0.0958266
R22291 vcm.n846 vcm 0.0958266
R22292 vcm.n809 vcm 0.0958266
R22293 vcm.n1039 vcm 0.0958266
R22294 vcm.n20 vcm 0.0958266
R22295 vcm.n81 vcm 0.0958266
R22296 vcm.n112 vcm 0.0958266
R22297 vcm.n238 vcm 0.0956149
R22298 vcm.n292 vcm 0.0956149
R22299 vcm.n382 vcm 0.0956149
R22300 vcm.n871 vcm 0.0956149
R22301 vcm.n1024 vcm 0.0956149
R22302 vcm.n812 vcm 0.0956149
R22303 vcm.n1111 vcm 0.0956149
R22304 vcm.n24 vcm 0.0956149
R22305 vcm.n45 vcm 0.0956149
R22306 vcm.n58 vcm 0.0956149
R22307 vcm.n91 vcm 0.0956149
R22308 vcm.n116 vcm 0.0956149
R22309 vcm.n676 vcm.n675 0.0955985
R22310 vcm.n1175 vcm.n1174 0.0915799
R22311 vcm.n489 vcm.n488 0.0915799
R22312 vcm.n713 vcm.n662 0.0915799
R22313 vcm.n1080 vcm.n1022 0.0915799
R22314 vcm.n942 vcm.n941 0.0915799
R22315 vcm.n793 vcm.n792 0.0915799
R22316 vcm.n1013 vcm.n1012 0.0915799
R22317 vcm.n1160 vcm.n1159 0.0915799
R22318 vcm.n122 vcm.n121 0.0915799
R22319 vcm.n101 vcm.n100 0.0914585
R22320 vcm.n89 vcm.n88 0.0914585
R22321 vcm.n55 vcm.n54 0.0914585
R22322 vcm.n377 vcm.n376 0.0914585
R22323 vcm.n484 vcm.n483 0.0914585
R22324 vcm.n258 vcm.n257 0.0914585
R22325 vcm.n182 vcm.n181 0.0914585
R22326 vcm.n236 vcm.n235 0.0914585
R22327 vcm.n225 vcm.n224 0.0914585
R22328 vcm.n164 vcm.n163 0.0914585
R22329 vcm.n173 vcm.n172 0.0914585
R22330 vcm.n247 vcm.n246 0.0914585
R22331 vcm.n191 vcm.n190 0.0914585
R22332 vcm.n312 vcm.n311 0.0914585
R22333 vcm.n323 vcm.n322 0.0914585
R22334 vcm.n334 vcm.n333 0.0914585
R22335 vcm.n419 vcm.n418 0.0914585
R22336 vcm.n405 vcm.n404 0.0914585
R22337 vcm.n476 vcm.n475 0.0914585
R22338 vcm.n468 vcm.n467 0.0914585
R22339 vcm.n460 vcm.n459 0.0914585
R22340 vcm.n531 vcm.n530 0.0914585
R22341 vcm.n520 vcm.n519 0.0914585
R22342 vcm.n301 vcm.n300 0.0914585
R22343 vcm.n391 vcm.n390 0.0914585
R22344 vcm.n542 vcm.n541 0.0914585
R22345 vcm.n553 vcm.n552 0.0914585
R22346 vcm.n710 vcm.n709 0.0914585
R22347 vcm.n648 vcm.n647 0.0914585
R22348 vcm.n634 vcm.n633 0.0914585
R22349 vcm.n702 vcm.n701 0.0914585
R22350 vcm.n693 vcm.n692 0.0914585
R22351 vcm.n626 vcm.n625 0.0914585
R22352 vcm.n612 vcm.n611 0.0914585
R22353 vcm.n685 vcm.n684 0.0914585
R22354 vcm.n931 vcm.n930 0.0914585
R22355 vcm.n939 vcm.n938 0.0914585
R22356 vcm.n789 vcm.n788 0.0914585
R22357 vcm.n841 vcm.n840 0.0914585
R22358 vcm.n855 vcm.n854 0.0914585
R22359 vcm.n869 vcm.n868 0.0914585
R22360 vcm.n996 vcm.n995 0.0914585
R22361 vcm.n1007 vcm.n1006 0.0914585
R22362 vcm.n1078 vcm.n1077 0.0914585
R22363 vcm.n1056 vcm.n1055 0.0914585
R22364 vcm.n1067 vcm.n1066 0.0914585
R22365 vcm.n1153 vcm.n1152 0.0914585
R22366 vcm.n1120 vcm.n1119 0.0914585
R22367 vcm.n1131 vcm.n1130 0.0914585
R22368 vcm.n1142 vcm.n1141 0.0914585
R22369 vcm.n781 vcm.n780 0.0914585
R22370 vcm.n773 vcm.n772 0.0914585
R22371 vcm.n764 vcm.n763 0.0914585
R22372 vcm.n833 vcm.n832 0.0914585
R22373 vcm.n915 vcm.n914 0.0914585
R22374 vcm.n923 vcm.n922 0.0914585
R22375 vcm.n988 vcm.n987 0.0914585
R22376 vcm.n977 vcm.n976 0.0914585
R22377 vcm.n1048 vcm.n1047 0.0914585
R22378 vcm.n43 vcm.n42 0.0914585
R22379 vcm.n32 vcm.n31 0.0914585
R22380 vcm.n79 vcm.n78 0.0914585
R22381 vcm.n66 vcm.n65 0.0914585
R22382 vcm.n110 vcm.n109 0.0914585
R22383 vcm.n196 vcm.n195 0.0888628
R22384 vcm.n1173 vcm.n1172 0.0888625
R22385 vcm.n500 vcm.n499 0.0888625
R22386 vcm.n487 vcm.n486 0.0888625
R22387 vcm.n423 vcm.n422 0.0888625
R22388 vcm.n267 vcm.n266 0.0888625
R22389 vcm.n341 vcm.n340 0.0888625
R22390 vcm.n715 vcm.n714 0.0888625
R22391 vcm.n898 vcm.n897 0.0888625
R22392 vcm.n804 vcm.n803 0.0888625
R22393 vcm.n120 vcm.n119 0.0888625
R22394 vcm.n674 vcm 0.0635002
R22395 vcm.n750 vcm 0.063
R22396 vcm.n729 vcm 0.0617502
R22397 vcm.n12 vcm.n11 0.049413
R22398 vcm.n907 vcm.n906 0.049413
R22399 vcm.n559 vcm.n558 0.049413
R22400 vcm.n290 vcm.n289 0.049413
R22401 vcm.n363 vcm.n362 0.049413
R22402 vcm.n194 vcm.n147 0.049413
R22403 vcm.n265 vcm.n264 0.049413
R22404 vcm.n155 vcm.n152 0.049413
R22405 vcm.n155 vcm.n154 0.049413
R22406 vcm.n214 vcm.n213 0.049413
R22407 vcm.n339 vcm.n281 0.049413
R22408 vcm.n452 vcm.n451 0.049413
R22409 vcm.n509 vcm.n508 0.049413
R22410 vcm.n598 vcm.n597 0.049413
R22411 vcm.n673 vcm.n672 0.049413
R22412 vcm.n878 vcm.n877 0.049413
R22413 vcm.n1109 vcm.n1108 0.049413
R22414 vcm.n748 vcm.n747 0.049413
R22415 vcm.n819 vcm.n818 0.049413
R22416 vcm.n966 vcm.n965 0.049413
R22417 vcm.n1037 vcm.n1036 0.049413
R22418 vcm.n18 vcm.n17 0.049413
R22419 vcm.n98 vcm.n0 0.0466957
R22420 vcm.n98 vcm.n97 0.0466957
R22421 vcm.n86 vcm.n70 0.0466957
R22422 vcm.n86 vcm.n85 0.0466957
R22423 vcm.n52 vcm.n4 0.0466957
R22424 vcm.n52 vcm.n51 0.0466957
R22425 vcm.n9 vcm.n8 0.0466957
R22426 vcm.n904 vcm.n903 0.0466957
R22427 vcm.n652 vcm.n651 0.0466957
R22428 vcm.n287 vcm.n286 0.0466957
R22429 vcm.n373 vcm.n358 0.0466957
R22430 vcm.n373 vcm.n372 0.0466957
R22431 vcm.n360 vcm.n359 0.0466957
R22432 vcm.n480 vcm.n444 0.0466957
R22433 vcm.n480 vcm.n479 0.0466957
R22434 vcm.n254 vcm.n206 0.0466957
R22435 vcm.n254 vcm.n253 0.0466957
R22436 vcm.n178 vcm.n149 0.0466957
R22437 vcm.n178 vcm.n177 0.0466957
R22438 vcm.n232 vcm.n208 0.0466957
R22439 vcm.n232 vcm.n231 0.0466957
R22440 vcm.n221 vcm.n209 0.0466957
R22441 vcm.n221 vcm.n220 0.0466957
R22442 vcm.n211 vcm.n210 0.0466957
R22443 vcm.n160 vcm.n159 0.0466957
R22444 vcm.n160 vcm.n151 0.0466957
R22445 vcm.n169 vcm.n168 0.0466957
R22446 vcm.n169 vcm.n150 0.0466957
R22447 vcm.n243 vcm.n242 0.0466957
R22448 vcm.n243 vcm.n207 0.0466957
R22449 vcm.n187 vcm.n186 0.0466957
R22450 vcm.n187 vcm.n148 0.0466957
R22451 vcm.n308 vcm.n307 0.0466957
R22452 vcm.n308 vcm.n284 0.0466957
R22453 vcm.n319 vcm.n318 0.0466957
R22454 vcm.n319 vcm.n283 0.0466957
R22455 vcm.n330 vcm.n329 0.0466957
R22456 vcm.n330 vcm.n282 0.0466957
R22457 vcm.n415 vcm.n355 0.0466957
R22458 vcm.n415 vcm.n414 0.0466957
R22459 vcm.n401 vcm.n400 0.0466957
R22460 vcm.n401 vcm.n356 0.0466957
R22461 vcm.n472 vcm.n445 0.0466957
R22462 vcm.n472 vcm.n471 0.0466957
R22463 vcm.n464 vcm.n446 0.0466957
R22464 vcm.n464 vcm.n463 0.0466957
R22465 vcm.n456 vcm.n447 0.0466957
R22466 vcm.n456 vcm.n455 0.0466957
R22467 vcm.n449 vcm.n448 0.0466957
R22468 vcm.n527 vcm.n503 0.0466957
R22469 vcm.n527 vcm.n526 0.0466957
R22470 vcm.n516 vcm.n504 0.0466957
R22471 vcm.n516 vcm.n515 0.0466957
R22472 vcm.n506 vcm.n505 0.0466957
R22473 vcm.n297 vcm.n296 0.0466957
R22474 vcm.n297 vcm.n285 0.0466957
R22475 vcm.n387 vcm.n386 0.0466957
R22476 vcm.n387 vcm.n357 0.0466957
R22477 vcm.n538 vcm.n537 0.0466957
R22478 vcm.n538 vcm.n502 0.0466957
R22479 vcm.n549 vcm.n548 0.0466957
R22480 vcm.n549 vcm.n501 0.0466957
R22481 vcm.n706 vcm.n705 0.0466957
R22482 vcm.n706 vcm.n663 0.0466957
R22483 vcm.n644 vcm.n584 0.0466957
R22484 vcm.n644 vcm.n643 0.0466957
R22485 vcm.n630 vcm.n629 0.0466957
R22486 vcm.n630 vcm.n585 0.0466957
R22487 vcm.n698 vcm.n665 0.0466957
R22488 vcm.n698 vcm.n697 0.0466957
R22489 vcm.n689 vcm.n688 0.0466957
R22490 vcm.n689 vcm.n666 0.0466957
R22491 vcm.n622 vcm.n592 0.0466957
R22492 vcm.n622 vcm.n621 0.0466957
R22493 vcm.n595 vcm.n594 0.0466957
R22494 vcm.n608 vcm.n607 0.0466957
R22495 vcm.n608 vcm.n593 0.0466957
R22496 vcm.n681 vcm.n668 0.0466957
R22497 vcm.n681 vcm.n680 0.0466957
R22498 vcm.n670 vcm.n669 0.0466957
R22499 vcm.n1082 vcm.n1081 0.0466957
R22500 vcm.n927 vcm.n926 0.0466957
R22501 vcm.n927 vcm.n900 0.0466957
R22502 vcm.n935 vcm.n934 0.0466957
R22503 vcm.n935 vcm.n899 0.0466957
R22504 vcm.n737 vcm.n736 0.0466957
R22505 vcm.n785 vcm.n784 0.0466957
R22506 vcm.n785 vcm.n738 0.0466957
R22507 vcm.n837 vcm.n836 0.0466957
R22508 vcm.n837 vcm.n807 0.0466957
R22509 vcm.n851 vcm.n850 0.0466957
R22510 vcm.n851 vcm.n806 0.0466957
R22511 vcm.n865 vcm.n864 0.0466957
R22512 vcm.n865 vcm.n805 0.0466957
R22513 vcm.n992 vcm.n991 0.0466957
R22514 vcm.n992 vcm.n956 0.0466957
R22515 vcm.n1003 vcm.n1002 0.0466957
R22516 vcm.n1003 vcm.n955 0.0466957
R22517 vcm.n1074 vcm.n1026 0.0466957
R22518 vcm.n1074 vcm.n1073 0.0466957
R22519 vcm.n1052 vcm.n1051 0.0466957
R22520 vcm.n1052 vcm.n1028 0.0466957
R22521 vcm.n1063 vcm.n1062 0.0466957
R22522 vcm.n1063 vcm.n1027 0.0466957
R22523 vcm.n1162 vcm.n1161 0.0466957
R22524 vcm.n1149 vcm.n1101 0.0466957
R22525 vcm.n1149 vcm.n1148 0.0466957
R22526 vcm.n1106 vcm.n1105 0.0466957
R22527 vcm.n1116 vcm.n1115 0.0466957
R22528 vcm.n1116 vcm.n1104 0.0466957
R22529 vcm.n1127 vcm.n1126 0.0466957
R22530 vcm.n1127 vcm.n1103 0.0466957
R22531 vcm.n1138 vcm.n1137 0.0466957
R22532 vcm.n1138 vcm.n1102 0.0466957
R22533 vcm.n777 vcm.n740 0.0466957
R22534 vcm.n777 vcm.n776 0.0466957
R22535 vcm.n769 vcm.n742 0.0466957
R22536 vcm.n769 vcm.n768 0.0466957
R22537 vcm.n745 vcm.n744 0.0466957
R22538 vcm.n760 vcm.n759 0.0466957
R22539 vcm.n760 vcm.n743 0.0466957
R22540 vcm.n829 vcm.n814 0.0466957
R22541 vcm.n829 vcm.n828 0.0466957
R22542 vcm.n816 vcm.n815 0.0466957
R22543 vcm.n911 vcm.n910 0.0466957
R22544 vcm.n911 vcm.n902 0.0466957
R22545 vcm.n919 vcm.n918 0.0466957
R22546 vcm.n919 vcm.n901 0.0466957
R22547 vcm.n984 vcm.n960 0.0466957
R22548 vcm.n984 vcm.n983 0.0466957
R22549 vcm.n963 vcm.n962 0.0466957
R22550 vcm.n973 vcm.n972 0.0466957
R22551 vcm.n973 vcm.n961 0.0466957
R22552 vcm.n1044 vcm.n1032 0.0466957
R22553 vcm.n1044 vcm.n1043 0.0466957
R22554 vcm.n1034 vcm.n1033 0.0466957
R22555 vcm.n40 vcm.n36 0.0466957
R22556 vcm.n40 vcm.n39 0.0466957
R22557 vcm.n15 vcm.n14 0.0466957
R22558 vcm.n29 vcm.n28 0.0466957
R22559 vcm.n29 vcm.n6 0.0466957
R22560 vcm.n76 vcm.n75 0.0466957
R22561 vcm.n76 vcm.n72 0.0466957
R22562 vcm.n63 vcm.n62 0.0466957
R22563 vcm.n63 vcm.n2 0.0466957
R22564 vcm.n107 vcm.n106 0.0466957
R22565 vcm.n107 vcm.n103 0.0466957
R22566 vcm.n559 vcm.n498 0.0394617
R22567 vcm.n425 vcm.n424 0.0394617
R22568 vcm.n147 vcm.n146 0.0394617
R22569 vcm.n264 vcm.n263 0.0394617
R22570 vcm.n281 vcm.n280 0.0394617
R22571 vcm.n878 vcm.n802 0.0394617
R22572 vcm.n1176 vcm.n1175 0.0385543
R22573 vcm.n654 vcm.n653 0.0385543
R22574 vcm.n490 vcm.n489 0.0385543
R22575 vcm.n1022 vcm.n1021 0.0385543
R22576 vcm.n943 vcm.n942 0.0385543
R22577 vcm.n794 vcm.n793 0.0385543
R22578 vcm.n1014 vcm.n1013 0.0385543
R22579 vcm.n1159 vcm.n1158 0.0385543
R22580 vcm.n1188 vcm.n122 0.0385543
R22581 vcm.n754 vcm.n753 0.0302414
R22582 vcm.n11 vcm.n10 0.0270767
R22583 vcm.n906 vcm.n905 0.0270767
R22584 vcm.n289 vcm.n288 0.0270767
R22585 vcm.n362 vcm.n361 0.0270767
R22586 vcm.n154 vcm.n153 0.0270767
R22587 vcm.n213 vcm.n212 0.0270767
R22588 vcm.n451 vcm.n450 0.0270767
R22589 vcm.n508 vcm.n507 0.0270767
R22590 vcm.n597 vcm.n596 0.0270767
R22591 vcm.n672 vcm.n671 0.0270767
R22592 vcm.n1108 vcm.n1107 0.0270767
R22593 vcm.n747 vcm.n746 0.0270767
R22594 vcm.n818 vcm.n817 0.0270767
R22595 vcm.n965 vcm.n964 0.0270767
R22596 vcm.n1036 vcm.n1035 0.0270767
R22597 vcm.n17 vcm.n16 0.0270767
R22598 vcm.n100 vcm 0.0209545
R22599 vcm.n88 vcm 0.0209545
R22600 vcm.n54 vcm 0.0209545
R22601 vcm.n376 vcm 0.0209545
R22602 vcm.n483 vcm 0.0209545
R22603 vcm.n257 vcm 0.0209545
R22604 vcm.n181 vcm 0.0209545
R22605 vcm.n235 vcm 0.0209545
R22606 vcm.n224 vcm 0.0209545
R22607 vcm.n163 vcm 0.0209545
R22608 vcm.n172 vcm 0.0209545
R22609 vcm.n246 vcm 0.0209545
R22610 vcm.n190 vcm 0.0209545
R22611 vcm.n311 vcm 0.0209545
R22612 vcm.n322 vcm 0.0209545
R22613 vcm.n333 vcm 0.0209545
R22614 vcm.n418 vcm 0.0209545
R22615 vcm.n404 vcm 0.0209545
R22616 vcm.n475 vcm 0.0209545
R22617 vcm.n467 vcm 0.0209545
R22618 vcm.n459 vcm 0.0209545
R22619 vcm.n530 vcm 0.0209545
R22620 vcm.n519 vcm 0.0209545
R22621 vcm.n300 vcm 0.0209545
R22622 vcm.n390 vcm 0.0209545
R22623 vcm.n541 vcm 0.0209545
R22624 vcm.n552 vcm 0.0209545
R22625 vcm.n709 vcm 0.0209545
R22626 vcm.n647 vcm 0.0209545
R22627 vcm.n633 vcm 0.0209545
R22628 vcm.n701 vcm 0.0209545
R22629 vcm.n692 vcm 0.0209545
R22630 vcm.n625 vcm 0.0209545
R22631 vcm.n611 vcm 0.0209545
R22632 vcm.n684 vcm 0.0209545
R22633 vcm.n930 vcm 0.0209545
R22634 vcm.n938 vcm 0.0209545
R22635 vcm.n788 vcm 0.0209545
R22636 vcm.n840 vcm 0.0209545
R22637 vcm.n854 vcm 0.0209545
R22638 vcm.n868 vcm 0.0209545
R22639 vcm.n995 vcm 0.0209545
R22640 vcm.n1006 vcm 0.0209545
R22641 vcm.n1077 vcm 0.0209545
R22642 vcm.n1055 vcm 0.0209545
R22643 vcm.n1066 vcm 0.0209545
R22644 vcm.n1152 vcm 0.0209545
R22645 vcm.n1119 vcm 0.0209545
R22646 vcm.n1130 vcm 0.0209545
R22647 vcm.n1141 vcm 0.0209545
R22648 vcm.n780 vcm 0.0209545
R22649 vcm.n772 vcm 0.0209545
R22650 vcm.n763 vcm 0.0209545
R22651 vcm.n832 vcm 0.0209545
R22652 vcm.n914 vcm 0.0209545
R22653 vcm.n922 vcm 0.0209545
R22654 vcm.n987 vcm 0.0209545
R22655 vcm.n976 vcm 0.0209545
R22656 vcm.n1047 vcm 0.0209545
R22657 vcm.n42 vcm 0.0209545
R22658 vcm.n31 vcm 0.0209545
R22659 vcm.n78 vcm 0.0209545
R22660 vcm.n65 vcm 0.0209545
R22661 vcm.n109 vcm 0.0209545
R22662 vcm.n753 vcm.n750 0.0197903
R22663 vcm vcm.n99 0.0150455
R22664 vcm vcm.n87 0.0150455
R22665 vcm vcm.n53 0.0150455
R22666 vcm.n374 vcm 0.0150455
R22667 vcm.n481 vcm 0.0150455
R22668 vcm.n255 vcm 0.0150455
R22669 vcm.n179 vcm 0.0150455
R22670 vcm.n233 vcm 0.0150455
R22671 vcm.n222 vcm 0.0150455
R22672 vcm.n161 vcm 0.0150455
R22673 vcm.n170 vcm 0.0150455
R22674 vcm.n244 vcm 0.0150455
R22675 vcm.n188 vcm 0.0150455
R22676 vcm.n309 vcm 0.0150455
R22677 vcm.n320 vcm 0.0150455
R22678 vcm.n331 vcm 0.0150455
R22679 vcm.n416 vcm 0.0150455
R22680 vcm.n402 vcm 0.0150455
R22681 vcm.n473 vcm 0.0150455
R22682 vcm.n465 vcm 0.0150455
R22683 vcm.n457 vcm 0.0150455
R22684 vcm.n528 vcm 0.0150455
R22685 vcm.n517 vcm 0.0150455
R22686 vcm.n298 vcm 0.0150455
R22687 vcm.n388 vcm 0.0150455
R22688 vcm.n539 vcm 0.0150455
R22689 vcm.n550 vcm 0.0150455
R22690 vcm.n707 vcm 0.0150455
R22691 vcm.n645 vcm 0.0150455
R22692 vcm.n631 vcm 0.0150455
R22693 vcm.n699 vcm 0.0150455
R22694 vcm.n690 vcm 0.0150455
R22695 vcm.n623 vcm 0.0150455
R22696 vcm.n609 vcm 0.0150455
R22697 vcm.n682 vcm 0.0150455
R22698 vcm.n928 vcm 0.0150455
R22699 vcm.n936 vcm 0.0150455
R22700 vcm.n786 vcm 0.0150455
R22701 vcm.n838 vcm 0.0150455
R22702 vcm.n852 vcm 0.0150455
R22703 vcm.n866 vcm 0.0150455
R22704 vcm.n993 vcm 0.0150455
R22705 vcm.n1004 vcm 0.0150455
R22706 vcm.n1075 vcm 0.0150455
R22707 vcm.n1053 vcm 0.0150455
R22708 vcm.n1064 vcm 0.0150455
R22709 vcm.n1150 vcm 0.0150455
R22710 vcm.n1117 vcm 0.0150455
R22711 vcm.n1128 vcm 0.0150455
R22712 vcm.n1139 vcm 0.0150455
R22713 vcm.n778 vcm 0.0150455
R22714 vcm.n770 vcm 0.0150455
R22715 vcm.n761 vcm 0.0150455
R22716 vcm.n830 vcm 0.0150455
R22717 vcm.n912 vcm 0.0150455
R22718 vcm.n920 vcm 0.0150455
R22719 vcm.n985 vcm 0.0150455
R22720 vcm.n974 vcm 0.0150455
R22721 vcm.n1045 vcm 0.0150455
R22722 vcm vcm.n41 0.0150455
R22723 vcm vcm.n30 0.0150455
R22724 vcm vcm.n77 0.0150455
R22725 vcm vcm.n64 0.0150455
R22726 vcm vcm.n108 0.0150455
R22727 vcm.n753 vcm.n752 0.00833208
R22728 vcm vcm 0.00640909
R22729 vcm vcm 0.00640909
R22730 vcm vcm 0.00640909
R22731 vcm vcm 0.00640909
R22732 vcm vcm 0.00640909
R22733 vcm vcm 0.00640909
R22734 vcm vcm 0.00640909
R22735 vcm vcm 0.00640909
R22736 vcm vcm 0.00640909
R22737 vcm vcm 0.00640909
R22738 vcm vcm 0.00640909
R22739 vcm vcm 0.00640909
R22740 vcm vcm 0.00640909
R22741 vcm vcm 0.00640909
R22742 vcm vcm 0.00640909
R22743 vcm vcm 0.00640909
R22744 vcm vcm 0.00640909
R22745 vcm vcm 0.00640909
R22746 vcm vcm 0.00640909
R22747 vcm vcm 0.00640909
R22748 vcm vcm 0.00640909
R22749 vcm vcm 0.00640909
R22750 vcm vcm 0.00640909
R22751 vcm vcm 0.00640909
R22752 vcm vcm 0.00640909
R22753 vcm vcm 0.00640909
R22754 vcm vcm 0.00640909
R22755 vcm vcm 0.00640909
R22756 vcm vcm 0.00640909
R22757 vcm vcm 0.00640909
R22758 vcm vcm 0.00640909
R22759 vcm vcm 0.00640909
R22760 vcm vcm 0.00640909
R22761 vcm vcm 0.00640909
R22762 vcm vcm 0.00640909
R22763 vcm vcm 0.00640909
R22764 vcm vcm 0.00640909
R22765 vcm vcm 0.00640909
R22766 vcm vcm 0.00640909
R22767 vcm vcm 0.00640909
R22768 vcm vcm 0.00640909
R22769 vcm vcm 0.00640909
R22770 vcm vcm 0.00640909
R22771 vcm vcm 0.00640909
R22772 vcm vcm 0.00640909
R22773 vcm vcm 0.00640909
R22774 vcm vcm 0.00640909
R22775 vcm vcm 0.00640909
R22776 vcm vcm 0.00640909
R22777 vcm vcm 0.00640909
R22778 vcm vcm 0.00640909
R22779 vcm vcm 0.00640909
R22780 vcm vcm 0.00640909
R22781 vcm vcm 0.00640909
R22782 vcm vcm 0.00640909
R22783 vcm vcm 0.00640909
R22784 vcm vcm 0.00640909
R22785 vcm vcm 0.00640909
R22786 vcm vcm 0.00640909
R22787 vcm vcm 0.00640909
R22788 vcm vcm 0.00640909
R22789 vcm vcm 0.00640909
R22790 vcm vcm 0.00640909
R22791 vcm vcm 0.00640909
R22792 vcm.n756 vcm.n755 0.00570833
R22793 vcm.n754 vcm.n749 0.00481034
R22794 vcm.n1174 vcm.n1173 0.00321739
R22795 vcm.n101 vcm.n0 0.00321739
R22796 vcm.n97 vcm.n96 0.00321739
R22797 vcm.n89 vcm.n70 0.00321739
R22798 vcm.n85 vcm.n84 0.00321739
R22799 vcm.n55 vcm.n4 0.00321739
R22800 vcm.n51 vcm.n50 0.00321739
R22801 vcm.n12 vcm.n9 0.00321739
R22802 vcm.n907 vcm.n904 0.00321739
R22803 vcm.n651 vcm.n650 0.00321739
R22804 vcm.n558 vcm.n500 0.00321739
R22805 vcm.n290 vcm.n287 0.00321739
R22806 vcm.n377 vcm.n358 0.00321739
R22807 vcm.n372 vcm.n371 0.00321739
R22808 vcm.n363 vcm.n360 0.00321739
R22809 vcm.n488 vcm.n487 0.00321739
R22810 vcm.n484 vcm.n444 0.00321739
R22811 vcm.n479 vcm.n478 0.00321739
R22812 vcm.n422 vcm.n421 0.00321739
R22813 vcm.n195 vcm.n194 0.00321739
R22814 vcm.n266 vcm.n265 0.00321739
R22815 vcm.n258 vcm.n206 0.00321739
R22816 vcm.n253 vcm.n252 0.00321739
R22817 vcm.n182 vcm.n149 0.00321739
R22818 vcm.n177 vcm.n176 0.00321739
R22819 vcm.n236 vcm.n208 0.00321739
R22820 vcm.n231 vcm.n230 0.00321739
R22821 vcm.n225 vcm.n209 0.00321739
R22822 vcm.n220 vcm.n219 0.00321739
R22823 vcm.n214 vcm.n211 0.00321739
R22824 vcm.n159 vcm.n158 0.00321739
R22825 vcm.n164 vcm.n151 0.00321739
R22826 vcm.n168 vcm.n167 0.00321739
R22827 vcm.n173 vcm.n150 0.00321739
R22828 vcm.n242 vcm.n241 0.00321739
R22829 vcm.n247 vcm.n207 0.00321739
R22830 vcm.n186 vcm.n185 0.00321739
R22831 vcm.n191 vcm.n148 0.00321739
R22832 vcm.n340 vcm.n339 0.00321739
R22833 vcm.n307 vcm.n306 0.00321739
R22834 vcm.n312 vcm.n284 0.00321739
R22835 vcm.n318 vcm.n317 0.00321739
R22836 vcm.n323 vcm.n283 0.00321739
R22837 vcm.n329 vcm.n328 0.00321739
R22838 vcm.n334 vcm.n282 0.00321739
R22839 vcm.n419 vcm.n355 0.00321739
R22840 vcm.n414 vcm.n413 0.00321739
R22841 vcm.n400 vcm.n399 0.00321739
R22842 vcm.n405 vcm.n356 0.00321739
R22843 vcm.n476 vcm.n445 0.00321739
R22844 vcm.n471 vcm.n470 0.00321739
R22845 vcm.n468 vcm.n446 0.00321739
R22846 vcm.n463 vcm.n462 0.00321739
R22847 vcm.n460 vcm.n447 0.00321739
R22848 vcm.n455 vcm.n454 0.00321739
R22849 vcm.n452 vcm.n449 0.00321739
R22850 vcm.n531 vcm.n503 0.00321739
R22851 vcm.n526 vcm.n525 0.00321739
R22852 vcm.n520 vcm.n504 0.00321739
R22853 vcm.n515 vcm.n514 0.00321739
R22854 vcm.n509 vcm.n506 0.00321739
R22855 vcm.n296 vcm.n295 0.00321739
R22856 vcm.n301 vcm.n285 0.00321739
R22857 vcm.n386 vcm.n385 0.00321739
R22858 vcm.n391 vcm.n357 0.00321739
R22859 vcm.n537 vcm.n536 0.00321739
R22860 vcm.n542 vcm.n502 0.00321739
R22861 vcm.n548 vcm.n547 0.00321739
R22862 vcm.n553 vcm.n501 0.00321739
R22863 vcm.n714 vcm.n713 0.00321739
R22864 vcm.n705 vcm.n704 0.00321739
R22865 vcm.n710 vcm.n663 0.00321739
R22866 vcm.n648 vcm.n584 0.00321739
R22867 vcm.n643 vcm.n642 0.00321739
R22868 vcm.n629 vcm.n628 0.00321739
R22869 vcm.n634 vcm.n585 0.00321739
R22870 vcm.n702 vcm.n665 0.00321739
R22871 vcm.n697 vcm.n696 0.00321739
R22872 vcm.n688 vcm.n687 0.00321739
R22873 vcm.n693 vcm.n666 0.00321739
R22874 vcm.n626 vcm.n592 0.00321739
R22875 vcm.n621 vcm.n620 0.00321739
R22876 vcm.n598 vcm.n595 0.00321739
R22877 vcm.n607 vcm.n606 0.00321739
R22878 vcm.n612 vcm.n593 0.00321739
R22879 vcm.n685 vcm.n668 0.00321739
R22880 vcm.n680 vcm.n679 0.00321739
R22881 vcm.n673 vcm.n670 0.00321739
R22882 vcm.n1081 vcm.n1080 0.00321739
R22883 vcm.n941 vcm.n898 0.00321739
R22884 vcm.n926 vcm.n925 0.00321739
R22885 vcm.n931 vcm.n900 0.00321739
R22886 vcm.n934 vcm.n933 0.00321739
R22887 vcm.n939 vcm.n899 0.00321739
R22888 vcm.n792 vcm.n737 0.00321739
R22889 vcm.n784 vcm.n783 0.00321739
R22890 vcm.n789 vcm.n738 0.00321739
R22891 vcm.n877 vcm.n804 0.00321739
R22892 vcm.n836 vcm.n835 0.00321739
R22893 vcm.n841 vcm.n807 0.00321739
R22894 vcm.n850 vcm.n849 0.00321739
R22895 vcm.n855 vcm.n806 0.00321739
R22896 vcm.n864 vcm.n863 0.00321739
R22897 vcm.n869 vcm.n805 0.00321739
R22898 vcm.n1012 vcm.n954 0.00321739
R22899 vcm.n991 vcm.n990 0.00321739
R22900 vcm.n996 vcm.n956 0.00321739
R22901 vcm.n1002 vcm.n1001 0.00321739
R22902 vcm.n1007 vcm.n955 0.00321739
R22903 vcm.n1078 vcm.n1026 0.00321739
R22904 vcm.n1073 vcm.n1072 0.00321739
R22905 vcm.n1051 vcm.n1050 0.00321739
R22906 vcm.n1056 vcm.n1028 0.00321739
R22907 vcm.n1062 vcm.n1061 0.00321739
R22908 vcm.n1067 vcm.n1027 0.00321739
R22909 vcm.n1161 vcm.n1160 0.00321739
R22910 vcm.n1153 vcm.n1101 0.00321739
R22911 vcm.n1148 vcm.n1147 0.00321739
R22912 vcm.n1109 vcm.n1106 0.00321739
R22913 vcm.n1115 vcm.n1114 0.00321739
R22914 vcm.n1120 vcm.n1104 0.00321739
R22915 vcm.n1126 vcm.n1125 0.00321739
R22916 vcm.n1131 vcm.n1103 0.00321739
R22917 vcm.n1137 vcm.n1136 0.00321739
R22918 vcm.n1142 vcm.n1102 0.00321739
R22919 vcm.n781 vcm.n740 0.00321739
R22920 vcm.n776 vcm.n775 0.00321739
R22921 vcm.n773 vcm.n742 0.00321739
R22922 vcm.n768 vcm.n767 0.00321739
R22923 vcm.n748 vcm.n745 0.00321739
R22924 vcm.n759 vcm.n758 0.00321739
R22925 vcm.n764 vcm.n743 0.00321739
R22926 vcm.n833 vcm.n814 0.00321739
R22927 vcm.n828 vcm.n827 0.00321739
R22928 vcm.n819 vcm.n816 0.00321739
R22929 vcm.n910 vcm.n909 0.00321739
R22930 vcm.n915 vcm.n902 0.00321739
R22931 vcm.n918 vcm.n917 0.00321739
R22932 vcm.n923 vcm.n901 0.00321739
R22933 vcm.n988 vcm.n960 0.00321739
R22934 vcm.n983 vcm.n982 0.00321739
R22935 vcm.n966 vcm.n963 0.00321739
R22936 vcm.n972 vcm.n971 0.00321739
R22937 vcm.n977 vcm.n961 0.00321739
R22938 vcm.n1048 vcm.n1032 0.00321739
R22939 vcm.n1043 vcm.n1042 0.00321739
R22940 vcm.n1037 vcm.n1034 0.00321739
R22941 vcm.n43 vcm.n36 0.00321739
R22942 vcm.n39 vcm.n38 0.00321739
R22943 vcm.n18 vcm.n15 0.00321739
R22944 vcm.n28 vcm.n27 0.00321739
R22945 vcm.n32 vcm.n6 0.00321739
R22946 vcm.n75 vcm.n74 0.00321739
R22947 vcm.n79 vcm.n72 0.00321739
R22948 vcm.n62 vcm.n61 0.00321739
R22949 vcm.n66 vcm.n2 0.00321739
R22950 vcm.n106 vcm.n105 0.00321739
R22951 vcm.n110 vcm.n103 0.00321739
R22952 vcm.n121 vcm.n120 0.00321739
R22953 vcm.n99 vcm.n1 0.00239652
R22954 vcm.n87 vcm.n71 0.00239652
R22955 vcm.n53 vcm.n5 0.00239652
R22956 vcm.n41 vcm.n37 0.00239652
R22957 vcm.n30 vcm.n7 0.00239652
R22958 vcm.n77 vcm.n73 0.00239652
R22959 vcm.n64 vcm.n3 0.00239652
R22960 vcm.n108 vcm.n104 0.00239652
R22961 vcm.n257 vcm.n256 0.00239442
R22962 vcm.n322 vcm.n321 0.00239442
R22963 vcm.n459 vcm.n458 0.00239442
R22964 vcm.n390 vcm.n389 0.00239442
R22965 vcm.n788 vcm.n787 0.00239442
R22966 vcm.n854 vcm.n853 0.00239442
R22967 vcm.n922 vcm.n921 0.00239442
R22968 vcm.n976 vcm.n975 0.00239442
R22969 vcm.n376 vcm.n375 0.00225049
R22970 vcm.n483 vcm.n482 0.00225049
R22971 vcm.n181 vcm.n180 0.00225049
R22972 vcm.n235 vcm.n234 0.00225049
R22973 vcm.n224 vcm.n223 0.00225049
R22974 vcm.n163 vcm.n162 0.00225049
R22975 vcm.n172 vcm.n171 0.00225049
R22976 vcm.n246 vcm.n245 0.00225049
R22977 vcm.n190 vcm.n189 0.00225049
R22978 vcm.n311 vcm.n310 0.00225049
R22979 vcm.n333 vcm.n332 0.00225049
R22980 vcm.n418 vcm.n417 0.00225049
R22981 vcm.n404 vcm.n403 0.00225049
R22982 vcm.n475 vcm.n474 0.00225049
R22983 vcm.n467 vcm.n466 0.00225049
R22984 vcm.n530 vcm.n529 0.00225049
R22985 vcm.n519 vcm.n518 0.00225049
R22986 vcm.n300 vcm.n299 0.00225049
R22987 vcm.n541 vcm.n540 0.00225049
R22988 vcm.n552 vcm.n551 0.00225049
R22989 vcm.n709 vcm.n708 0.00225049
R22990 vcm.n647 vcm.n646 0.00225049
R22991 vcm.n633 vcm.n632 0.00225049
R22992 vcm.n701 vcm.n700 0.00225049
R22993 vcm.n692 vcm.n691 0.00225049
R22994 vcm.n625 vcm.n624 0.00225049
R22995 vcm.n611 vcm.n610 0.00225049
R22996 vcm.n684 vcm.n683 0.00225049
R22997 vcm.n930 vcm.n929 0.00225049
R22998 vcm.n938 vcm.n937 0.00225049
R22999 vcm.n840 vcm.n839 0.00225049
R23000 vcm.n868 vcm.n867 0.00225049
R23001 vcm.n995 vcm.n994 0.00225049
R23002 vcm.n1006 vcm.n1005 0.00225049
R23003 vcm.n1077 vcm.n1076 0.00225049
R23004 vcm.n1055 vcm.n1054 0.00225049
R23005 vcm.n1066 vcm.n1065 0.00225049
R23006 vcm.n1152 vcm.n1151 0.00225049
R23007 vcm.n1119 vcm.n1118 0.00225049
R23008 vcm.n1130 vcm.n1129 0.00225049
R23009 vcm.n1141 vcm.n1140 0.00225049
R23010 vcm.n780 vcm.n779 0.00225049
R23011 vcm.n772 vcm.n771 0.00225049
R23012 vcm.n763 vcm.n762 0.00225049
R23013 vcm.n832 vcm.n831 0.00225049
R23014 vcm.n914 vcm.n913 0.00225049
R23015 vcm.n987 vcm.n986 0.00225049
R23016 vcm.n1047 vcm.n1046 0.00225049
R23017 vcm.n261 vcm.n260 0.00149648
R23018 vcm.n337 vcm.n336 0.00149648
R23019 vcm.n354 vcm.n353 0.00149648
R23020 vcm.n411 vcm.n410 0.00149648
R23021 vcm.n408 vcm.n407 0.00149648
R23022 vcm.n512 vcm.n511 0.00149648
R23023 vcm.n397 vcm.n396 0.00149648
R23024 vcm.n394 vcm.n393 0.00149648
R23025 vcm.n556 vcm.n555 0.00149648
R23026 vcm.n583 vcm.n582 0.00149648
R23027 vcm.n640 vcm.n639 0.00149648
R23028 vcm.n637 vcm.n636 0.00149648
R23029 vcm.n591 vcm.n590 0.00149648
R23030 vcm.n618 vcm.n617 0.00149648
R23031 vcm.n615 vcm.n614 0.00149648
R23032 vcm.n601 vcm.n600 0.00149648
R23033 vcm.n1070 vcm.n1069 0.00149648
R23034 vcm.n999 vcm.n998 0.00149648
R23035 vcm.n858 vcm.n857 0.00149648
R23036 vcm.n825 vcm.n824 0.00149648
R23037 vcm.n822 vcm.n821 0.00149648
R23038 vcm.n844 vcm.n843 0.00149648
R23039 vcm.n959 vcm.n958 0.00149648
R23040 vcm.n980 vcm.n979 0.00149648
R23041 vcm.n1031 vcm.n1030 0.00149648
R23042 vcm.n260 vcm.n259 0.00149647
R23043 vcm.n336 vcm.n335 0.00149647
R23044 vcm.n353 vcm.n352 0.00149647
R23045 vcm.n410 vcm.n409 0.00149647
R23046 vcm.n407 vcm.n406 0.00149647
R23047 vcm.n511 vcm.n510 0.00149647
R23048 vcm.n396 vcm.n395 0.00149647
R23049 vcm.n393 vcm.n392 0.00149647
R23050 vcm.n555 vcm.n554 0.00149647
R23051 vcm.n582 vcm.n581 0.00149647
R23052 vcm.n639 vcm.n638 0.00149647
R23053 vcm.n636 vcm.n635 0.00149647
R23054 vcm.n590 vcm.n589 0.00149647
R23055 vcm.n617 vcm.n616 0.00149647
R23056 vcm.n614 vcm.n613 0.00149647
R23057 vcm.n600 vcm.n599 0.00149647
R23058 vcm.n1069 vcm.n1068 0.00149647
R23059 vcm.n998 vcm.n997 0.00149647
R23060 vcm.n857 vcm.n856 0.00149647
R23061 vcm.n824 vcm.n823 0.00149647
R23062 vcm.n821 vcm.n820 0.00149647
R23063 vcm.n843 vcm.n842 0.00149647
R23064 vcm.n958 vcm.n957 0.00149647
R23065 vcm.n979 vcm.n978 0.00149647
R23066 vcm.n1030 vcm.n1029 0.00149647
R23067 vcm.n239 vcm.n238 0.00145928
R23068 vcm.n293 vcm.n292 0.00145928
R23069 vcm.n383 vcm.n382 0.00145928
R23070 vcm.n872 vcm.n871 0.00145928
R23071 vcm.n1025 vcm.n1024 0.00145928
R23072 vcm.n813 vcm.n812 0.00145928
R23073 vcm.n1112 vcm.n1111 0.00145928
R23074 vcm.n25 vcm.n24 0.00145928
R23075 vcm.n46 vcm.n45 0.00145928
R23076 vcm.n59 vcm.n58 0.00145928
R23077 vcm.n92 vcm.n91 0.00145928
R23078 vcm.n117 vcm.n116 0.00145928
R23079 vcm.n238 vcm.n237 0.00139285
R23080 vcm.n292 vcm.n291 0.00139285
R23081 vcm.n382 vcm.n381 0.00139285
R23082 vcm.n871 vcm.n870 0.00139285
R23083 vcm.n1024 vcm.n1023 0.00139285
R23084 vcm.n812 vcm.n811 0.00139285
R23085 vcm.n1111 vcm.n1110 0.00139285
R23086 vcm.n24 vcm.n23 0.00139285
R23087 vcm.n45 vcm.n44 0.00139285
R23088 vcm.n58 vcm.n57 0.00139285
R23089 vcm.n91 vcm.n90 0.00139285
R23090 vcm.n116 vcm.n115 0.00139285
R23091 vcm.n145 vcm.n143 0.00114214
R23092 vcm.n888 vcm.n887 0.00104325
R23093 vcm.n435 vcm.n434 0.00104325
R23094 vcm.n569 vcm.n568 0.00104325
R23095 vcm.n726 vcm.n725 0.00104325
R23096 vcm.n659 vcm.n577 0.00103325
R23097 vcm.n495 vcm.n443 0.00103325
R23098 vcm.n346 vcm.n279 0.00103325
R23099 vcm.n1093 vcm.n1092 0.00103325
R23100 vcm.n948 vcm.n896 0.00103325
R23101 vcm.n799 vcm.n735 0.00103325
R23102 vcm.n1167 vcm.n1100 0.00103325
R23103 vcm.n799 vcm.n798 0.00103325
R23104 vcm.n948 vcm.n947 0.00103325
R23105 vcm.n1019 vcm.n1018 0.00103325
R23106 vcm.n1167 vcm.n1166 0.00103325
R23107 vcm.n1181 vcm.n1180 0.00103325
R23108 vcm.n272 vcm.n271 0.00103325
R23109 vcm.n346 vcm.n345 0.00103325
R23110 vcm.n495 vcm.n494 0.00103325
R23111 vcm.n659 vcm.n658 0.00103325
R23112 vcm.n568 vcm.n567 0.00103323
R23113 vcm.n434 vcm.n433 0.00103323
R23114 vcm.n142 vcm.n141 0.00103323
R23115 vcm.n725 vcm.n724 0.00103323
R23116 vcm.n887 vcm.n886 0.00103323
R23117 vcm.n1171 vcm.n1169 0.00103319
R23118 vcm.n1097 vcm.n1095 0.00103319
R23119 vcm.n1089 vcm.n1087 0.00103319
R23120 vcm.n952 vcm.n950 0.00103319
R23121 vcm.n893 vcm.n891 0.00103319
R23122 vcm.n732 vcm.n730 0.00103319
R23123 vcm.n574 vcm.n572 0.00103319
R23124 vcm.n440 vcm.n438 0.00103319
R23125 vcm.n276 vcm.n274 0.00103319
R23126 vcm.n205 vcm.n203 0.00103319
R23127 vcm.n1182 vcm.n1171 0.00103319
R23128 vcm.n1168 vcm.n1097 0.00103319
R23129 vcm.n1094 vcm.n1089 0.00103319
R23130 vcm.n1020 vcm.n952 0.00103319
R23131 vcm.n949 vcm.n893 0.00103319
R23132 vcm.n800 vcm.n732 0.00103319
R23133 vcm.n660 vcm.n574 0.00103319
R23134 vcm.n496 vcm.n440 0.00103319
R23135 vcm.n347 vcm.n276 0.00103319
R23136 vcm.n273 vcm.n205 0.00103319
R23137 vcm.n128 vcm.n127 0.00103293
R23138 vcm.n202 vcm.n145 0.00103293
R23139 vcm.n201 vcm.n200 0.00102352
R23140 vcm.n883 vcm.n882 0.00102352
R23141 vcm.n430 vcm.n429 0.00102352
R23142 vcm.n564 vcm.n563 0.00102352
R23143 vcm.n721 vcm.n720 0.00102352
R23144 vcm.n890 vcm.n889 0.00102346
R23145 vcm.n437 vcm.n436 0.00102346
R23146 vcm.n571 vcm.n570 0.00102346
R23147 vcm.n728 vcm.n727 0.00102346
R23148 vcm.n889 vcm.n888 0.00101835
R23149 vcm.n727 vcm.n726 0.00101835
R23150 vcm.n570 vcm.n569 0.00101835
R23151 vcm.n436 vcm.n435 0.00101835
R23152 vcm.n890 vcm.n883 0.0010183
R23153 vcm.n728 vcm.n721 0.0010183
R23154 vcm.n571 vcm.n564 0.0010183
R23155 vcm.n437 vcm.n430 0.0010183
R23156 vcm.n202 vcm.n201 0.0010183
R23157 vcm.n125 vcm.n124 0.00100588
R23158 vcm.n131 vcm.n130 0.00100116
R23159 vcm.n576 vcm.n575 0.00100116
R23160 vcm.n566 vcm.n565 0.00100116
R23161 vcm.n442 vcm.n441 0.00100116
R23162 vcm.n432 vcm.n431 0.00100116
R23163 vcm.n140 vcm.n139 0.00100116
R23164 vcm.n137 vcm.n136 0.00100116
R23165 vcm.n278 vcm.n277 0.00100116
R23166 vcm.n723 vcm.n722 0.00100116
R23167 vcm.n1091 vcm.n1090 0.00100116
R23168 vcm.n895 vcm.n894 0.00100116
R23169 vcm.n734 vcm.n733 0.00100116
R23170 vcm.n885 vcm.n884 0.00100116
R23171 vcm.n134 vcm.n133 0.00100116
R23172 vcm.n1099 vcm.n1098 0.00100116
R23173 vcm.n127 vcm.n126 0.00100034
R23174 vcm.n145 vcm.n144 0.00100034
R23175 vcm.n256 vcm.n255 0.0010003
R23176 vcm.n321 vcm.n320 0.0010003
R23177 vcm.n458 vcm.n457 0.0010003
R23178 vcm.n389 vcm.n388 0.0010003
R23179 vcm.n787 vcm.n786 0.0010003
R23180 vcm.n853 vcm.n852 0.0010003
R23181 vcm.n921 vcm.n920 0.0010003
R23182 vcm.n975 vcm.n974 0.0010003
R23183 vcm.n375 vcm.n374 0.00100024
R23184 vcm.n482 vcm.n481 0.00100024
R23185 vcm.n180 vcm.n179 0.00100024
R23186 vcm.n234 vcm.n233 0.00100024
R23187 vcm.n223 vcm.n222 0.00100024
R23188 vcm.n162 vcm.n161 0.00100024
R23189 vcm.n171 vcm.n170 0.00100024
R23190 vcm.n245 vcm.n244 0.00100024
R23191 vcm.n189 vcm.n188 0.00100024
R23192 vcm.n310 vcm.n309 0.00100024
R23193 vcm.n332 vcm.n331 0.00100024
R23194 vcm.n417 vcm.n416 0.00100024
R23195 vcm.n403 vcm.n402 0.00100024
R23196 vcm.n474 vcm.n473 0.00100024
R23197 vcm.n466 vcm.n465 0.00100024
R23198 vcm.n529 vcm.n528 0.00100024
R23199 vcm.n518 vcm.n517 0.00100024
R23200 vcm.n299 vcm.n298 0.00100024
R23201 vcm.n540 vcm.n539 0.00100024
R23202 vcm.n551 vcm.n550 0.00100024
R23203 vcm.n708 vcm.n707 0.00100024
R23204 vcm.n646 vcm.n645 0.00100024
R23205 vcm.n632 vcm.n631 0.00100024
R23206 vcm.n700 vcm.n699 0.00100024
R23207 vcm.n691 vcm.n690 0.00100024
R23208 vcm.n624 vcm.n623 0.00100024
R23209 vcm.n610 vcm.n609 0.00100024
R23210 vcm.n683 vcm.n682 0.00100024
R23211 vcm.n929 vcm.n928 0.00100024
R23212 vcm.n937 vcm.n936 0.00100024
R23213 vcm.n839 vcm.n838 0.00100024
R23214 vcm.n867 vcm.n866 0.00100024
R23215 vcm.n994 vcm.n993 0.00100024
R23216 vcm.n1005 vcm.n1004 0.00100024
R23217 vcm.n1076 vcm.n1075 0.00100024
R23218 vcm.n1054 vcm.n1053 0.00100024
R23219 vcm.n1065 vcm.n1064 0.00100024
R23220 vcm.n1151 vcm.n1150 0.00100024
R23221 vcm.n1118 vcm.n1117 0.00100024
R23222 vcm.n1129 vcm.n1128 0.00100024
R23223 vcm.n1140 vcm.n1139 0.00100024
R23224 vcm.n779 vcm.n778 0.00100024
R23225 vcm.n771 vcm.n770 0.00100024
R23226 vcm.n762 vcm.n761 0.00100024
R23227 vcm.n831 vcm.n830 0.00100024
R23228 vcm.n913 vcm.n912 0.00100024
R23229 vcm.n986 vcm.n985 0.00100024
R23230 vcm.n1046 vcm.n1045 0.00100024
R23231 vcm.n100 vcm.n1 0.00100019
R23232 vcm.n88 vcm.n71 0.00100019
R23233 vcm.n54 vcm.n5 0.00100019
R23234 vcm.n42 vcm.n37 0.00100019
R23235 vcm.n31 vcm.n7 0.00100019
R23236 vcm.n78 vcm.n73 0.00100019
R23237 vcm.n65 vcm.n3 0.00100019
R23238 vcm.n109 vcm.n104 0.00100019
R23239 vcm.n675 vcm.n674 0.00100017
R23240 vcm.n1171 vcm.n1170 0.00100008
R23241 vcm.n1097 vcm.n1096 0.00100008
R23242 vcm.n1089 vcm.n1088 0.00100008
R23243 vcm.n952 vcm.n951 0.00100008
R23244 vcm.n893 vcm.n892 0.00100008
R23245 vcm.n732 vcm.n731 0.00100008
R23246 vcm.n574 vcm.n573 0.00100008
R23247 vcm.n440 vcm.n439 0.00100008
R23248 vcm.n276 vcm.n275 0.00100008
R23249 vcm.n205 vcm.n204 0.00100008
R23250 vcm.n143 vcm.n142 0.00100006
R23251 vcm.n1183 vcm.n129 0.00100006
R23252 vcm.n217 vcm.n216 0.00100005
R23253 vcm.n228 vcm.n227 0.00100005
R23254 vcm.n315 vcm.n314 0.00100005
R23255 vcm.n326 vcm.n325 0.00100005
R23256 vcm.n250 vcm.n249 0.00100005
R23257 vcm.n351 vcm.n350 0.00100005
R23258 vcm.n545 vcm.n544 0.00100005
R23259 vcm.n604 vcm.n603 0.00100005
R23260 vcm.n366 vcm.n365 0.00100005
R23261 vcm.n369 vcm.n368 0.00100005
R23262 vcm.n304 vcm.n303 0.00100005
R23263 vcm.n523 vcm.n522 0.00100005
R23264 vcm.n380 vcm.n379 0.00100005
R23265 vcm.n534 vcm.n533 0.00100005
R23266 vcm.n580 vcm.n579 0.00100005
R23267 vcm.n588 vcm.n587 0.00100005
R23268 vcm.n875 vcm.n874 0.00100005
R23269 vcm.n1010 vcm.n1009 0.00100005
R23270 vcm.n1156 vcm.n1155 0.00100005
R23271 vcm.n1145 vcm.n1144 0.00100005
R23272 vcm.n861 vcm.n860 0.00100005
R23273 vcm.n847 vcm.n846 0.00100005
R23274 vcm.n810 vcm.n809 0.00100005
R23275 vcm.n969 vcm.n968 0.00100005
R23276 vcm.n1134 vcm.n1133 0.00100005
R23277 vcm.n1059 vcm.n1058 0.00100005
R23278 vcm.n1123 vcm.n1122 0.00100005
R23279 vcm.n1040 vcm.n1039 0.00100005
R23280 vcm.n21 vcm.n20 0.00100005
R23281 vcm.n82 vcm.n81 0.00100005
R23282 vcm.n113 vcm.n112 0.00100005
R23283 vcm.n48 vcm.n35 0.00100005
R23284 vcm.n94 vcm.n69 0.00100005
R23285 vcm.n1182 vcm.n1181 0.00100005
R23286 vcm.n1168 vcm.n1167 0.00100005
R23287 vcm.n1094 vcm.n1093 0.00100005
R23288 vcm.n1020 vcm.n1019 0.00100005
R23289 vcm.n949 vcm.n948 0.00100005
R23290 vcm.n800 vcm.n799 0.00100005
R23291 vcm.n660 vcm.n659 0.00100005
R23292 vcm.n496 vcm.n495 0.00100005
R23293 vcm.n347 vcm.n346 0.00100005
R23294 vcm.n273 vcm.n272 0.00100005
R23295 vcm.n35 vcm.n34 0.00100004
R23296 vcm.n69 vcm.n68 0.00100004
R23297 vcm.n216 vcm.n215 0.00100004
R23298 vcm.n227 vcm.n226 0.00100004
R23299 vcm.n314 vcm.n313 0.00100004
R23300 vcm.n325 vcm.n324 0.00100004
R23301 vcm.n249 vcm.n248 0.00100004
R23302 vcm.n350 vcm.n349 0.00100004
R23303 vcm.n544 vcm.n543 0.00100004
R23304 vcm.n603 vcm.n602 0.00100004
R23305 vcm.n365 vcm.n364 0.00100004
R23306 vcm.n368 vcm.n367 0.00100004
R23307 vcm.n303 vcm.n302 0.00100004
R23308 vcm.n522 vcm.n521 0.00100004
R23309 vcm.n379 vcm.n378 0.00100004
R23310 vcm.n533 vcm.n532 0.00100004
R23311 vcm.n579 vcm.n578 0.00100004
R23312 vcm.n587 vcm.n586 0.00100004
R23313 vcm.n874 vcm.n873 0.00100004
R23314 vcm.n1009 vcm.n1008 0.00100004
R23315 vcm.n1155 vcm.n1154 0.00100004
R23316 vcm.n1144 vcm.n1143 0.00100004
R23317 vcm.n860 vcm.n859 0.00100004
R23318 vcm.n846 vcm.n845 0.00100004
R23319 vcm.n809 vcm.n808 0.00100004
R23320 vcm.n968 vcm.n967 0.00100004
R23321 vcm.n1133 vcm.n1132 0.00100004
R23322 vcm.n1058 vcm.n1057 0.00100004
R23323 vcm.n1122 vcm.n1121 0.00100004
R23324 vcm.n1039 vcm.n1038 0.00100004
R23325 vcm.n20 vcm.n19 0.00100004
R23326 vcm.n81 vcm.n80 0.00100004
R23327 vcm.n112 vcm.n111 0.00100004
R23328 vcm.n128 vcm.n123 0.000533349
R23329 vcm.n1184 vcm.n128 0.000533349
R23330 vcm.n882 vcm.n801 0.000533349
R23331 vcm.n950 vcm.n135 0.000533349
R23332 vcm.n1087 vcm.n1086 0.000533349
R23333 vcm.n1169 vcm.n132 0.000533349
R23334 vcm.n203 vcm.n138 0.000533349
R23335 vcm.n429 vcm.n348 0.000533349
R23336 vcm.n563 vcm.n497 0.000533349
R23337 vcm.n720 vcm.n661 0.000533349
R23338 vcm.n1184 vcm.n1183 0.000533349
R23339 vcm.n567 vcm.n566 0.00050467
R23340 vcm.n433 vcm.n432 0.00050467
R23341 vcm.n141 vcm.n140 0.00050467
R23342 vcm.n724 vcm.n723 0.00050467
R23343 vcm.n886 vcm.n885 0.00050467
R23344 vcm.n200 vcm.n199 0.00050467
R23345 vcm.n735 vcm.n734 0.00050467
R23346 vcm.n798 vcm.n797 0.00050467
R23347 vcm.n882 vcm.n881 0.00050467
R23348 vcm.n896 vcm.n895 0.00050467
R23349 vcm.n947 vcm.n946 0.00050467
R23350 vcm.n135 vcm.n134 0.00050467
R23351 vcm.n1018 vcm.n1017 0.00050467
R23352 vcm.n1092 vcm.n1091 0.00050467
R23353 vcm.n1086 vcm.n1085 0.00050467
R23354 vcm.n1100 vcm.n1099 0.00050467
R23355 vcm.n1166 vcm.n1165 0.00050467
R23356 vcm.n132 vcm.n131 0.00050467
R23357 vcm.n1180 vcm.n1179 0.00050467
R23358 vcm.n138 vcm.n137 0.00050467
R23359 vcm.n271 vcm.n270 0.00050467
R23360 vcm.n279 vcm.n278 0.00050467
R23361 vcm.n345 vcm.n344 0.00050467
R23362 vcm.n429 vcm.n428 0.00050467
R23363 vcm.n443 vcm.n442 0.00050467
R23364 vcm.n494 vcm.n493 0.00050467
R23365 vcm.n563 vcm.n562 0.00050467
R23366 vcm.n577 vcm.n576 0.00050467
R23367 vcm.n658 vcm.n657 0.00050467
R23368 vcm.n720 vcm.n719 0.00050467
R23369 vcm.n126 vcm.n125 0.00050467
R23370 vcm.n1185 vcm.n1184 0.00050467
R23371 vcm.n199 vcm.n198 0.000502311
R23372 vcm.n1186 vcm.n1185 0.000502311
R23373 vcm.n1179 vcm.n1178 0.000502311
R23374 vcm.n657 vcm.n656 0.000502311
R23375 vcm.n562 vcm.n561 0.000502311
R23376 vcm.n493 vcm.n492 0.000502311
R23377 vcm.n428 vcm.n427 0.000502311
R23378 vcm.n270 vcm.n269 0.000502311
R23379 vcm.n344 vcm.n343 0.000502311
R23380 vcm.n719 vcm.n718 0.000502311
R23381 vcm.n1085 vcm.n1084 0.000502311
R23382 vcm.n946 vcm.n945 0.000502311
R23383 vcm.n797 vcm.n796 0.000502311
R23384 vcm.n881 vcm.n880 0.000502311
R23385 vcm.n1017 vcm.n1016 0.000502311
R23386 vcm.n1165 vcm.n1164 0.000502311
R23387 vcm.n752 vcm.n751 0.000500172
R23388 vcm.n755 vcm.n754 0.000500095
R23389 vcm.n677 vcm.n676 0.000500095
C0 phi2_n mimtop2 0.0586f
C1 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 2.7e-20
C2 sky130_fd_sc_hd__buf_4_1/a_27_47# VDD 0.0671f
C3 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VDD 0.0203f
C4 mimtop1 phi2 0.0428f
C5 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# VDD 0.00178f
C6 mimtop1 sky130_fd_sc_hd__inv_1_3/Y 0.00363f
C7 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VDD 0.00498f
C8 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# vcm 0.037f
C9 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# VDD -2.7e-19
C10 VDD clk 0.172f
C11 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# VDD -0.00242f
C12 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# VDD 0.00475f
C13 mimbot1 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.028f
C14 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.00112f
C15 phi2 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.103f
C16 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.045f
C17 mimtop1 sky130_fd_sc_hd__inv_1_2/Y 0.00212f
C18 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.0578f
C19 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.0244f
C20 VDD vcm 46.2f
C21 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.0029f
C22 mimbot1 clk 0.00965f
C23 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.0067f
C24 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.0174f
C25 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__buf_4_3/a_27_47# 2.28e-19
C26 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 1.02e-19
C27 mimbot1 vcm 1.65f
C28 phi2_n sky130_fd_sc_hd__inv_1_1/A 6.18e-21
C29 phi2 sky130_fd_sc_hd__inv_1_3/A 0.00259f
C30 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.0584f
C31 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_3/Y 0.174f
C32 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.0137f
C33 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_1/A 0.0104f
C34 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_2/A 4.25e-19
C35 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 4.05e-19
C36 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 8.42e-20
C37 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 1.12e-19
C38 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 1.31e-20
C39 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_1/A 0.00778f
C40 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 2.97e-20
C41 phi1 sky130_fd_sc_hd__buf_4_1/a_27_47# 0.0991f
C42 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00335f
C43 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 1.32e-20
C44 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.0126f
C45 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.0126f
C46 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.0137f
C47 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 2.42e-19
C48 sky130_fd_sc_hd__nand2_1_1/a_113_47# vcm 2.3e-19
C49 sky130_fd_sc_hd__dlymetal6s6s_1_5/A sky130_fd_sc_hd__buf_4_0/a_27_47# 3.61e-19
C50 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 2.92e-21
C51 phi1_n sky130_fd_sc_hd__inv_1_4/Y 9.78e-20
C52 sky130_fd_sc_hd__nand2_1_0/Y phi1_n 0.00628f
C53 sky130_fd_sc_hd__nand2_1_1/Y VDD 0.106f
C54 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VDD 0.0184f
C55 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VDD 0.00342f
C56 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# vcm 0.0198f
C57 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# VDD -2.73e-19
C58 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# VDD 0.00766f
C59 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 4.65e-19
C60 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# VDD 0.00326f
C61 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/A 6.15e-19
C62 phi1 vcm 0.197f
C63 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 5.61e-19
C64 mimtop1 sky130_fd_sc_hd__buf_4_1/a_27_47# 1.48e-20
C65 mimbot1 sky130_fd_sc_hd__nand2_1_1/Y 9.9e-19
C66 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00195f
C67 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_4/A -7.45e-27
C68 VDD sky130_fd_sc_hd__buf_4_0/a_27_47# 0.0181f
C69 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.0122f
C70 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00152f
C71 mimtop1 clk 0.175f
C72 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.00204f
C73 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00101f
C74 phi1_n sky130_fd_sc_hd__inv_1_3/Y 0.0056f
C75 phi1_n sky130_fd_sc_hd__inv_1_2/A -4.02e-25
C76 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 1.86e-19
C77 mimbot1 sky130_fd_sc_hd__buf_4_0/a_27_47# 0.00827f
C78 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.0884f
C79 mimtop1 vcm 4.59f
C80 sky130_fd_sc_hd__inv_1_2/Y phi1_n 0.0108f
C81 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1_1/Y 4.69e-19
C82 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.0541f
C83 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.0012f
C84 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 2.17e-19
C85 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00223f
C86 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.0647f
C87 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 2.97e-20
C88 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 2.48e-19
C89 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# sky130_fd_sc_hd__inv_1_1/A 0.0211f
C90 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00883f
C91 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 3.29e-20
C92 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_3/A 7.55e-19
C93 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00232f
C94 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 3.52e-21
C95 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 4.65e-19
C96 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 4.65e-19
C97 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 6.18e-20
C98 phi2_n VDD 0.449f
C99 sky130_fd_sc_hd__inv_1_0/A VDD 0.256f
C100 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# VDD 0.00244f
C101 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# VDD 0.00764f
C102 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# mimtop2 0.00635f
C103 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# vcm 0.00609f
C104 phi1 sky130_fd_sc_hd__buf_4_0/a_27_47# 0.0148f
C105 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# VDD 0.00334f
C106 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 2.42e-19
C107 sky130_fd_sc_hd__buf_4_2/a_27_47# VDD 0.0172f
C108 mimbot1 phi2_n 0.152f
C109 mimtop1 sky130_fd_sc_hd__nand2_1_1/Y 0.0297f
C110 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00858f
C111 VDD mimtop2 1.66f
C112 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 3.99e-19
C113 sky130_fd_sc_hd__nand2_1_0/a_113_47# VDD -1.75e-19
C114 mimbot1 sky130_fd_sc_hd__buf_4_2/a_27_47# 7.45e-19
C115 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00736f
C116 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.0576f
C117 sky130_fd_sc_hd__buf_4_1/a_27_47# phi1_n 0.0184f
C118 mimbot1 mimtop2 1.54f
C119 mimbot1 sky130_fd_sc_hd__nand2_1_0/a_113_47# 4.99e-20
C120 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_4/A 3.28e-19
C121 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00211f
C122 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 7.06e-20
C123 phi1_n clk 0.00371f
C124 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 1.2e-19
C125 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.00629f
C126 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.00865f
C127 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 0.0467f
C128 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 3.81e-19
C129 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 8.17e-20
C130 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.0137f
C131 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 4.65e-19
C132 sky130_fd_sc_hd__dlymetal6s6s_1_2/A clk -6.85e-25
C133 phi1 sky130_fd_sc_hd__inv_1_0/A 0.00225f
C134 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 0.0111f
C135 phi1_n vcm 0.225f
C136 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 1.37e-19
C137 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.0126f
C138 phi1 sky130_fd_sc_hd__buf_4_2/a_27_47# 3.94e-20
C139 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# vcm 0.0611f
C140 sky130_fd_sc_hd__inv_1_1/A VDD 0.254f
C141 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# VDD 0.00492f
C142 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__buf_4_0/a_27_47# 3.37e-20
C143 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# VDD 0.00333f
C144 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# mimtop2 0.0175f
C145 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# vcm 5.29e-19
C146 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 2.37e-19
C147 phi1 mimtop2 0.0481f
C148 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# VDD 0.0493f
C149 mimtop1 phi2_n 0.0722f
C150 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00549f
C151 phi2_n sky130_fd_sc_hd__buf_4_3/a_27_47# 0.0174f
C152 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_4/Y 7.79e-19
C153 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# -1.06e-34
C154 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00449f
C155 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00768f
C156 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.0595f
C157 mimtop1 mimtop2 0.0211f
C158 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__buf_4_3/a_27_47# 6.05e-19
C159 sky130_fd_sc_hd__nand2_1_1/Y phi1_n 2.53e-19
C160 mimtop1 sky130_fd_sc_hd__nand2_1_0/a_113_47# 2.18e-19
C161 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00426f
C162 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00905f
C163 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.0654f
C164 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.0525f
C165 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 4.65e-19
C166 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.0171f
C167 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 2.56e-19
C168 sky130_fd_sc_hd__buf_4_3/a_27_47# mimtop2 4.27e-20
C169 phi2_n sky130_fd_sc_hd__inv_1_3/A 3.13e-25
C170 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.0126f
C171 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.0126f
C172 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_3/Y 0.234f
C173 phi1_n sky130_fd_sc_hd__buf_4_0/a_27_47# 8.88e-21
C174 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# 8.38e-19
C175 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.0204f
C176 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_4/Y 0.00111f
C177 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VDD 0.0184f
C178 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# vcm 0.0366f
C179 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__inv_1_2/Y 6.3e-20
C180 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# VDD 0.00717f
C181 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# mimtop2 0.0392f
C182 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 1.44e-19
C183 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VDD -0.00379f
C184 phi2 sky130_fd_sc_hd__inv_1_3/Y 0.248f
C185 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.00154f
C186 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00172f
C187 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 1.81e-19
C188 phi2 sky130_fd_sc_hd__inv_1_2/Y 2.22e-20
C189 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__inv_1_1/A 1.58e-20
C190 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_3/Y 0.279f
C191 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_2/A 0.172f
C192 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.00358f
C193 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.0141f
C194 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.0039f
C195 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.0536f
C196 phi2_n phi1_n 0.00349f
C197 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_2/A 0.00231f
C198 phi1_n sky130_fd_sc_hd__inv_1_0/A 1.03e-20
C199 mimbot1 VDD 1.69f
C200 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.00574f
C201 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_2/A 3.23e-19
C202 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.00736f
C203 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00146f
C204 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00151f
C205 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.0138f
C206 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 0.00445f
C207 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.0447f
C208 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 1.28e-19
C209 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 7.12e-19
C210 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_1/A 0.0512f
C211 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 2.14e-19
C212 phi1_n mimtop2 0.0612f
C213 sky130_fd_sc_hd__nand2_1_1/a_113_47# VDD -1.55e-19
C214 sky130_fd_sc_hd__dlymetal6s6s_1_2/A mimtop2 6.84e-19
C215 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# vcm 0.0173f
C216 sky130_fd_sc_hd__inv_1_4/Y clk 0.0432f
C217 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# mimtop2 0.0398f
C218 sky130_fd_sc_hd__nand2_1_0/Y clk 0.0401f
C219 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 1.52e-19
C220 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# VDD -0.00169f
C221 phi1 VDD 0.198f
C222 mimbot1 sky130_fd_sc_hd__nand2_1_1/a_113_47# 4.07e-20
C223 vcm sky130_fd_sc_hd__inv_1_4/Y 0.00464f
C224 sky130_fd_sc_hd__nand2_1_0/Y vcm 0.179f
C225 phi2 sky130_fd_sc_hd__buf_4_1/a_27_47# 3.43e-21
C226 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 6.64e-20
C227 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00381f
C228 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 6.37e-19
C229 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/A 4.55e-19
C230 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_2/A 7.06e-21
C231 mimbot1 phi1 0.0816f
C232 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 1.22e-19
C233 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00188f
C234 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.00384f
C235 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.00678f
C236 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00255f
C237 sky130_fd_sc_hd__inv_1_3/Y clk 8.23e-19
C238 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.0607f
C239 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__inv_1_2/A 2.42e-19
C240 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__inv_1_2/A 0.0111f
C241 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__buf_4_1/a_27_47# 0.0372f
C242 mimtop1 VDD 1.51f
C243 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 7.18e-20
C244 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 0.00468f
C245 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.0667f
C246 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.00449f
C247 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.0631f
C248 phi2 vcm 0.0265f
C249 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 3.08e-19
C250 sky130_fd_sc_hd__inv_1_2/Y clk 2.81e-19
C251 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.105f
C252 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# 0.00169f
C253 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# sky130_fd_sc_hd__inv_1_0/A 6.92e-21
C254 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.0267f
C255 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00117f
C256 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.00446f
C257 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.0533f
C258 sky130_fd_sc_hd__inv_1_3/Y vcm 0.21f
C259 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00865f
C260 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.0137f
C261 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 0.0137f
C262 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 7.12e-19
C263 sky130_fd_sc_hd__buf_4_3/a_27_47# VDD 0.0648f
C264 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 0.0126f
C265 mimbot1 mimtop1 1.31f
C266 sky130_fd_sc_hd__inv_1_2/Y vcm 0.216f
C267 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__buf_4_0/a_27_47# 0.00416f
C268 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_4/Y 0.0222f
C269 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# mimtop2 0.00804f
C270 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# vcm 0.00547f
C271 mimbot1 sky130_fd_sc_hd__buf_4_3/a_27_47# 0.00895f
C272 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_1/Y 0.0147f
C273 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 7.34e-20
C274 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# VDD -0.0021f
C275 sky130_fd_sc_hd__inv_1_3/A VDD 0.169f
C276 mimtop1 sky130_fd_sc_hd__nand2_1_1/a_113_47# 2.3e-19
C277 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.002f
C278 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.0012f
C279 mimbot1 sky130_fd_sc_hd__inv_1_3/A 2.31e-19
C280 mimtop1 phi1 0.074f
C281 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_3/Y 7.86e-19
C282 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.0176f
C283 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.00644f
C284 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 0.00493f
C285 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 0.00181f
C286 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.063f
C287 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_2/A 3.52e-21
C288 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__inv_1_2/A 8.38e-19
C289 phi1 sky130_fd_sc_hd__buf_4_3/a_27_47# 1.79e-21
C290 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__nand2_1_1/Y 0.259f
C291 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00594f
C292 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00283f
C293 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# 0.00358f
C294 phi2 sky130_fd_sc_hd__buf_4_0/a_27_47# 4.02e-20
C295 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 0.0474f
C296 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 0.105f
C297 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 4.65e-19
C298 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 3.38e-19
C299 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__inv_1_0/A 0.00215f
C300 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# 6.66e-19
C301 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__inv_1_0/A 1.91e-20
C302 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# 0.0222f
C303 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00117f
C304 sky130_fd_sc_hd__dlymetal6s6s_1_4/A clk -3.91e-26
C305 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.005f
C306 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.0171f
C307 sky130_fd_sc_hd__buf_4_0/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.0201f
C308 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 4.65e-19
C309 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 4.65e-19
C310 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 4.65e-19
C311 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 4.65e-19
C312 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 1.92e-19
C313 sky130_fd_sc_hd__buf_4_1/a_27_47# vcm 0.00117f
C314 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__buf_4_0/a_27_47# 0.171f
C315 sky130_fd_sc_hd__dlymetal6s6s_1_4/A vcm -4.89e-24
C316 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__buf_4_0/a_27_47# 1.92e-19
C317 sky130_fd_sc_hd__nand2_1_0/Y phi2_n 2.59e-20
C318 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__buf_4_0/a_27_47# 7.18e-20
C319 phi1_n VDD 0.532f
C320 vcm clk 0.00409f
C321 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# mimtop2 0.0188f
C322 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# vcm 3.01e-20
C323 mimtop1 sky130_fd_sc_hd__buf_4_3/a_27_47# 2.61e-19
C324 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# VDD 0.0529f
C325 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VDD 0.00998f
C326 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# VDD -0.00122f
C327 mimbot1 phi1_n 0.14f
C328 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# -5.66e-37
C329 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.0575f
C330 sky130_fd_sc_hd__nand2_1_0/Y mimtop2 6.91e-19
C331 phi2 phi2_n 0.647f
C332 phi2_n sky130_fd_sc_hd__inv_1_3/Y 0.00875f
C333 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1_0/Y 5.19e-19
C334 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 5.19e-19
C335 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.0178f
C336 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_0/A 0.0075f
C337 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 4.88e-20
C338 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_2/A 0.04f
C339 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.00861f
C340 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# 0.00309f
C341 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 0.00134f
C342 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# sky130_fd_sc_hd__inv_1_2/A 1.37e-19
C343 phi2 sky130_fd_sc_hd__buf_4_2/a_27_47# 0.0172f
C344 sky130_fd_sc_hd__inv_1_2/Y phi2_n 1.74e-19
C345 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__inv_1_2/A 1.97e-19
C346 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.174f
C347 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 1.21e-19
C348 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_0/A 0.0271f
C349 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__inv_1_2/A 3.37e-20
C350 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/A 6.68e-19
C351 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00678f
C352 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 1.85e-19
C353 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.0548f
C354 phi2 mimtop2 0.0606f
C355 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# 1.31e-19
C356 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# sky130_fd_sc_hd__inv_1_0/A 0.00325f
C357 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# 7.49e-19
C358 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__inv_1_0/A 1.31e-20
C359 sky130_fd_sc_hd__nand2_1_1/Y clk 0.00909f
C360 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.00865f
C361 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 4.28e-19
C362 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00322f
C363 sky130_fd_sc_hd__inv_1_3/Y mimtop2 0.0818f
C364 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.0126f
C365 phi1 phi1_n 0.785f
C366 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# 0.0126f
C367 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__buf_4_0/a_27_47# 6.05e-19
C368 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# 0.00416f
C369 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 0.0137f
C370 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/A 2e-20
C371 sky130_fd_sc_hd__inv_1_2/Y mimtop2 0.08f
C372 sky130_fd_sc_hd__nand2_1_1/Y vcm 0.171f
C373 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# mimtop2 0.0419f
C374 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# VDD -0.0028f
C375 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VDD 0.0039f
C376 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.0386f
C377 mimtop1 phi1_n 0.0579f
C378 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.0295f
C379 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 2.14e-21
C380 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 8.06e-19
C381 phi1_n sky130_fd_sc_hd__buf_4_3/a_27_47# 1.3e-20
C382 phi2 sky130_fd_sc_hd__inv_1_1/A 0.00236f
C383 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 5.6e-19
C384 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_1/A 0.0364f
C385 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 4.84e-21
C386 sky130_fd_sc_hd__buf_4_1/a_27_47# phi2_n 1.3e-20
C387 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.021f
C388 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 0.00242f
C389 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 0.0542f
C390 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__inv_1_0/A 1.89e-19
C391 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_4/A 0.00187f
C392 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 5.64e-19
C393 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 1.02e-19
C394 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_1/A 8.25e-20
C395 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# 0.00393f
C396 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 4.65e-19
C397 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__inv_1_1/A 0.00215f
C398 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 2.65e-19
C399 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.0413f
C400 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 1.72e-19
C401 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# sky130_fd_sc_hd__inv_1_0/A 0.00429f
C402 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__inv_1_0/A 1.2e-19
C403 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/A 0.0171f
C404 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# 0.00489f
C405 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 7.12e-19
C406 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 3.29e-20
C407 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# 7.18e-20
C408 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 4.65e-19
C409 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 4.65e-19
C410 phi2_n vcm 0.031f
C411 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00865f
C412 sky130_fd_sc_hd__buf_4_1/a_27_47# mimtop2 4.98e-20
C413 phi1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 5.55e-20
C414 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__buf_4_0/a_27_47# 0.00883f
C415 sky130_fd_sc_hd__dlymetal6s6s_1_4/A mimtop2 4.9e-19
C416 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# mimtop2 0.0383f
C417 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# VDD 0.00405f
C418 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VDD -0.00386f
C419 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# VDD 0.00288f
C420 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.00493f
C421 vcm mimtop2 3.21f
C422 sky130_fd_sc_hd__nand2_1_0/a_113_47# vcm 2.27e-19
C423 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# 0.00163f
C424 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 0.0137f
C425 mimtop1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 3.04e-20
C426 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.00194f
C427 VDD sky130_fd_sc_hd__inv_1_4/Y 0.0709f
C428 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_5/A 7.55e-19
C429 sky130_fd_sc_hd__nand2_1_0/Y VDD 0.0452f
C430 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.0282f
C431 phi2 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 6.99e-20
C432 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.0273f
C433 sky130_fd_sc_hd__nand2_1_1/Y phi2_n 0.00587f
C434 mimbot1 sky130_fd_sc_hd__inv_1_4/Y 0.00182f
C435 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 0.0599f
C436 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 4.05e-19
C437 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.003f
C438 mimbot1 sky130_fd_sc_hd__nand2_1_0/Y 0.0025f
C439 sky130_fd_sc_hd__buf_4_1/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 1.86e-19
C440 sky130_fd_sc_hd__dlymetal6s6s_1_3/A sky130_fd_sc_hd__inv_1_0/A 0.00211f
C441 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# 1.73e-19
C442 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.00235f
C443 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/A 0.105f
C444 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# 6.92e-21
C445 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# sky130_fd_sc_hd__inv_1_1/A 0.00325f
C446 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 1.19e-19
C447 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 0.0264f
C448 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__inv_1_0/A 0.00778f
C449 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__inv_1_0/A 4.96e-19
C450 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# 0.00604f
C451 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# 1.32e-20
C452 phi2 VDD 0.262f
C453 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 0.0137f
C454 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# 0.0137f
C455 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_3/A 3.61e-19
C456 sky130_fd_sc_hd__inv_1_3/Y VDD 0.62f
C457 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 7.12e-19
C458 VDD sky130_fd_sc_hd__inv_1_2/A 0.134f
C459 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# 0.0126f
C460 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/A 0.0171f
C461 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__buf_4_0/a_27_47# 0.00343f
C462 sky130_fd_sc_hd__nand2_1_1/Y mimtop2 5.76e-19
C463 sky130_fd_sc_hd__inv_1_2/Y VDD 0.366f
C464 mimbot1 phi2 0.118f
C465 mimbot1 sky130_fd_sc_hd__inv_1_3/Y 0.134f
C466 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# VDD 0.00405f
C467 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# vcm 0.0628f
C468 sky130_fd_sc_hd__buf_4_2/a_27_47# sky130_fd_sc_hd__buf_4_0/a_27_47# 0.00102f
C469 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VDD 0.005f
C470 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# VDD -0.0022f
C471 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# VDD 0.00408f
C472 mimbot1 sky130_fd_sc_hd__inv_1_2/A 0.00628f
C473 sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.00169f
C474 mimbot1 sky130_fd_sc_hd__inv_1_2/Y 0.165f
C475 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# 0.00226f
C476 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# 0.0119f
C477 mimbot1 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# 0.00109f
C478 sky130_fd_sc_hd__buf_4_3/a_27_47# sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# 1.21e-19
C479 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_2/Y 1.16e-19
C480 phi2 phi1 1e-23
C481 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 0.0535f
C482 mimtop1 sky130_fd_sc_hd__inv_1_4/Y 0.0294f
C483 phi1 sky130_fd_sc_hd__inv_1_3/Y 1.81e-19
C484 phi2_n sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# 0.0012f
C485 sky130_fd_sc_hd__dlymetal6s6s_1_4/A sky130_fd_sc_hd__dlymetal6s6s_1_5/A 1.91e-24
C486 mimtop1 sky130_fd_sc_hd__nand2_1_0/Y 0.0311f
C487 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 6.38e-19
C488 phi1_n sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# 2.36e-19
C489 phi1 sky130_fd_sc_hd__inv_1_2/A 0.00226f
C490 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# 1.91e-20
C491 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# sky130_fd_sc_hd__inv_1_1/A 0.00429f
C492 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 1.74e-19
C493 phi2_n sky130_fd_sc_hd__buf_4_2/a_27_47# 8.34e-21
C494 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__inv_1_0/A 0.0211f
C495 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# 3.29e-20
C496 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# 4.65e-19
C497 sky130_fd_sc_hd__dlymetal6s6s_1_2/A sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# 0.105f
C498 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# 4.65e-19
C499 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# 4.65e-19
C500 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# 4.65e-19
C501 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# 4.65e-19
C502 sky130_fd_sc_hd__inv_1_2/Y phi1 0.252f
C503 vcm.n0 VSS 2.37f
C504 vcm.n1 VSS 0.242f
C505 vcm.n2 VSS 2.37f
C506 vcm.n3 VSS 0.242f
C507 vcm.n4 VSS 2.37f
C508 vcm.n5 VSS 0.242f
C509 vcm.n6 VSS 2.37f
C510 vcm.n7 VSS 0.242f
C511 vcm.t47 VSS 7.36f
C512 vcm.n8 VSS 0.502f
C513 vcm.n9 VSS 2.37f
C514 vcm.n10 VSS 0.251f
C515 vcm.n11 VSS 0.0569f
C516 vcm.n12 VSS -0.398f
C517 vcm.n13 VSS 0.0142f
C518 vcm.n14 VSS 0.502f
C519 vcm.n15 VSS 2.37f
C520 vcm.n16 VSS 0.251f
C521 vcm.n17 VSS 0.0569f
C522 vcm.n18 VSS -0.398f
C523 vcm.n19 VSS 0.404f
C524 vcm.n20 VSS -0.0314f
C525 vcm.n21 VSS -0.341f
C526 vcm.n22 VSS -0.287f
C527 vcm.n23 VSS 0.427f
C528 vcm.n24 VSS -0.0315f
C529 vcm.n25 VSS -0.364f
C530 vcm.n26 VSS -0.287f
C531 vcm.n27 VSS -0.356f
C532 vcm.n28 VSS 2.37f
C533 vcm.n29 VSS 1f
C534 vcm.n30 VSS 0.242f
C535 vcm.n31 VSS 0.157f
C536 vcm.n32 VSS -0.356f
C537 vcm.n33 VSS 0.0139f
C538 vcm.n34 VSS 0.404f
C539 vcm.n35 VSS -0.0312f
C540 vcm.n36 VSS 2.37f
C541 vcm.n37 VSS 0.242f
C542 vcm.n38 VSS -0.356f
C543 vcm.t46 VSS 7.36f
C544 vcm.n39 VSS 2.37f
C545 vcm.n40 VSS 1f
C546 vcm.n41 VSS 0.242f
C547 vcm.n42 VSS 0.157f
C548 vcm.n43 VSS -0.356f
C549 vcm.n44 VSS 0.426f
C550 vcm.n45 VSS -0.0315f
C551 vcm.n46 VSS -0.364f
C552 vcm.n47 VSS -0.287f
C553 vcm.n48 VSS -0.341f
C554 vcm.n49 VSS -0.287f
C555 vcm.n50 VSS -0.356f
C556 vcm.t55 VSS 7.36f
C557 vcm.n51 VSS 2.37f
C558 vcm.n52 VSS 1f
C559 vcm.n53 VSS 0.242f
C560 vcm.n54 VSS 0.157f
C561 vcm.n55 VSS -0.356f
C562 vcm.n56 VSS 0.0142f
C563 vcm.n57 VSS 0.427f
C564 vcm.n58 VSS -0.0315f
C565 vcm.n59 VSS -0.364f
C566 vcm.n60 VSS -0.287f
C567 vcm.n61 VSS -0.356f
C568 vcm.t63 VSS 7.36f
C569 vcm.n62 VSS 2.37f
C570 vcm.n63 VSS 1f
C571 vcm.n64 VSS 0.242f
C572 vcm.n65 VSS 0.157f
C573 vcm.n66 VSS -0.356f
C574 vcm.n67 VSS 0.0139f
C575 vcm.n68 VSS 0.404f
C576 vcm.n69 VSS -0.0312f
C577 vcm.n70 VSS 2.37f
C578 vcm.n71 VSS 0.242f
C579 vcm.n72 VSS 2.37f
C580 vcm.n73 VSS 0.242f
C581 vcm.n74 VSS -0.356f
C582 vcm.t54 VSS 7.36f
C583 vcm.n75 VSS 2.37f
C584 vcm.n76 VSS 1f
C585 vcm.n77 VSS 0.242f
C586 vcm.n78 VSS 0.157f
C587 vcm.n79 VSS -0.356f
C588 vcm.n80 VSS 0.404f
C589 vcm.n81 VSS -0.0314f
C590 vcm.n82 VSS -0.341f
C591 vcm.n83 VSS -0.287f
C592 vcm.n84 VSS -0.356f
C593 vcm.t62 VSS 7.36f
C594 vcm.n85 VSS 2.37f
C595 vcm.n86 VSS 1f
C596 vcm.n87 VSS 0.242f
C597 vcm.n88 VSS 0.157f
C598 vcm.n89 VSS -0.356f
C599 vcm.n90 VSS 0.426f
C600 vcm.n91 VSS -0.0315f
C601 vcm.n92 VSS -0.364f
C602 vcm.n93 VSS -0.287f
C603 vcm.n94 VSS -0.341f
C604 vcm.n95 VSS -0.287f
C605 vcm.n96 VSS -0.356f
C606 vcm.t71 VSS 7.36f
C607 vcm.n97 VSS 2.37f
C608 vcm.n98 VSS 1f
C609 vcm.n99 VSS 0.242f
C610 vcm.n100 VSS 0.157f
C611 vcm.n101 VSS -0.356f
C612 vcm.n102 VSS 0.0142f
C613 vcm.n103 VSS 2.37f
C614 vcm.n104 VSS 0.242f
C615 vcm.n105 VSS -0.356f
C616 vcm.t70 VSS 7.36f
C617 vcm.n106 VSS 2.37f
C618 vcm.n107 VSS 1f
C619 vcm.n108 VSS 0.242f
C620 vcm.n109 VSS 0.157f
C621 vcm.n110 VSS -0.356f
C622 vcm.n111 VSS 0.404f
C623 vcm.n112 VSS -0.0314f
C624 vcm.n113 VSS -0.341f
C625 vcm.n114 VSS -0.287f
C626 vcm.n115 VSS 0.427f
C627 vcm.n116 VSS -0.0315f
C628 vcm.n117 VSS -0.364f
C629 vcm.n118 VSS -0.287f
C630 vcm.n119 VSS 0.331f
C631 vcm.t79 VSS 7.36f
C632 vcm.n120 VSS 2.39f
C633 vcm.n121 VSS -0.379f
C634 vcm.n122 VSS 0.156f
C635 vcm.n123 VSS 0.146f
C636 vcm.n124 VSS 0.0526f
C637 vcm.n125 VSS 0.0393f
C638 vcm.n126 VSS 0.0393f
C639 vcm.n128 VSS 1.01f
C640 vcm.n130 VSS 0.0526f
C641 vcm.n131 VSS 0.0393f
C642 vcm.n132 VSS 0.0393f
C643 vcm.n133 VSS 0.0526f
C644 vcm.n134 VSS 0.0393f
C645 vcm.n135 VSS 0.0393f
C646 vcm.n136 VSS 0.0526f
C647 vcm.n137 VSS 0.0393f
C648 vcm.n138 VSS 0.0393f
C649 vcm.n139 VSS 0.0526f
C650 vcm.n140 VSS 0.0393f
C651 vcm.n141 VSS 0.0393f
C652 vcm.n143 VSS 1.09f
C653 vcm.n144 VSS 0.146f
C654 vcm.n146 VSS 0.242f
C655 vcm.n147 VSS 0.0585f
C656 vcm.n148 VSS 2.37f
C657 vcm.t24 VSS 7.36f
C658 vcm.n149 VSS 2.37f
C659 vcm.n150 VSS 2.37f
C660 vcm.t8 VSS 7.36f
C661 vcm.n151 VSS 2.37f
C662 vcm.t0 VSS 16.7f
C663 vcm.n152 VSS 0.446f
C664 vcm.n153 VSS 0.251f
C665 vcm.n154 VSS 0.0569f
C666 vcm.n155 VSS -1.34f
C667 vcm.n156 VSS 0.0144f
C668 vcm.n157 VSS -0.288f
C669 vcm.n158 VSS -0.356f
C670 vcm.n159 VSS -0.332f
C671 vcm.n160 VSS 1f
C672 vcm.n161 VSS 0.158f
C673 vcm.n162 VSS 0.241f
C674 vcm.n163 VSS 0.241f
C675 vcm.n164 VSS -0.356f
C676 vcm.n165 VSS 0.0144f
C677 vcm.n166 VSS -0.288f
C678 vcm.n167 VSS -0.356f
C679 vcm.n168 VSS 2.37f
C680 vcm.n169 VSS 1f
C681 vcm.n170 VSS 0.158f
C682 vcm.n171 VSS 0.241f
C683 vcm.n172 VSS 0.241f
C684 vcm.n173 VSS -0.356f
C685 vcm.n174 VSS 0.0144f
C686 vcm.n175 VSS -0.288f
C687 vcm.n176 VSS -0.356f
C688 vcm.t16 VSS 7.36f
C689 vcm.n177 VSS 2.37f
C690 vcm.n178 VSS 1f
C691 vcm.n179 VSS 0.158f
C692 vcm.n180 VSS 0.241f
C693 vcm.n181 VSS 0.241f
C694 vcm.n182 VSS -0.356f
C695 vcm.n183 VSS 0.0144f
C696 vcm.n184 VSS -0.288f
C697 vcm.n185 VSS -0.356f
C698 vcm.n186 VSS 2.37f
C699 vcm.n187 VSS 1f
C700 vcm.n188 VSS 0.158f
C701 vcm.n189 VSS 0.241f
C702 vcm.n190 VSS 0.241f
C703 vcm.n191 VSS -0.356f
C704 vcm.n192 VSS 0.0144f
C705 vcm.n193 VSS -0.288f
C706 vcm.n194 VSS -0.398f
C707 vcm.t32 VSS 7.36f
C708 vcm.n195 VSS 2.39f
C709 vcm.n196 VSS 0.323f
C710 vcm.n197 VSS 0.193f
C711 vcm.n198 VSS 0.21f
C712 vcm.n199 VSS 0.0444f
C713 vcm.n200 VSS 0.0444f
C714 vcm.n202 VSS 1f
C715 vcm.n203 VSS 1f
C716 vcm.n204 VSS 0.146f
C717 vcm.n206 VSS 2.37f
C718 vcm.n207 VSS 2.37f
C719 vcm.t17 VSS 7.36f
C720 vcm.n208 VSS 2.37f
C721 vcm.n209 VSS 2.37f
C722 vcm.n210 VSS 0.502f
C723 vcm.n211 VSS 2.37f
C724 vcm.n212 VSS 0.251f
C725 vcm.n213 VSS 0.0569f
C726 vcm.n214 VSS -0.398f
C727 vcm.n215 VSS 0.404f
C728 vcm.n216 VSS -0.0314f
C729 vcm.n217 VSS -0.341f
C730 vcm.n218 VSS -0.287f
C731 vcm.n219 VSS -0.356f
C732 vcm.t1 VSS 7.36f
C733 vcm.n220 VSS 2.37f
C734 vcm.n221 VSS 1f
C735 vcm.n222 VSS 0.158f
C736 vcm.n223 VSS 0.241f
C737 vcm.n224 VSS 0.241f
C738 vcm.n225 VSS -0.356f
C739 vcm.n226 VSS 0.404f
C740 vcm.n227 VSS -0.0314f
C741 vcm.n228 VSS -0.341f
C742 vcm.n229 VSS -0.287f
C743 vcm.n230 VSS -0.356f
C744 vcm.t9 VSS 7.36f
C745 vcm.n231 VSS 2.37f
C746 vcm.n232 VSS 1f
C747 vcm.n233 VSS 0.158f
C748 vcm.n234 VSS 0.241f
C749 vcm.n235 VSS 0.241f
C750 vcm.n236 VSS -0.356f
C751 vcm.n237 VSS 0.427f
C752 vcm.n238 VSS -0.0315f
C753 vcm.n239 VSS -0.364f
C754 vcm.n240 VSS -0.287f
C755 vcm.n241 VSS -0.356f
C756 vcm.n242 VSS 2.37f
C757 vcm.n243 VSS 1f
C758 vcm.n244 VSS 0.158f
C759 vcm.n245 VSS 0.241f
C760 vcm.n246 VSS 0.241f
C761 vcm.n247 VSS -0.356f
C762 vcm.n248 VSS 0.404f
C763 vcm.n249 VSS -0.0314f
C764 vcm.n250 VSS -0.341f
C765 vcm.n251 VSS -0.287f
C766 vcm.n252 VSS -0.356f
C767 vcm.t25 VSS 7.36f
C768 vcm.n253 VSS 2.37f
C769 vcm.n254 VSS 1f
C770 vcm.n255 VSS 0.149f
C771 vcm.n256 VSS 0.243f
C772 vcm.n257 VSS 0.248f
C773 vcm.n258 VSS -0.356f
C774 vcm.n259 VSS 0.403f
C775 vcm.n260 VSS -0.0296f
C776 vcm.n261 VSS -0.34f
C777 vcm.n262 VSS -0.287f
C778 vcm.n263 VSS 0.242f
C779 vcm.n264 VSS 0.0585f
C780 vcm.n265 VSS -0.398f
C781 vcm.t33 VSS 7.36f
C782 vcm.n266 VSS 2.39f
C783 vcm.n267 VSS 0.323f
C784 vcm.n268 VSS 0.192f
C785 vcm.n269 VSS 0.21f
C786 vcm.n270 VSS 0.0444f
C787 vcm.n271 VSS 0.0444f
C788 vcm.n273 VSS 1f
C789 vcm.n274 VSS 1f
C790 vcm.n275 VSS 0.146f
C791 vcm.n277 VSS 0.0526f
C792 vcm.n278 VSS 0.0393f
C793 vcm.n279 VSS 0.0393f
C794 vcm.n280 VSS 0.242f
C795 vcm.n281 VSS 0.0587f
C796 vcm.n282 VSS 2.37f
C797 vcm.t26 VSS 7.36f
C798 vcm.n283 VSS 2.37f
C799 vcm.t18 VSS 7.36f
C800 vcm.n284 VSS 2.37f
C801 vcm.t10 VSS 7.36f
C802 vcm.n285 VSS 2.37f
C803 vcm.t2 VSS 7.36f
C804 vcm.n286 VSS 0.502f
C805 vcm.n287 VSS 2.37f
C806 vcm.n288 VSS 0.251f
C807 vcm.n289 VSS 0.0569f
C808 vcm.n290 VSS -0.398f
C809 vcm.n291 VSS 0.426f
C810 vcm.n292 VSS -0.0315f
C811 vcm.n293 VSS -0.364f
C812 vcm.n294 VSS -0.287f
C813 vcm.n295 VSS -0.356f
C814 vcm.n296 VSS 2.37f
C815 vcm.n297 VSS 1f
C816 vcm.n298 VSS 0.158f
C817 vcm.n299 VSS 0.241f
C818 vcm.n300 VSS 0.241f
C819 vcm.n301 VSS -0.356f
C820 vcm.n302 VSS 0.404f
C821 vcm.n303 VSS -0.0314f
C822 vcm.n304 VSS -0.341f
C823 vcm.n305 VSS -0.287f
C824 vcm.n306 VSS -0.356f
C825 vcm.n307 VSS 2.37f
C826 vcm.n308 VSS 1f
C827 vcm.n309 VSS 0.158f
C828 vcm.n310 VSS 0.241f
C829 vcm.n311 VSS 0.241f
C830 vcm.n312 VSS -0.356f
C831 vcm.n313 VSS 0.404f
C832 vcm.n314 VSS -0.0314f
C833 vcm.n315 VSS -0.341f
C834 vcm.n316 VSS -0.287f
C835 vcm.n317 VSS -0.356f
C836 vcm.n318 VSS 2.37f
C837 vcm.n319 VSS 1f
C838 vcm.n320 VSS 0.149f
C839 vcm.n321 VSS 0.243f
C840 vcm.n322 VSS 0.248f
C841 vcm.n323 VSS -0.356f
C842 vcm.n324 VSS 0.403f
C843 vcm.n325 VSS -0.0297f
C844 vcm.n326 VSS -0.34f
C845 vcm.n327 VSS -0.287f
C846 vcm.n328 VSS -0.356f
C847 vcm.n329 VSS 2.37f
C848 vcm.n330 VSS 1f
C849 vcm.n331 VSS 0.158f
C850 vcm.n332 VSS 0.241f
C851 vcm.n333 VSS 0.241f
C852 vcm.n334 VSS -0.356f
C853 vcm.n335 VSS 0.403f
C854 vcm.n336 VSS -0.0296f
C855 vcm.n337 VSS -0.34f
C856 vcm.n338 VSS -0.287f
C857 vcm.n339 VSS -0.398f
C858 vcm.t34 VSS 7.36f
C859 vcm.n340 VSS 2.39f
C860 vcm.n341 VSS 0.323f
C861 vcm.n342 VSS 0.193f
C862 vcm.n343 VSS 0.21f
C863 vcm.n344 VSS 0.0444f
C864 vcm.n345 VSS 0.0444f
C865 vcm.n347 VSS 0.993f
C866 vcm.n348 VSS 0.993f
C867 vcm.t35 VSS 7.36f
C868 vcm.n349 VSS 0.403f
C869 vcm.n350 VSS -0.0297f
C870 vcm.n351 VSS -0.34f
C871 vcm.n352 VSS 0.403f
C872 vcm.n353 VSS -0.0296f
C873 vcm.n354 VSS -0.34f
C874 vcm.n355 VSS 2.37f
C875 vcm.n356 VSS 2.37f
C876 vcm.t19 VSS 7.36f
C877 vcm.n357 VSS 2.37f
C878 vcm.n358 VSS 2.37f
C879 vcm.n359 VSS 0.502f
C880 vcm.n360 VSS 2.37f
C881 vcm.n361 VSS 0.251f
C882 vcm.n362 VSS 0.0569f
C883 vcm.n363 VSS -0.398f
C884 vcm.n364 VSS 0.404f
C885 vcm.n365 VSS -0.0314f
C886 vcm.n366 VSS -0.341f
C887 vcm.n367 VSS 0.404f
C888 vcm.n368 VSS -0.0314f
C889 vcm.n369 VSS -0.341f
C890 vcm.n370 VSS -0.287f
C891 vcm.n371 VSS -0.356f
C892 vcm.t3 VSS 7.36f
C893 vcm.n372 VSS 2.37f
C894 vcm.n373 VSS 1f
C895 vcm.n374 VSS 0.158f
C896 vcm.n375 VSS 0.241f
C897 vcm.n376 VSS 0.241f
C898 vcm.n377 VSS -0.356f
C899 vcm.n378 VSS 0.403f
C900 vcm.n379 VSS -0.0297f
C901 vcm.n380 VSS -0.34f
C902 vcm.n381 VSS 0.426f
C903 vcm.n382 VSS -0.0315f
C904 vcm.n383 VSS -0.364f
C905 vcm.n384 VSS -0.287f
C906 vcm.n385 VSS -0.356f
C907 vcm.t11 VSS 7.36f
C908 vcm.n386 VSS 2.37f
C909 vcm.n387 VSS 1f
C910 vcm.n388 VSS 0.149f
C911 vcm.n389 VSS 0.243f
C912 vcm.n390 VSS 0.248f
C913 vcm.n391 VSS -0.356f
C914 vcm.n392 VSS 0.403f
C915 vcm.n393 VSS -0.0296f
C916 vcm.n394 VSS -0.34f
C917 vcm.n395 VSS 0.403f
C918 vcm.n396 VSS -0.0296f
C919 vcm.n397 VSS -0.34f
C920 vcm.n398 VSS -0.287f
C921 vcm.n399 VSS -0.356f
C922 vcm.n400 VSS 2.37f
C923 vcm.n401 VSS 1f
C924 vcm.n402 VSS 0.158f
C925 vcm.n403 VSS 0.241f
C926 vcm.n404 VSS 0.241f
C927 vcm.n405 VSS -0.356f
C928 vcm.n406 VSS 0.403f
C929 vcm.n407 VSS -0.0296f
C930 vcm.n408 VSS -0.34f
C931 vcm.n409 VSS 0.403f
C932 vcm.n410 VSS -0.0296f
C933 vcm.n411 VSS -0.34f
C934 vcm.n412 VSS -0.287f
C935 vcm.n413 VSS -0.356f
C936 vcm.t27 VSS 7.36f
C937 vcm.n414 VSS 2.37f
C938 vcm.n415 VSS 1f
C939 vcm.n416 VSS 0.158f
C940 vcm.n417 VSS 0.241f
C941 vcm.n418 VSS 0.241f
C942 vcm.n419 VSS -0.356f
C943 vcm.n420 VSS -0.287f
C944 vcm.n421 VSS -0.398f
C945 vcm.n422 VSS 2.39f
C946 vcm.n423 VSS 0.325f
C947 vcm.n424 VSS 0.242f
C948 vcm.n425 VSS 0.0581f
C949 vcm.n426 VSS 0.191f
C950 vcm.n427 VSS 0.21f
C951 vcm.n428 VSS 0.0444f
C952 vcm.n429 VSS 0.0444f
C953 vcm.n431 VSS 0.0526f
C954 vcm.n432 VSS 0.0393f
C955 vcm.n433 VSS 0.0393f
C956 vcm.n435 VSS 0.146f
C957 vcm.n437 VSS 0.956f
C958 vcm.n438 VSS 0.956f
C959 vcm.n439 VSS 0.146f
C960 vcm.n441 VSS 0.0526f
C961 vcm.n442 VSS 0.0393f
C962 vcm.n443 VSS 0.0393f
C963 vcm.n444 VSS 2.37f
C964 vcm.t28 VSS 7.36f
C965 vcm.n445 VSS 2.37f
C966 vcm.n446 VSS 2.37f
C967 vcm.t12 VSS 7.36f
C968 vcm.n447 VSS 2.37f
C969 vcm.n448 VSS 0.502f
C970 vcm.n449 VSS 2.37f
C971 vcm.n450 VSS 0.251f
C972 vcm.n451 VSS 0.0569f
C973 vcm.n452 VSS -0.398f
C974 vcm.n453 VSS -0.287f
C975 vcm.n454 VSS -0.356f
C976 vcm.t4 VSS 7.36f
C977 vcm.n455 VSS 2.37f
C978 vcm.n456 VSS 1f
C979 vcm.n457 VSS 0.149f
C980 vcm.n458 VSS 0.243f
C981 vcm.n459 VSS 0.248f
C982 vcm.n460 VSS -0.356f
C983 vcm.n461 VSS -0.287f
C984 vcm.n462 VSS -0.356f
C985 vcm.n463 VSS 2.37f
C986 vcm.n464 VSS 1f
C987 vcm.n465 VSS 0.158f
C988 vcm.n466 VSS 0.241f
C989 vcm.n467 VSS 0.241f
C990 vcm.n468 VSS -0.356f
C991 vcm.n469 VSS -0.287f
C992 vcm.n470 VSS -0.356f
C993 vcm.t20 VSS 7.36f
C994 vcm.n471 VSS 2.37f
C995 vcm.n472 VSS 1f
C996 vcm.n473 VSS 0.158f
C997 vcm.n474 VSS 0.241f
C998 vcm.n475 VSS 0.241f
C999 vcm.n476 VSS -0.356f
C1000 vcm.n477 VSS -0.287f
C1001 vcm.n478 VSS -0.356f
C1002 vcm.n479 VSS 2.37f
C1003 vcm.n480 VSS 1f
C1004 vcm.n481 VSS 0.158f
C1005 vcm.n482 VSS 0.241f
C1006 vcm.n483 VSS 0.241f
C1007 vcm.n484 VSS -0.356f
C1008 vcm.n485 VSS -0.287f
C1009 vcm.n486 VSS 0.331f
C1010 vcm.t36 VSS 7.36f
C1011 vcm.n487 VSS 2.39f
C1012 vcm.n488 VSS -0.379f
C1013 vcm.n489 VSS 0.156f
C1014 vcm.n490 VSS 0.176f
C1015 vcm.n491 VSS 0.193f
C1016 vcm.n492 VSS 0.21f
C1017 vcm.n493 VSS 0.0444f
C1018 vcm.n494 VSS 0.0444f
C1019 vcm.n496 VSS 1.03f
C1020 vcm.n497 VSS 1.03f
C1021 vcm.n498 VSS 0.242f
C1022 vcm.n499 VSS 0.328f
C1023 vcm.t37 VSS 7.36f
C1024 vcm.n500 VSS 2.39f
C1025 vcm.n501 VSS 2.37f
C1026 vcm.t29 VSS 7.36f
C1027 vcm.n502 VSS 2.37f
C1028 vcm.t21 VSS 7.36f
C1029 vcm.n503 VSS 2.37f
C1030 vcm.n504 VSS 2.37f
C1031 vcm.n505 VSS 0.502f
C1032 vcm.n506 VSS 2.37f
C1033 vcm.n507 VSS 0.251f
C1034 vcm.n508 VSS 0.0569f
C1035 vcm.n509 VSS -0.398f
C1036 vcm.n510 VSS 0.403f
C1037 vcm.n511 VSS -0.0296f
C1038 vcm.n512 VSS -0.34f
C1039 vcm.n513 VSS -0.287f
C1040 vcm.n514 VSS -0.356f
C1041 vcm.t5 VSS 7.36f
C1042 vcm.n515 VSS 2.37f
C1043 vcm.n516 VSS 1f
C1044 vcm.n517 VSS 0.158f
C1045 vcm.n518 VSS 0.241f
C1046 vcm.n519 VSS 0.241f
C1047 vcm.n520 VSS -0.356f
C1048 vcm.n521 VSS 0.403f
C1049 vcm.n522 VSS -0.0297f
C1050 vcm.n523 VSS -0.34f
C1051 vcm.n524 VSS -0.287f
C1052 vcm.n525 VSS -0.356f
C1053 vcm.t13 VSS 7.36f
C1054 vcm.n526 VSS 2.37f
C1055 vcm.n527 VSS 1f
C1056 vcm.n528 VSS 0.158f
C1057 vcm.n529 VSS 0.241f
C1058 vcm.n530 VSS 0.241f
C1059 vcm.n531 VSS -0.356f
C1060 vcm.n532 VSS 0.403f
C1061 vcm.n533 VSS -0.0297f
C1062 vcm.n534 VSS -0.34f
C1063 vcm.n535 VSS -0.287f
C1064 vcm.n536 VSS -0.356f
C1065 vcm.n537 VSS 2.37f
C1066 vcm.n538 VSS 1f
C1067 vcm.n539 VSS 0.158f
C1068 vcm.n540 VSS 0.241f
C1069 vcm.n541 VSS 0.241f
C1070 vcm.n542 VSS -0.356f
C1071 vcm.n543 VSS 0.403f
C1072 vcm.n544 VSS -0.0297f
C1073 vcm.n545 VSS -0.34f
C1074 vcm.n546 VSS -0.287f
C1075 vcm.n547 VSS -0.356f
C1076 vcm.n548 VSS 2.37f
C1077 vcm.n549 VSS 1f
C1078 vcm.n550 VSS 0.158f
C1079 vcm.n551 VSS 0.241f
C1080 vcm.n552 VSS 0.241f
C1081 vcm.n553 VSS -0.356f
C1082 vcm.n554 VSS 0.403f
C1083 vcm.n555 VSS -0.0296f
C1084 vcm.n556 VSS -0.34f
C1085 vcm.n557 VSS -0.287f
C1086 vcm.n558 VSS -0.398f
C1087 vcm.n559 VSS 0.0567f
C1088 vcm.n560 VSS 0.19f
C1089 vcm.n561 VSS 0.21f
C1090 vcm.n562 VSS 0.0444f
C1091 vcm.n563 VSS 0.0444f
C1092 vcm.n565 VSS 0.0526f
C1093 vcm.n566 VSS 0.0393f
C1094 vcm.n567 VSS 0.0393f
C1095 vcm.n569 VSS 0.146f
C1096 vcm.n571 VSS 0.949f
C1097 vcm.n572 VSS 0.949f
C1098 vcm.n573 VSS 0.146f
C1099 vcm.n575 VSS 0.0526f
C1100 vcm.n576 VSS 0.0393f
C1101 vcm.n577 VSS 0.0393f
C1102 vcm.t38 VSS 7.36f
C1103 vcm.n578 VSS 0.403f
C1104 vcm.n579 VSS -0.0297f
C1105 vcm.n580 VSS -0.34f
C1106 vcm.n581 VSS 0.403f
C1107 vcm.n582 VSS -0.0296f
C1108 vcm.n583 VSS -0.34f
C1109 vcm.n584 VSS 2.37f
C1110 vcm.n585 VSS 2.37f
C1111 vcm.t22 VSS 7.36f
C1112 vcm.n586 VSS 0.403f
C1113 vcm.n587 VSS -0.0297f
C1114 vcm.n588 VSS -0.34f
C1115 vcm.n589 VSS 0.403f
C1116 vcm.n590 VSS -0.0296f
C1117 vcm.n591 VSS -0.34f
C1118 vcm.n592 VSS 2.37f
C1119 vcm.n593 VSS 2.37f
C1120 vcm.t6 VSS 7.36f
C1121 vcm.n594 VSS 0.502f
C1122 vcm.n595 VSS 2.37f
C1123 vcm.n596 VSS 0.251f
C1124 vcm.n597 VSS 0.0569f
C1125 vcm.n598 VSS -0.398f
C1126 vcm.n599 VSS 0.403f
C1127 vcm.n600 VSS -0.0296f
C1128 vcm.n601 VSS -0.34f
C1129 vcm.n602 VSS 0.403f
C1130 vcm.n603 VSS -0.0297f
C1131 vcm.n604 VSS -0.34f
C1132 vcm.n605 VSS -0.287f
C1133 vcm.n606 VSS -0.356f
C1134 vcm.n607 VSS 2.37f
C1135 vcm.n608 VSS 1f
C1136 vcm.n609 VSS 0.158f
C1137 vcm.n610 VSS 0.241f
C1138 vcm.n611 VSS 0.241f
C1139 vcm.n612 VSS -0.356f
C1140 vcm.n613 VSS 0.403f
C1141 vcm.n614 VSS -0.0296f
C1142 vcm.n615 VSS -0.34f
C1143 vcm.n616 VSS 0.403f
C1144 vcm.n617 VSS -0.0296f
C1145 vcm.n618 VSS -0.34f
C1146 vcm.n619 VSS -0.287f
C1147 vcm.n620 VSS -0.356f
C1148 vcm.t14 VSS 7.36f
C1149 vcm.n621 VSS 2.37f
C1150 vcm.n622 VSS 1f
C1151 vcm.n623 VSS 0.158f
C1152 vcm.n624 VSS 0.241f
C1153 vcm.n625 VSS 0.241f
C1154 vcm.n626 VSS -0.356f
C1155 vcm.n627 VSS -0.287f
C1156 vcm.n628 VSS -0.356f
C1157 vcm.n629 VSS 2.37f
C1158 vcm.n630 VSS 1f
C1159 vcm.n631 VSS 0.158f
C1160 vcm.n632 VSS 0.241f
C1161 vcm.n633 VSS 0.241f
C1162 vcm.n634 VSS -0.356f
C1163 vcm.n635 VSS 0.403f
C1164 vcm.n636 VSS -0.0296f
C1165 vcm.n637 VSS -0.34f
C1166 vcm.n638 VSS 0.403f
C1167 vcm.n639 VSS -0.0296f
C1168 vcm.n640 VSS -0.34f
C1169 vcm.n641 VSS -0.287f
C1170 vcm.n642 VSS -0.356f
C1171 vcm.t30 VSS 7.36f
C1172 vcm.n643 VSS 2.37f
C1173 vcm.n644 VSS 1f
C1174 vcm.n645 VSS 0.158f
C1175 vcm.n646 VSS 0.241f
C1176 vcm.n647 VSS 0.241f
C1177 vcm.n648 VSS -0.356f
C1178 vcm.n649 VSS -0.287f
C1179 vcm.n650 VSS -0.379f
C1180 vcm.n651 VSS 2.37f
C1181 vcm.n652 VSS 0.503f
C1182 vcm.n653 VSS 0.193f
C1183 vcm.n654 VSS 0.174f
C1184 vcm.n655 VSS 0.184f
C1185 vcm.n656 VSS 0.21f
C1186 vcm.n657 VSS 0.0444f
C1187 vcm.n658 VSS 0.0444f
C1188 vcm.n660 VSS 1.04f
C1189 vcm.n661 VSS 1.04f
C1190 vcm.n662 VSS 0.156f
C1191 vcm.n663 VSS 2.37f
C1192 vcm.t31 VSS 7.36f
C1193 vcm.n664 VSS 0.0142f
C1194 vcm.n665 VSS 2.37f
C1195 vcm.n666 VSS 2.37f
C1196 vcm.t15 VSS 7.36f
C1197 vcm.n667 VSS 0.0142f
C1198 vcm.n668 VSS 2.37f
C1199 vcm.n669 VSS 0.502f
C1200 vcm.n670 VSS 2.37f
C1201 vcm.n671 VSS 0.251f
C1202 vcm.n672 VSS 0.0569f
C1203 vcm.n673 VSS -0.398f
C1204 vcm.n674 VSS 0.13f
C1205 vcm.n675 VSS 3.19f
C1206 vcm.n676 VSS 0.188f
C1207 vcm.n677 VSS -0.135f
C1208 vcm.n678 VSS -0.287f
C1209 vcm.n679 VSS -0.356f
C1210 vcm.t7 VSS 7.36f
C1211 vcm.n680 VSS 2.37f
C1212 vcm.n681 VSS 1f
C1213 vcm.n682 VSS 0.158f
C1214 vcm.n683 VSS 0.241f
C1215 vcm.n684 VSS 0.241f
C1216 vcm.n685 VSS -0.356f
C1217 vcm.n686 VSS -0.287f
C1218 vcm.n687 VSS -0.356f
C1219 vcm.n688 VSS 2.37f
C1220 vcm.n689 VSS 1f
C1221 vcm.n690 VSS 0.158f
C1222 vcm.n691 VSS 0.241f
C1223 vcm.n692 VSS 0.241f
C1224 vcm.n693 VSS -0.356f
C1225 vcm.n694 VSS 0.0139f
C1226 vcm.n695 VSS -0.287f
C1227 vcm.n696 VSS -0.356f
C1228 vcm.t23 VSS 7.36f
C1229 vcm.n697 VSS 2.37f
C1230 vcm.n698 VSS 1f
C1231 vcm.n699 VSS 0.158f
C1232 vcm.n700 VSS 0.241f
C1233 vcm.n701 VSS 0.241f
C1234 vcm.n702 VSS -0.356f
C1235 vcm.n703 VSS -0.287f
C1236 vcm.n704 VSS -0.356f
C1237 vcm.n705 VSS 2.37f
C1238 vcm.n706 VSS 1f
C1239 vcm.n707 VSS 0.158f
C1240 vcm.n708 VSS 0.241f
C1241 vcm.n709 VSS 0.241f
C1242 vcm.n710 VSS -0.356f
C1243 vcm.n711 VSS 0.0139f
C1244 vcm.n712 VSS -0.287f
C1245 vcm.n713 VSS -0.379f
C1246 vcm.t39 VSS 7.36f
C1247 vcm.n714 VSS 2.39f
C1248 vcm.n715 VSS 0.33f
C1249 vcm.n716 VSS 0.177f
C1250 vcm.n717 VSS 0.194f
C1251 vcm.n718 VSS 0.21f
C1252 vcm.n719 VSS 0.0444f
C1253 vcm.n720 VSS 0.0444f
C1254 vcm.n722 VSS 0.0526f
C1255 vcm.n723 VSS 0.0393f
C1256 vcm.n724 VSS 0.0393f
C1257 vcm.n726 VSS 0.146f
C1258 vcm.n728 VSS 1.71f
C1259 vcm.n729 VSS 4.35f
C1260 vcm.n730 VSS 2.57f
C1261 vcm.n731 VSS 0.146f
C1262 vcm.n733 VSS 0.0526f
C1263 vcm.n734 VSS 0.0393f
C1264 vcm.n735 VSS 0.0393f
C1265 vcm.n736 VSS 0.504f
C1266 vcm.t72 VSS 7.36f
C1267 vcm.n737 VSS 2.37f
C1268 vcm.n738 VSS 2.37f
C1269 vcm.t64 VSS 7.36f
C1270 vcm.n739 VSS 0.0144f
C1271 vcm.n740 VSS 2.37f
C1272 vcm.t56 VSS 7.36f
C1273 vcm.n741 VSS 0.0144f
C1274 vcm.n742 VSS 2.37f
C1275 vcm.n743 VSS 2.37f
C1276 vcm.t40 VSS 7.36f
C1277 vcm.n744 VSS 0.502f
C1278 vcm.n745 VSS 2.37f
C1279 vcm.n746 VSS 0.251f
C1280 vcm.n747 VSS 0.0569f
C1281 vcm.n748 VSS -0.398f
C1282 vcm.n749 VSS 0.196f
C1283 vcm.n750 VSS 0.078f
C1284 vcm.n751 VSS 0.0766f
C1285 vcm.n752 VSS 3.43f
C1286 vcm.n753 VSS -0.473f
C1287 vcm.n754 VSS 0.0143f
C1288 vcm.n755 VSS 0.0451f
C1289 vcm.n756 VSS -0.177f
C1290 vcm.n757 VSS -0.287f
C1291 vcm.n758 VSS -0.356f
C1292 vcm.n759 VSS 2.37f
C1293 vcm.n760 VSS 1f
C1294 vcm.n761 VSS 0.158f
C1295 vcm.n762 VSS 0.241f
C1296 vcm.n763 VSS 0.241f
C1297 vcm.n764 VSS -0.356f
C1298 vcm.n765 VSS 0.0144f
C1299 vcm.n766 VSS -0.288f
C1300 vcm.n767 VSS -0.356f
C1301 vcm.t48 VSS 7.36f
C1302 vcm.n768 VSS 2.37f
C1303 vcm.n769 VSS 1f
C1304 vcm.n770 VSS 0.158f
C1305 vcm.n771 VSS 0.241f
C1306 vcm.n772 VSS 0.241f
C1307 vcm.n773 VSS -0.356f
C1308 vcm.n774 VSS -0.288f
C1309 vcm.n775 VSS -0.356f
C1310 vcm.n776 VSS 2.37f
C1311 vcm.n777 VSS 1f
C1312 vcm.n778 VSS 0.158f
C1313 vcm.n779 VSS 0.241f
C1314 vcm.n780 VSS 0.241f
C1315 vcm.n781 VSS -0.356f
C1316 vcm.n782 VSS -0.288f
C1317 vcm.n783 VSS -0.356f
C1318 vcm.n784 VSS 2.37f
C1319 vcm.n785 VSS 1f
C1320 vcm.n786 VSS 0.149f
C1321 vcm.n787 VSS 0.243f
C1322 vcm.n788 VSS 0.248f
C1323 vcm.n789 VSS -0.356f
C1324 vcm.n790 VSS 0.0144f
C1325 vcm.n791 VSS -0.288f
C1326 vcm.n792 VSS -0.379f
C1327 vcm.n793 VSS 0.193f
C1328 vcm.n794 VSS 0.173f
C1329 vcm.n795 VSS 0.184f
C1330 vcm.n796 VSS 0.21f
C1331 vcm.n797 VSS 0.0444f
C1332 vcm.n798 VSS 0.0444f
C1333 vcm.n800 VSS 1.07f
C1334 vcm.n801 VSS 1.07f
C1335 vcm.n802 VSS 0.242f
C1336 vcm.n803 VSS 0.329f
C1337 vcm.t73 VSS 7.36f
C1338 vcm.n804 VSS 2.39f
C1339 vcm.n805 VSS 2.37f
C1340 vcm.t65 VSS 7.36f
C1341 vcm.n806 VSS 2.37f
C1342 vcm.t57 VSS 7.36f
C1343 vcm.n807 VSS 2.37f
C1344 vcm.t49 VSS 7.36f
C1345 vcm.n808 VSS 0.404f
C1346 vcm.n809 VSS -0.0314f
C1347 vcm.n810 VSS -0.341f
C1348 vcm.n811 VSS 0.427f
C1349 vcm.n812 VSS -0.0315f
C1350 vcm.n813 VSS -0.364f
C1351 vcm.n814 VSS 2.37f
C1352 vcm.n815 VSS 0.502f
C1353 vcm.n816 VSS 2.37f
C1354 vcm.n817 VSS 0.251f
C1355 vcm.n818 VSS 0.0569f
C1356 vcm.n819 VSS -0.398f
C1357 vcm.n820 VSS 0.403f
C1358 vcm.n821 VSS -0.0296f
C1359 vcm.n822 VSS -0.34f
C1360 vcm.n823 VSS 0.403f
C1361 vcm.n824 VSS -0.0296f
C1362 vcm.n825 VSS -0.34f
C1363 vcm.n826 VSS -0.287f
C1364 vcm.n827 VSS -0.356f
C1365 vcm.t41 VSS 7.36f
C1366 vcm.n828 VSS 2.37f
C1367 vcm.n829 VSS 1f
C1368 vcm.n830 VSS 0.158f
C1369 vcm.n831 VSS 0.241f
C1370 vcm.n832 VSS 0.241f
C1371 vcm.n833 VSS -0.356f
C1372 vcm.n834 VSS -0.287f
C1373 vcm.n835 VSS -0.356f
C1374 vcm.n836 VSS 2.37f
C1375 vcm.n837 VSS 1f
C1376 vcm.n838 VSS 0.158f
C1377 vcm.n839 VSS 0.241f
C1378 vcm.n840 VSS 0.241f
C1379 vcm.n841 VSS -0.356f
C1380 vcm.n842 VSS 0.403f
C1381 vcm.n843 VSS -0.0296f
C1382 vcm.n844 VSS -0.34f
C1383 vcm.n845 VSS 0.404f
C1384 vcm.n846 VSS -0.0314f
C1385 vcm.n847 VSS -0.341f
C1386 vcm.n848 VSS -0.287f
C1387 vcm.n849 VSS -0.356f
C1388 vcm.n850 VSS 2.37f
C1389 vcm.n851 VSS 1f
C1390 vcm.n852 VSS 0.149f
C1391 vcm.n853 VSS 0.243f
C1392 vcm.n854 VSS 0.248f
C1393 vcm.n855 VSS -0.356f
C1394 vcm.n856 VSS 0.403f
C1395 vcm.n857 VSS -0.0296f
C1396 vcm.n858 VSS -0.34f
C1397 vcm.n859 VSS 0.403f
C1398 vcm.n860 VSS -0.0297f
C1399 vcm.n861 VSS -0.34f
C1400 vcm.n862 VSS -0.287f
C1401 vcm.n863 VSS -0.356f
C1402 vcm.n864 VSS 2.37f
C1403 vcm.n865 VSS 1f
C1404 vcm.n866 VSS 0.158f
C1405 vcm.n867 VSS 0.241f
C1406 vcm.n868 VSS 0.241f
C1407 vcm.n869 VSS -0.356f
C1408 vcm.n870 VSS 0.426f
C1409 vcm.n871 VSS -0.0315f
C1410 vcm.n872 VSS -0.364f
C1411 vcm.n873 VSS 0.404f
C1412 vcm.n874 VSS -0.0314f
C1413 vcm.n875 VSS -0.341f
C1414 vcm.n876 VSS -0.287f
C1415 vcm.n877 VSS -0.398f
C1416 vcm.n878 VSS 0.0562f
C1417 vcm.n879 VSS 0.189f
C1418 vcm.n880 VSS 0.21f
C1419 vcm.n881 VSS 0.0444f
C1420 vcm.n882 VSS 0.0444f
C1421 vcm.n884 VSS 0.0526f
C1422 vcm.n885 VSS 0.0393f
C1423 vcm.n886 VSS 0.0393f
C1424 vcm.n888 VSS 0.146f
C1425 vcm.n890 VSS 0.982f
C1426 vcm.n891 VSS 0.982f
C1427 vcm.n892 VSS 0.146f
C1428 vcm.n894 VSS 0.0526f
C1429 vcm.n895 VSS 0.0393f
C1430 vcm.n896 VSS 0.0393f
C1431 vcm.n897 VSS 0.331f
C1432 vcm.t74 VSS 7.36f
C1433 vcm.n898 VSS 2.39f
C1434 vcm.n899 VSS 2.37f
C1435 vcm.t66 VSS 7.36f
C1436 vcm.n900 VSS 2.37f
C1437 vcm.t58 VSS 7.36f
C1438 vcm.n901 VSS 2.37f
C1439 vcm.t50 VSS 7.36f
C1440 vcm.n902 VSS 2.37f
C1441 vcm.t42 VSS 7.36f
C1442 vcm.n903 VSS 0.502f
C1443 vcm.n904 VSS 2.37f
C1444 vcm.n905 VSS 0.251f
C1445 vcm.n906 VSS 0.0569f
C1446 vcm.n907 VSS -0.398f
C1447 vcm.n908 VSS -0.287f
C1448 vcm.n909 VSS -0.356f
C1449 vcm.n910 VSS 2.37f
C1450 vcm.n911 VSS 1f
C1451 vcm.n912 VSS 0.158f
C1452 vcm.n913 VSS 0.241f
C1453 vcm.n914 VSS 0.241f
C1454 vcm.n915 VSS -0.356f
C1455 vcm.n916 VSS -0.287f
C1456 vcm.n917 VSS -0.356f
C1457 vcm.n918 VSS 2.37f
C1458 vcm.n919 VSS 1f
C1459 vcm.n920 VSS 0.149f
C1460 vcm.n921 VSS 0.243f
C1461 vcm.n922 VSS 0.248f
C1462 vcm.n923 VSS -0.356f
C1463 vcm.n924 VSS -0.287f
C1464 vcm.n925 VSS -0.356f
C1465 vcm.n926 VSS 2.37f
C1466 vcm.n927 VSS 1f
C1467 vcm.n928 VSS 0.158f
C1468 vcm.n929 VSS 0.241f
C1469 vcm.n930 VSS 0.241f
C1470 vcm.n931 VSS -0.356f
C1471 vcm.n932 VSS -0.287f
C1472 vcm.n933 VSS -0.356f
C1473 vcm.n934 VSS 2.37f
C1474 vcm.n935 VSS 1f
C1475 vcm.n936 VSS 0.158f
C1476 vcm.n937 VSS 0.241f
C1477 vcm.n938 VSS 0.241f
C1478 vcm.n939 VSS -0.356f
C1479 vcm.n940 VSS -0.287f
C1480 vcm.n941 VSS -0.379f
C1481 vcm.n942 VSS 0.156f
C1482 vcm.n943 VSS 0.176f
C1483 vcm.n944 VSS 0.193f
C1484 vcm.n945 VSS 0.21f
C1485 vcm.n946 VSS 0.0444f
C1486 vcm.n947 VSS 0.0444f
C1487 vcm.n949 VSS 1.01f
C1488 vcm.n950 VSS 1.01f
C1489 vcm.n951 VSS 0.146f
C1490 vcm.n953 VSS 0.331f
C1491 vcm.t75 VSS 7.36f
C1492 vcm.n954 VSS 2.39f
C1493 vcm.n955 VSS 2.37f
C1494 vcm.t67 VSS 7.36f
C1495 vcm.n956 VSS 2.37f
C1496 vcm.t59 VSS 7.36f
C1497 vcm.n957 VSS 0.403f
C1498 vcm.n958 VSS -0.0296f
C1499 vcm.n959 VSS -0.34f
C1500 vcm.n960 VSS 2.37f
C1501 vcm.n961 VSS 2.37f
C1502 vcm.t43 VSS 7.36f
C1503 vcm.n962 VSS 0.502f
C1504 vcm.n963 VSS 2.37f
C1505 vcm.n964 VSS 0.251f
C1506 vcm.n965 VSS 0.0569f
C1507 vcm.n966 VSS -0.398f
C1508 vcm.n967 VSS 0.403f
C1509 vcm.n968 VSS -0.0297f
C1510 vcm.n969 VSS -0.34f
C1511 vcm.n970 VSS -0.287f
C1512 vcm.n971 VSS -0.356f
C1513 vcm.n972 VSS 2.37f
C1514 vcm.n973 VSS 1f
C1515 vcm.n974 VSS 0.149f
C1516 vcm.n975 VSS 0.243f
C1517 vcm.n976 VSS 0.248f
C1518 vcm.n977 VSS -0.356f
C1519 vcm.n978 VSS 0.403f
C1520 vcm.n979 VSS -0.0296f
C1521 vcm.n980 VSS -0.34f
C1522 vcm.n981 VSS -0.287f
C1523 vcm.n982 VSS -0.356f
C1524 vcm.t51 VSS 7.36f
C1525 vcm.n983 VSS 2.37f
C1526 vcm.n984 VSS 1f
C1527 vcm.n985 VSS 0.158f
C1528 vcm.n986 VSS 0.241f
C1529 vcm.n987 VSS 0.241f
C1530 vcm.n988 VSS -0.356f
C1531 vcm.n989 VSS -0.287f
C1532 vcm.n990 VSS -0.356f
C1533 vcm.n991 VSS 2.37f
C1534 vcm.n992 VSS 1f
C1535 vcm.n993 VSS 0.158f
C1536 vcm.n994 VSS 0.241f
C1537 vcm.n995 VSS 0.241f
C1538 vcm.n996 VSS -0.356f
C1539 vcm.n997 VSS 0.403f
C1540 vcm.n998 VSS -0.0296f
C1541 vcm.n999 VSS -0.34f
C1542 vcm.n1000 VSS -0.287f
C1543 vcm.n1001 VSS -0.356f
C1544 vcm.n1002 VSS 2.37f
C1545 vcm.n1003 VSS 1f
C1546 vcm.n1004 VSS 0.158f
C1547 vcm.n1005 VSS 0.241f
C1548 vcm.n1006 VSS 0.241f
C1549 vcm.n1007 VSS -0.356f
C1550 vcm.n1008 VSS 0.404f
C1551 vcm.n1009 VSS -0.0314f
C1552 vcm.n1010 VSS -0.341f
C1553 vcm.n1011 VSS -0.287f
C1554 vcm.n1012 VSS -0.379f
C1555 vcm.n1013 VSS 0.156f
C1556 vcm.n1014 VSS 0.177f
C1557 vcm.n1015 VSS 0.194f
C1558 vcm.n1016 VSS 0.21f
C1559 vcm.n1017 VSS 0.0444f
C1560 vcm.n1018 VSS 0.0444f
C1561 vcm.n1020 VSS 0.992f
C1562 vcm.t76 VSS 7.36f
C1563 vcm.n1021 VSS 0.176f
C1564 vcm.n1022 VSS 0.193f
C1565 vcm.n1023 VSS 0.426f
C1566 vcm.n1024 VSS -0.0315f
C1567 vcm.n1025 VSS -0.364f
C1568 vcm.n1026 VSS 2.37f
C1569 vcm.n1027 VSS 2.37f
C1570 vcm.t60 VSS 7.36f
C1571 vcm.n1028 VSS 2.37f
C1572 vcm.t52 VSS 7.36f
C1573 vcm.n1029 VSS 0.403f
C1574 vcm.n1030 VSS -0.0296f
C1575 vcm.n1031 VSS -0.34f
C1576 vcm.n1032 VSS 2.37f
C1577 vcm.n1033 VSS 0.502f
C1578 vcm.n1034 VSS 2.37f
C1579 vcm.n1035 VSS 0.251f
C1580 vcm.n1036 VSS 0.0569f
C1581 vcm.n1037 VSS -0.398f
C1582 vcm.n1038 VSS 0.404f
C1583 vcm.n1039 VSS -0.0314f
C1584 vcm.n1040 VSS -0.341f
C1585 vcm.n1041 VSS -0.287f
C1586 vcm.n1042 VSS -0.356f
C1587 vcm.t44 VSS 7.36f
C1588 vcm.n1043 VSS 2.37f
C1589 vcm.n1044 VSS 1f
C1590 vcm.n1045 VSS 0.158f
C1591 vcm.n1046 VSS 0.241f
C1592 vcm.n1047 VSS 0.241f
C1593 vcm.n1048 VSS -0.356f
C1594 vcm.n1049 VSS -0.287f
C1595 vcm.n1050 VSS -0.356f
C1596 vcm.n1051 VSS 2.37f
C1597 vcm.n1052 VSS 1f
C1598 vcm.n1053 VSS 0.158f
C1599 vcm.n1054 VSS 0.241f
C1600 vcm.n1055 VSS 0.241f
C1601 vcm.n1056 VSS -0.356f
C1602 vcm.n1057 VSS 0.403f
C1603 vcm.n1058 VSS -0.0297f
C1604 vcm.n1059 VSS -0.34f
C1605 vcm.n1060 VSS -0.287f
C1606 vcm.n1061 VSS -0.356f
C1607 vcm.n1062 VSS 2.37f
C1608 vcm.n1063 VSS 1f
C1609 vcm.n1064 VSS 0.158f
C1610 vcm.n1065 VSS 0.241f
C1611 vcm.n1066 VSS 0.241f
C1612 vcm.n1067 VSS -0.356f
C1613 vcm.n1068 VSS 0.403f
C1614 vcm.n1069 VSS -0.0296f
C1615 vcm.n1070 VSS -0.34f
C1616 vcm.n1071 VSS -0.287f
C1617 vcm.n1072 VSS -0.356f
C1618 vcm.t68 VSS 7.36f
C1619 vcm.n1073 VSS 2.37f
C1620 vcm.n1074 VSS 1f
C1621 vcm.n1075 VSS 0.158f
C1622 vcm.n1076 VSS 0.241f
C1623 vcm.n1077 VSS 0.241f
C1624 vcm.n1078 VSS -0.356f
C1625 vcm.n1079 VSS -0.287f
C1626 vcm.n1080 VSS -0.379f
C1627 vcm.n1081 VSS 2.37f
C1628 vcm.n1082 VSS 0.501f
C1629 vcm.n1083 VSS 0.184f
C1630 vcm.n1084 VSS 0.21f
C1631 vcm.n1085 VSS 0.0444f
C1632 vcm.n1086 VSS 0.0444f
C1633 vcm.n1087 VSS 0.992f
C1634 vcm.n1088 VSS 0.146f
C1635 vcm.n1090 VSS 0.0526f
C1636 vcm.n1091 VSS 0.0393f
C1637 vcm.n1092 VSS 0.0393f
C1638 vcm.n1094 VSS 1f
C1639 vcm.n1095 VSS 1f
C1640 vcm.n1096 VSS 0.146f
C1641 vcm.n1098 VSS 0.0526f
C1642 vcm.n1099 VSS 0.0393f
C1643 vcm.n1100 VSS 0.0393f
C1644 vcm.n1101 VSS 2.37f
C1645 vcm.n1102 VSS 2.37f
C1646 vcm.t61 VSS 7.36f
C1647 vcm.n1103 VSS 2.37f
C1648 vcm.t53 VSS 7.36f
C1649 vcm.n1104 VSS 2.37f
C1650 vcm.t45 VSS 7.36f
C1651 vcm.n1105 VSS 0.502f
C1652 vcm.n1106 VSS 2.37f
C1653 vcm.n1107 VSS 0.251f
C1654 vcm.n1108 VSS 0.0569f
C1655 vcm.n1109 VSS -0.398f
C1656 vcm.n1110 VSS 0.426f
C1657 vcm.n1111 VSS -0.0315f
C1658 vcm.n1112 VSS -0.364f
C1659 vcm.n1113 VSS -0.287f
C1660 vcm.n1114 VSS -0.356f
C1661 vcm.n1115 VSS 2.37f
C1662 vcm.n1116 VSS 1f
C1663 vcm.n1117 VSS 0.158f
C1664 vcm.n1118 VSS 0.241f
C1665 vcm.n1119 VSS 0.241f
C1666 vcm.n1120 VSS -0.356f
C1667 vcm.n1121 VSS 0.403f
C1668 vcm.n1122 VSS -0.0297f
C1669 vcm.n1123 VSS -0.34f
C1670 vcm.n1124 VSS -0.287f
C1671 vcm.n1125 VSS -0.356f
C1672 vcm.n1126 VSS 2.37f
C1673 vcm.n1127 VSS 1f
C1674 vcm.n1128 VSS 0.158f
C1675 vcm.n1129 VSS 0.241f
C1676 vcm.n1130 VSS 0.241f
C1677 vcm.n1131 VSS -0.356f
C1678 vcm.n1132 VSS 0.403f
C1679 vcm.n1133 VSS -0.0297f
C1680 vcm.n1134 VSS -0.34f
C1681 vcm.n1135 VSS -0.287f
C1682 vcm.n1136 VSS -0.356f
C1683 vcm.n1137 VSS 2.37f
C1684 vcm.n1138 VSS 1f
C1685 vcm.n1139 VSS 0.158f
C1686 vcm.n1140 VSS 0.241f
C1687 vcm.n1141 VSS 0.241f
C1688 vcm.n1142 VSS -0.356f
C1689 vcm.n1143 VSS 0.403f
C1690 vcm.n1144 VSS -0.0297f
C1691 vcm.n1145 VSS -0.34f
C1692 vcm.n1146 VSS -0.287f
C1693 vcm.n1147 VSS -0.356f
C1694 vcm.t69 VSS 7.36f
C1695 vcm.n1148 VSS 2.37f
C1696 vcm.n1149 VSS 1f
C1697 vcm.n1150 VSS 0.158f
C1698 vcm.n1151 VSS 0.241f
C1699 vcm.n1152 VSS 0.241f
C1700 vcm.n1153 VSS -0.356f
C1701 vcm.n1154 VSS 0.404f
C1702 vcm.n1155 VSS -0.0314f
C1703 vcm.n1156 VSS -0.341f
C1704 vcm.n1157 VSS -0.287f
C1705 vcm.n1158 VSS 0.176f
C1706 vcm.n1159 VSS 0.193f
C1707 vcm.n1160 VSS -0.379f
C1708 vcm.t77 VSS 7.36f
C1709 vcm.n1161 VSS 2.37f
C1710 vcm.n1162 VSS 0.501f
C1711 vcm.n1163 VSS 0.184f
C1712 vcm.n1164 VSS 0.21f
C1713 vcm.n1165 VSS 0.0444f
C1714 vcm.n1166 VSS 0.0444f
C1715 vcm.n1168 VSS 1f
C1716 vcm.n1169 VSS 1f
C1717 vcm.n1170 VSS 0.146f
C1718 vcm.n1172 VSS 0.331f
C1719 vcm.t78 VSS 7.36f
C1720 vcm.n1173 VSS 2.39f
C1721 vcm.n1174 VSS -0.379f
C1722 vcm.n1175 VSS 0.156f
C1723 vcm.n1176 VSS 0.176f
C1724 vcm.n1177 VSS 0.193f
C1725 vcm.n1178 VSS 0.21f
C1726 vcm.n1179 VSS 0.0444f
C1727 vcm.n1180 VSS 0.0444f
C1728 vcm.n1182 VSS 1f
C1729 vcm.n1183 VSS 1f
C1730 vcm.n1184 VSS 0.0444f
C1731 vcm.n1185 VSS 0.0444f
C1732 vcm.n1186 VSS 0.21f
C1733 vcm.n1187 VSS 0.193f
C1734 vcm.n1188 VSS 0.176f
C1735 VDD.n0 VSS 0.00279f
C1736 VDD.n1 VSS 0.0028f
C1737 VDD.n3 VSS 6.43e-19
C1738 VDD.n4 VSS 0.00406f
C1739 VDD.n5 VSS 0.00253f
C1740 VDD.n6 VSS 0.00406f
C1741 VDD.n7 VSS 6.6e-19
C1742 VDD.n8 VSS 0.00805f
C1743 VDD.n9 VSS 1.92f
C1744 VDD.n10 VSS 0.0034f
C1745 VDD.n11 VSS 6.75e-19
C1746 VDD.n12 VSS 0.00226f
C1747 VDD.n13 VSS 6.75e-19
C1748 VDD.n14 VSS 0.00226f
C1749 VDD.n15 VSS 0.00157f
C1750 VDD.n16 VSS 0.00226f
C1751 VDD.n17 VSS 0.00201f
C1752 VDD.n18 VSS 0.00519f
C1753 VDD.n19 VSS 0.00226f
C1754 VDD.n20 VSS 0.00254f
C1755 VDD.n21 VSS 0.0017f
C1756 VDD.n22 VSS 0.0017f
C1757 VDD.n23 VSS 0.00175f
C1758 VDD.n24 VSS 0.00157f
C1759 VDD.n25 VSS 0.00118f
C1760 VDD.n26 VSS 0.0103f
C1761 VDD.n27 VSS 0.0463f
C1762 VDD.n28 VSS 0.0131f
C1763 VDD.n29 VSS 7.75e-19
C1764 VDD.n30 VSS 0.00356f
C1765 VDD.n31 VSS 0.00424f
C1766 VDD.n32 VSS 0.00205f
C1767 VDD.n33 VSS 0.0017f
C1768 VDD.n34 VSS 7.75e-19
C1769 VDD.n35 VSS 0.00369f
C1770 VDD.n36 VSS 0.00385f
C1771 VDD.n37 VSS 0.00205f
C1772 VDD.n38 VSS 0.0017f
C1773 VDD.n39 VSS 7.87e-19
C1774 VDD.n40 VSS 4.79e-19
C1775 VDD.n41 VSS 0.00587f
C1776 VDD.n42 VSS 0.00204f
C1777 VDD.n43 VSS 0.00226f
C1778 VDD.n44 VSS 0.00139f
C1779 VDD.n45 VSS 0.00656f
C1780 VDD.n46 VSS 7.23e-19
C1781 VDD.n47 VSS 0.00809f
C1782 VDD.n48 VSS 0.0017f
C1783 VDD.n49 VSS 7.87e-19
C1784 VDD.n50 VSS 1.44e-19
C1785 VDD.n51 VSS 0.00567f
C1786 VDD.n52 VSS 0.00204f
C1787 VDD.n53 VSS 0.00226f
C1788 VDD.n54 VSS 0.00226f
C1789 VDD.n55 VSS 0.006f
C1790 VDD.n56 VSS 7.88e-19
C1791 VDD.n57 VSS 0.00804f
C1792 VDD.n58 VSS 0.0017f
C1793 VDD.n59 VSS 9.22e-19
C1794 VDD.n60 VSS 8.24e-19
C1795 VDD.n61 VSS 8.01e-19
C1796 VDD.n62 VSS 8.01e-19
C1797 VDD.n63 VSS 0.0017f
C1798 VDD.n64 VSS 0.00226f
C1799 VDD.n65 VSS 0.00226f
C1800 VDD.n66 VSS 0.00118f
C1801 VDD.n67 VSS 8.01e-19
C1802 VDD.n68 VSS 0.00162f
C1803 VDD.n69 VSS 0.00226f
C1804 VDD.n70 VSS 0.00226f
C1805 VDD.n71 VSS 0.00226f
C1806 VDD.n72 VSS 8.01e-19
C1807 VDD.n73 VSS 0.00112f
C1808 VDD.n74 VSS 0.00961f
C1809 VDD.n75 VSS 0.00226f
C1810 VDD.n76 VSS 0.00139f
C1811 VDD.n77 VSS 0.0017f
C1812 VDD.n78 VSS 0.00673f
C1813 VDD.n79 VSS 5.83e-19
C1814 VDD.n80 VSS 0.00698f
C1815 VDD.n81 VSS 0.00135f
C1816 VDD.n82 VSS 0.0017f
C1817 VDD.n83 VSS 7.75e-19
C1818 VDD.n84 VSS 0.00143f
C1819 VDD.n85 VSS 0.00667f
C1820 VDD.n86 VSS 0.0196f
C1821 VDD.n87 VSS 0.0119f
C1822 VDD.n88 VSS 0.00548f
C1823 VDD.n89 VSS 0.00729f
C1824 VDD.n90 VSS 8.61e-19
C1825 VDD.n91 VSS 0.0141f
C1826 VDD.n92 VSS 0.00279f
C1827 VDD.n93 VSS 0.0028f
C1828 VDD.n94 VSS 0.0028f
C1829 VDD.n95 VSS 6.75e-19
C1830 VDD.n96 VSS 0.00209f
C1831 VDD.n97 VSS 0.0537f
C1832 VDD.n98 VSS 0.00804f
C1833 VDD.n99 VSS 0.00244f
C1834 VDD.n101 VSS 0.00118f
C1835 VDD.n102 VSS 0.00248f
C1836 VDD.n103 VSS 0.00356f
C1837 VDD.n104 VSS 0.00408f
C1838 VDD.n105 VSS 0.00408f
C1839 VDD.n106 VSS 0.00408f
C1840 VDD.n107 VSS 3.73f
C1841 VDD.n108 VSS 0.00408f
C1842 VDD.n109 VSS 0.00408f
C1843 VDD.n110 VSS 0.00408f
C1844 VDD.n111 VSS 1.77f
C1845 VDD.n112 VSS 0.00408f
C1846 VDD.n113 VSS 0.00408f
C1847 VDD.n114 VSS 0.00408f
C1848 VDD.n115 VSS 0.00408f
C1849 VDD.n116 VSS 0.00408f
C1850 VDD.n117 VSS 0.0045f
C1851 VDD.n118 VSS 0.00408f
C1852 VDD.n119 VSS 0.00418f
C1853 VDD.n120 VSS 0.00408f
C1854 VDD.n121 VSS 0.00408f
C1855 VDD.n122 VSS 0.00408f
C1856 VDD.n123 VSS 0.00408f
C1857 VDD.n124 VSS 0.00511f
C1858 VDD.n125 VSS 0.0585f
C1859 VDD.n126 VSS 0.00133f
C1860 VDD.n127 VSS -0.0588f
C1861 VDD.n128 VSS 0.205f
C1862 VDD.n129 VSS 0.00133f
C1863 VDD.n130 VSS -0.0588f
C1864 VDD.n131 VSS 0.205f
C1865 VDD.n132 VSS 0.00133f
C1866 VDD.n133 VSS -0.0588f
C1867 VDD.n134 VSS 0.103f
C1868 VDD.n135 VSS 0.0512f
C1869 VDD.n136 VSS 0.0116f
C1870 VDD.n137 VSS -0.0814f
C1871 VDD.n138 VSS 0.484f
C1872 VDD.t0 VSS 1.51f
C1873 VDD.n139 VSS 0.484f
C1874 VDD.n140 VSS -0.0729f
C1875 VDD.n141 VSS 0.0304f
C1876 VDD.n142 VSS 0.0498f
C1877 VDD.n143 VSS 0.0508f
C1878 VDD.n144 VSS -0.0729f
C1879 VDD.n145 VSS 0.484f
C1880 VDD.t2 VSS 1.51f
C1881 VDD.n146 VSS 0.484f
C1882 VDD.n147 VSS -0.0729f
C1883 VDD.n148 VSS 0.0304f
C1884 VDD.n149 VSS 0.0498f
C1885 VDD.n150 VSS 0.0508f
C1886 VDD.n151 VSS -0.0729f
C1887 VDD.n152 VSS 0.484f
C1888 VDD.t4 VSS 1.51f
C1889 VDD.n153 VSS 0.488f
C1890 VDD.n154 VSS -0.0814f
C1891 VDD.n155 VSS 0.0115f
C1892 VDD.n156 VSS 0.0427f
C1893 VDD.n157 VSS 0.0151f
C1894 VDD.n158 VSS 0.00408f
C1895 VDD.n159 VSS 0.00238f
C1896 VDD.n160 VSS 0.0316f
C1897 VDD.t5 VSS 4.74f
C1898 VDD.t3 VSS 4.74f
C1899 VDD.t1 VSS 5.4f
C1900 VDD.n161 VSS 1.71f
C1901 VDD.n162 VSS 1.71f
C1902 VDD.n163 VSS 0.759f
C1903 VDD.n164 VSS 0.038f
C1904 VDD.n165 VSS 0.0512f
C1905 VDD.n166 VSS 0.00516f
C1906 VDD.n167 VSS 0.00532f
C1907 VDD.n168 VSS 0.00238f
C1908 VDD.n169 VSS 0.00408f
C1909 VDD.n170 VSS 0.00408f
C1910 VDD.n171 VSS 0.00408f
C1911 VDD.n172 VSS 0.00408f
C1912 VDD.n173 VSS 0.00408f
C1913 VDD.n174 VSS 0.00408f
C1914 VDD.n175 VSS 0.00408f
C1915 VDD.n176 VSS 0.0147f
C1916 VDD.n177 VSS 0.0237f
C1917 VDD.n178 VSS 0.0237f
C1918 VDD.n179 VSS 0.00474f
C1919 VDD.n180 VSS 0.00474f
C1920 VDD.n181 VSS 0.00408f
C1921 VDD.n182 VSS 0.00408f
C1922 VDD.n183 VSS 0.00408f
C1923 VDD.n184 VSS 0.00408f
C1924 VDD.n185 VSS 0.00412f
C1925 VDD.n186 VSS 0.00417f
C1926 VDD.n187 VSS 0.0151f
C1927 VDD.n188 VSS 0.259f
C1928 VDD.n189 VSS 0.00408f
C1929 VDD.n190 VSS 0.00408f
C1930 VDD.n191 VSS 0.0151f
C1931 VDD.n192 VSS 0.00408f
C1932 VDD.n193 VSS 0.00417f
C1933 VDD.n194 VSS 0.00412f
C1934 VDD.n195 VSS 0.00408f
C1935 VDD.n196 VSS 0.00408f
C1936 VDD.n197 VSS 0.00408f
C1937 VDD.n198 VSS 0.259f
C1938 VDD.n199 VSS 0.00474f
C1939 VDD.n200 VSS 0.00474f
C1940 VDD.n201 VSS 0.694f
C1941 VDD.n202 VSS 0.698f
C1942 VDD.n203 VSS 0.00359f
C1943 VDD.n204 VSS 0.00247f
C1944 VDD.n205 VSS 0.00694f
C1945 VDD.n206 VSS 0.00694f
C1946 VDD.n207 VSS 0.00359f
C1947 VDD.n208 VSS 0.00115f
C1948 VDD.n209 VSS 0.00115f
C1949 VDD.n210 VSS 0.00816f
C1950 VDD.n211 VSS 0.01f
C1951 VDD.n212 VSS 0.00108f
C1952 VDD.n214 VSS 3.72f
C1953 VDD.n215 VSS 0.00811f
C1954 VDD.n216 VSS 0.0571f
C1955 VDD.n217 VSS 0.0537f
C1956 VDD.n218 VSS 6.5e-19
C1957 VDD.n219 VSS 0.00188f
C1958 VDD.n220 VSS 0.0537f
C1959 VDD.n221 VSS 0.0028f
C1960 VDD.n222 VSS 0.0028f
C1961 VDD.n223 VSS 0.015f
C1962 VDD.n224 VSS 0.0066f
C1963 VDD.n225 VSS 7.62e-19
C1964 VDD.n226 VSS 0.00519f
C1965 VDD.n227 VSS 0.0017f
C1966 VDD.n228 VSS 0.0017f
C1967 VDD.n229 VSS 0.00175f
C1968 VDD.n230 VSS 0.00157f
C1969 VDD.n231 VSS 0.00118f
C1970 VDD.n232 VSS 0.0484f
C1971 VDD.n233 VSS 0.0131f
C1972 VDD.n234 VSS 7.75e-19
C1973 VDD.n235 VSS 0.00356f
C1974 VDD.n236 VSS 0.00424f
C1975 VDD.n237 VSS 0.00205f
C1976 VDD.n238 VSS 0.0017f
C1977 VDD.n239 VSS 7.75e-19
C1978 VDD.n240 VSS 0.00369f
C1979 VDD.n241 VSS 0.00385f
C1980 VDD.n242 VSS 0.00205f
C1981 VDD.n243 VSS 0.0017f
C1982 VDD.n244 VSS 7.87e-19
C1983 VDD.n245 VSS 4.79e-19
C1984 VDD.n246 VSS 0.00587f
C1985 VDD.n247 VSS 0.00204f
C1986 VDD.n248 VSS 0.00226f
C1987 VDD.n249 VSS 0.00139f
C1988 VDD.n250 VSS 0.00656f
C1989 VDD.n251 VSS 7.23e-19
C1990 VDD.n252 VSS 0.00809f
C1991 VDD.n253 VSS 0.0017f
C1992 VDD.n254 VSS 7.87e-19
C1993 VDD.n255 VSS 1.44e-19
C1994 VDD.n256 VSS 0.00567f
C1995 VDD.n257 VSS 0.00204f
C1996 VDD.n258 VSS 0.00254f
C1997 VDD.n259 VSS 0.00226f
C1998 VDD.n260 VSS 0.006f
C1999 VDD.n261 VSS 0.00226f
C2000 VDD.n262 VSS 7.88e-19
C2001 VDD.n263 VSS 0.00226f
C2002 VDD.n264 VSS 0.00804f
C2003 VDD.n265 VSS 0.0017f
C2004 VDD.n266 VSS 9.22e-19
C2005 VDD.n267 VSS 8.24e-19
C2006 VDD.n268 VSS 8.01e-19
C2007 VDD.n269 VSS 8.01e-19
C2008 VDD.n270 VSS 0.0017f
C2009 VDD.n271 VSS 0.00201f
C2010 VDD.n272 VSS 0.00226f
C2011 VDD.n273 VSS 0.00118f
C2012 VDD.n274 VSS 0.00226f
C2013 VDD.n275 VSS 8.01e-19
C2014 VDD.n276 VSS 0.00226f
C2015 VDD.n277 VSS 0.00162f
C2016 VDD.n278 VSS 0.00226f
C2017 VDD.n279 VSS 0.00157f
C2018 VDD.n280 VSS 0.00226f
C2019 VDD.n281 VSS 8.01e-19
C2020 VDD.n282 VSS 0.00226f
C2021 VDD.n283 VSS 0.00123f
C2022 VDD.n284 VSS 0.00226f
C2023 VDD.n285 VSS 0.00196f
C2024 VDD.n286 VSS 0.00226f
C2025 VDD.n287 VSS 0.00139f
C2026 VDD.n288 VSS 6.75e-19
C2027 VDD.n289 VSS 0.00698f
C2028 VDD.n290 VSS 5.83e-19
C2029 VDD.n291 VSS 0.00207f
C2030 VDD.n292 VSS 0.0017f
C2031 VDD.n293 VSS 8.61e-19
C2032 VDD.n294 VSS 0.00387f
C2033 VDD.n295 VSS 0.0457f
C2034 VDD.n296 VSS 0.0355f
C2035 phi1 VSS 1.58f
C2036 sky130_fd_sc_hd__nand2_1_1/Y VSS 0.159f
C2037 sky130_fd_sc_hd__inv_1_2/Y VSS 1.4f
C2038 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 4.74e-20
C2039 phi2 VSS 1.24f
C2040 sky130_fd_sc_hd__nand2_1_0/Y VSS 0.311f
C2041 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS 8.14e-20
C2042 mimtop1 VSS 47.8f
C2043 mimbot1 VSS 67.1f
C2044 mimtop2 VSS 49.8f
C2045 vcm VSS 75.6f
C2046 VDD VSS 0.161p
C2047 sky130_fd_sc_hd__dlymetal6s6s_1_5/A VSS 0.157f
C2048 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_629_47# VSS 0.124f
C2049 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_523_47# VSS 0.149f
C2050 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_346_47# VSS 0.0937f
C2051 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_240_47# VSS 0.138f
C2052 sky130_fd_sc_hd__dlymetal6s6s_1_4/a_63_47# VSS 0.149f
C2053 sky130_fd_sc_hd__inv_1_1/A VSS 0.466f
C2054 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_629_47# VSS 0.132f
C2055 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_523_47# VSS 0.164f
C2056 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_346_47# VSS 0.11f
C2057 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_240_47# VSS 0.153f
C2058 sky130_fd_sc_hd__dlymetal6s6s_1_5/a_63_47# VSS 0.167f
C2059 sky130_fd_sc_hd__inv_1_0/A VSS 0.464f
C2060 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_629_47# VSS 0.132f
C2061 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_523_47# VSS 0.164f
C2062 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_346_47# VSS 0.11f
C2063 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_240_47# VSS 0.153f
C2064 sky130_fd_sc_hd__dlymetal6s6s_1_3/a_63_47# VSS 0.167f
C2065 sky130_fd_sc_hd__dlymetal6s6s_1_3/A VSS 0.157f
C2066 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_629_47# VSS 0.127f
C2067 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_523_47# VSS 0.159f
C2068 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_346_47# VSS 0.106f
C2069 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_240_47# VSS 0.149f
C2070 sky130_fd_sc_hd__dlymetal6s6s_1_2/a_63_47# VSS 0.163f
C2071 sky130_fd_sc_hd__dlymetal6s6s_1_4/A VSS 0.14f
C2072 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_629_47# VSS 0.113f
C2073 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_523_47# VSS 0.148f
C2074 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_346_47# VSS 0.0949f
C2075 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_240_47# VSS 0.139f
C2076 sky130_fd_sc_hd__dlymetal6s6s_1_1/a_63_47# VSS 0.149f
C2077 sky130_fd_sc_hd__dlymetal6s6s_1_2/A VSS 0.156f
C2078 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_629_47# VSS 0.126f
C2079 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_523_47# VSS 0.159f
C2080 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_346_47# VSS 0.107f
C2081 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_240_47# VSS 0.15f
C2082 sky130_fd_sc_hd__dlymetal6s6s_1_0/a_63_47# VSS 0.211f
C2083 sky130_fd_sc_hd__inv_1_3/Y VSS 0.98f
C2084 sky130_fd_sc_hd__buf_4_3/a_27_47# VSS 0.485f
C2085 sky130_fd_sc_hd__inv_1_3/A VSS 0.373f
C2086 sky130_fd_sc_hd__buf_4_2/a_27_47# VSS 0.444f
C2087 phi1_n VSS 0.843f
C2088 phi2_n VSS 0.581f
C2089 sky130_fd_sc_hd__buf_4_1/a_27_47# VSS 0.483f
C2090 sky130_fd_sc_hd__inv_1_2/A VSS 0.338f
C2091 sky130_fd_sc_hd__buf_4_0/a_27_47# VSS 0.443f
C2092 sky130_fd_sc_hd__inv_1_4/Y VSS 0.182f
C2093 clk VSS 0.68f
.ends

