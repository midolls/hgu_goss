* NGSPICE file created from hgu_delay_no_code_flat.ext - technology: sky130A

.subckt hgu_delay_no_code_flat IN OUT code[3] code[1] code[2] code[0] code_offset
+ VSS VDD
X0 Uc x10.Y.t2 x5[7].floating.t7 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1 Uc code[2].t0 x4[3].floating VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2 x5[7].floating.t6 x10.Y.t3 Uc VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3 Uc code_offset.t0 x7.floating VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4 a_15703_1340# OUT.t2 VDD.t9 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 x3[1].floating code[1].t0 Uc VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X6 a_9893_879# IN.t0 nstack_lab5 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X7 nstack_lab2 IN.t1 a_9893_465# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 pstack_lab4 IN.t2 pstack_lab5 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X9 nstack_lab6 IN.t3 a_9893_1017# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 pstack_lab2 IN.t4 pstack_lab1 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_15703_1340# Uc VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X12 a_15703_1681# Uc OUT.t0 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X13 x4[3].floating code[2].t1 Uc VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X14 VDD.t15 OUT.t3 a_15703_1340# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_9893_465# IN.t5 nstack_lab1 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X16 VDD.t12 code_offset.t1 x6.SW VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X17 VSS.t5 IN.t6 a_9893_327# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 Uc x10.Y.t4 x5[7].floating.t5 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X19 x5[7].floating.t4 x10.Y.t5 Uc VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X20 pstack_lab2 IN.t7 pstack_lab3 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X21 Uc code[1].t1 x3[1].floating VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X22 nstack_lab4 IN.t8 a_9893_741# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 a_9893_327# IN.t9 nstack_lab1 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X24 x10.Y.t0 code[3].t0 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X25 a_15703_1681# Uc VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X26 Uc x6.SW x6.floating VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 VSS.t10 code_offset.t2 x6.SW VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X28 a_9893_1293# IN.t10 nstack_lab7 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x5[7].floating.t3 x10.Y.t6 Uc VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X30 a_15703_1681# OUT.t4 VSS.t12 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_9893_741# IN.t11 nstack_lab3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X32 Uc IN.t12 pstack_lab5 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X33 x5[7].floating.t2 x10.Y.t7 Uc VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X34 Uc x10.Y.t8 x5[7].floating.t1 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X35 Uc code[2].t2 x4[3].floating VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X36 nstack_lab2 IN.t13 a_9893_603# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X37 pstack_lab4 IN.t14 pstack_lab3 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X38 x4[3].floating code[2].t3 Uc VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X39 a_15703_1340# Uc OUT.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X40 Uc IN.t15 a_9893_1293# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 x10.Y.t1 code[3].t1 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X42 a_9893_1155# IN.t16 nstack_lab7 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X43 VDD.t4 IN.t17 pstack_lab1 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X44 Uc x10.Y.t9 x5[7].floating.t0 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X45 VSS.t11 OUT.t5 a_15703_1681# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X46 x2.floating code[0].t0 Uc VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X47 a_9893_603# IN.t18 nstack_lab3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X48 nstack_lab6 IN.t19 a_9893_1155# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 nstack_lab4 IN.t20 a_9893_879# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X50 a_9893_1017# IN.t21 nstack_lab5 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
R0 x10.Y x10.Y.t6 154.847
R1 x10.Y x10.Y.t8 154.8
R2 x10.Y x10.Y.t7 154.8
R3 x10.Y x10.Y.t2 154.8
R4 x10.Y x10.Y.t3 154.8
R5 x10.Y x10.Y.t4 154.8
R6 x10.Y x10.Y.t5 154.8
R7 x10.Y x10.Y.t9 154.8
R8 x10.Y.n0 x10.Y 134.239
R9 x10.Y x10.Y.t1 106.635
R10 x10.Y.n2 x10.Y.t0 24.6567
R11 x10.Y.n5 x10.Y.n4 12.4089
R12 x10.Y.n3 x10.Y.n2 9.12522
R13 x10.Y.n4 x10.Y.n3 7.34048
R14 x10.Y.n5 x10.Y 2.22659
R15 x10.Y.n2 x10.Y.n1 1.93377
R16 x10.Y x10.Y.n5 1.55202
R17 x10.Y.n3 x10.Y.n0 0.69928
R18 x5[7].floating.n95 x5[7].floating.t7 68.0345
R19 x5[7].floating.n24 x5[7].floating.t2 68.0345
R20 x5[7].floating.n42 x5[7].floating.t1 68.0345
R21 x5[7].floating.n54 x5[7].floating.t3 68.0345
R22 x5[7].floating.n154 x5[7].floating.t0 68.0345
R23 x5[7].floating.n142 x5[7].floating.t4 68.0345
R24 x5[7].floating.n12 x5[7].floating.t5 68.0345
R25 x5[7].floating.n109 x5[7].floating.t6 68.0345
R26 x5[7].floating.n73 x5[7].floating.n35 0.660401
R27 x5[7].floating.n91 x5[7].floating.n90 0.660401
R28 x5[7].floating.n130 x5[7].floating.n20 0.660401
R29 x5[7].floating.n139 x5[7].floating.n5 0.660401
R30 x5[7].floating.n121 x5[7].floating.n120 0.660401
R31 x5[7].floating.n60 x5[7].floating.n59 0.320345
R32 x5[7].floating.n160 x5[7].floating.n159 0.308269
R33 x5[7].floating.n161 x5[7].floating.n160 0.173084
R34 x5[7].floating.n61 x5[7].floating.n60 0.162103
R35 x5[7].floating.n160 x5[7].floating 0.100688
R36 x5[7].floating.n60 x5[7].floating 0.0755007
R37 x5[7].floating.n36 x5[7].floating.n35 0.0716912
R38 x5[7].floating.n35 x5[7].floating.n34 0.0716912
R39 x5[7].floating.n6 x5[7].floating.n5 0.0716912
R40 x5[7].floating.n5 x5[7].floating.n4 0.0716912
R41 x5[7].floating.n74 x5[7].floating.n73 0.0716912
R42 x5[7].floating.n122 x5[7].floating.n121 0.0716912
R43 x5[7].floating.n140 x5[7].floating.n139 0.0716912
R44 x5[7].floating.n120 x5[7].floating.n105 0.0716912
R45 x5[7].floating.n120 x5[7].floating.n119 0.0716912
R46 x5[7].floating.n40 x5[7].floating.n39 0.0557941
R47 x5[7].floating.n39 x5[7].floating.n38 0.0557941
R48 x5[7].floating.n38 x5[7].floating.n37 0.0557941
R49 x5[7].floating.n37 x5[7].floating.n36 0.0557941
R50 x5[7].floating.n34 x5[7].floating.n33 0.0557941
R51 x5[7].floating.n33 x5[7].floating.n32 0.0557941
R52 x5[7].floating.n32 x5[7].floating.n31 0.0557941
R53 x5[7].floating.n31 x5[7].floating.n30 0.0557941
R54 x5[7].floating.n10 x5[7].floating.n9 0.0557941
R55 x5[7].floating.n9 x5[7].floating.n8 0.0557941
R56 x5[7].floating.n8 x5[7].floating.n7 0.0557941
R57 x5[7].floating.n7 x5[7].floating.n6 0.0557941
R58 x5[7].floating.n4 x5[7].floating.n3 0.0557941
R59 x5[7].floating.n3 x5[7].floating.n2 0.0557941
R60 x5[7].floating.n2 x5[7].floating.n1 0.0557941
R61 x5[7].floating.n1 x5[7].floating.n0 0.0557941
R62 x5[7].floating.n69 x5[7].floating.n68 0.0557941
R63 x5[7].floating.n70 x5[7].floating.n69 0.0557941
R64 x5[7].floating.n71 x5[7].floating.n70 0.0557941
R65 x5[7].floating.n72 x5[7].floating.n71 0.0557941
R66 x5[7].floating.n76 x5[7].floating.n75 0.0557941
R67 x5[7].floating.n77 x5[7].floating.n76 0.0557941
R68 x5[7].floating.n78 x5[7].floating.n77 0.0557941
R69 x5[7].floating.n86 x5[7].floating.n85 0.0557941
R70 x5[7].floating.n85 x5[7].floating.n84 0.0557941
R71 x5[7].floating.n84 x5[7].floating.n83 0.0557941
R72 x5[7].floating.n83 x5[7].floating.n82 0.0557941
R73 x5[7].floating.n124 x5[7].floating.n123 0.0557941
R74 x5[7].floating.n125 x5[7].floating.n124 0.0557941
R75 x5[7].floating.n126 x5[7].floating.n125 0.0557941
R76 x5[7].floating.n135 x5[7].floating.n134 0.0557941
R77 x5[7].floating.n136 x5[7].floating.n135 0.0557941
R78 x5[7].floating.n137 x5[7].floating.n136 0.0557941
R79 x5[7].floating.n138 x5[7].floating.n137 0.0557941
R80 x5[7].floating.n171 x5[7].floating.n170 0.0557941
R81 x5[7].floating.n170 x5[7].floating.n169 0.0557941
R82 x5[7].floating.n169 x5[7].floating.n168 0.0557941
R83 x5[7].floating.n102 x5[7].floating.n101 0.0557941
R84 x5[7].floating.n103 x5[7].floating.n102 0.0557941
R85 x5[7].floating.n104 x5[7].floating.n103 0.0557941
R86 x5[7].floating.n105 x5[7].floating.n104 0.0557941
R87 x5[7].floating.n119 x5[7].floating.n118 0.0557941
R88 x5[7].floating.n118 x5[7].floating.n117 0.0557941
R89 x5[7].floating.n117 x5[7].floating.n116 0.0557941
R90 x5[7].floating.n116 x5[7].floating.n115 0.0557941
R91 x5[7].floating.n65 x5[7].floating.n64 0.0537206
R92 x5[7].floating.n90 x5[7].floating.n89 0.0537206
R93 x5[7].floating.n131 x5[7].floating.n130 0.0537206
R94 x5[7].floating.n164 x5[7].floating.n163 0.0537206
R95 x5[7].floating.n64 x5[7].floating.n63 0.0530294
R96 x5[7].floating.n90 x5[7].floating.n81 0.0530294
R97 x5[7].floating.n130 x5[7].floating.n129 0.0530294
R98 x5[7].floating.n165 x5[7].floating.n164 0.0530294
R99 x5[7].floating.n92 x5[7].floating.n91 0.0529559
R100 x5[7].floating.n50 x5[7].floating.n49 0.0529559
R101 x5[7].floating.n20 x5[7].floating.n19 0.0529559
R102 x5[7].floating.n151 x5[7].floating.n150 0.0529559
R103 x5[7].floating.n51 x5[7].floating.n50 0.0524559
R104 x5[7].floating.n91 x5[7].floating.n21 0.0524559
R105 x5[7].floating.n106 x5[7].floating.n20 0.0524559
R106 x5[7].floating.n150 x5[7].floating.n149 0.0524559
R107 x5[7].floating.n79 x5[7].floating.n78 0.0523382
R108 x5[7].floating.n127 x5[7].floating.n126 0.0523382
R109 x5[7].floating.n168 x5[7].floating.n167 0.0523382
R110 x5[7].floating.n68 x5[7].floating.n67 0.0516471
R111 x5[7].floating.n87 x5[7].floating.n86 0.0516471
R112 x5[7].floating.n134 x5[7].floating.n133 0.0516471
R113 x5[7].floating.n73 x5[7].floating 0.0495735
R114 x5[7].floating.n121 x5[7].floating 0.0495735
R115 x5[7].floating.n139 x5[7].floating 0.0495735
R116 x5[7].floating.n98 x5[7].floating.n97 0.0408846
R117 x5[7].floating.n45 x5[7].floating.n44 0.0408846
R118 x5[7].floating.n157 x5[7].floating.n156 0.0408846
R119 x5[7].floating.n15 x5[7].floating.n14 0.0408846
R120 x5[7].floating.n75 x5[7].floating 0.0336765
R121 x5[7].floating.n123 x5[7].floating 0.0336765
R122 x5[7].floating x5[7].floating.n171 0.0336765
R123 x5[7].floating.n30 x5[7].floating.n29 0.0271618
R124 x5[7].floating.n115 x5[7].floating.n114 0.0271618
R125 x5[7].floating.n101 x5[7].floating.n100 0.0266618
R126 x5[7].floating.n41 x5[7].floating.n40 0.0266618
R127 x5[7].floating.n11 x5[7].floating.n10 0.0266618
R128 x5[7].floating x5[7].floating.n72 0.0226176
R129 x5[7].floating x5[7].floating.n74 0.0226176
R130 x5[7].floating.n82 x5[7].floating 0.0226176
R131 x5[7].floating x5[7].floating.n122 0.0226176
R132 x5[7].floating x5[7].floating.n138 0.0226176
R133 x5[7].floating x5[7].floating.n140 0.0226176
R134 x5[7].floating.n63 x5[7].floating.n62 0.0191618
R135 x5[7].floating.n81 x5[7].floating.n80 0.0191618
R136 x5[7].floating.n129 x5[7].floating.n128 0.0191618
R137 x5[7].floating.n166 x5[7].floating.n165 0.0191618
R138 x5[7].floating.n66 x5[7].floating.n65 0.0184706
R139 x5[7].floating.n89 x5[7].floating.n88 0.0184706
R140 x5[7].floating.n132 x5[7].floating.n131 0.0184706
R141 x5[7].floating.n163 x5[7].floating.n162 0.0184706
R142 x5[7].floating.n100 x5[7].floating.n99 0.014
R143 x5[7].floating.n52 x5[7].floating.n51 0.014
R144 x5[7].floating.n46 x5[7].floating.n41 0.014
R145 x5[7].floating.n22 x5[7].floating.n21 0.014
R146 x5[7].floating.n16 x5[7].floating.n11 0.014
R147 x5[7].floating.n149 x5[7].floating.n148 0.014
R148 x5[7].floating.n159 x5[7].floating.n158 0.014
R149 x5[7].floating.n107 x5[7].floating.n106 0.014
R150 x5[7].floating.n93 x5[7].floating.n92 0.0135
R151 x5[7].floating.n59 x5[7].floating.n58 0.0135
R152 x5[7].floating.n49 x5[7].floating.n48 0.0135
R153 x5[7].floating.n29 x5[7].floating.n28 0.0135
R154 x5[7].floating.n19 x5[7].floating.n18 0.0135
R155 x5[7].floating.n146 x5[7].floating.n141 0.0135
R156 x5[7].floating.n152 x5[7].floating.n151 0.0135
R157 x5[7].floating.n114 x5[7].floating.n113 0.0135
R158 x5[7].floating.n27 x5[7].floating.n26 0.0120385
R159 x5[7].floating.n57 x5[7].floating.n56 0.0120385
R160 x5[7].floating.n145 x5[7].floating.n144 0.0120385
R161 x5[7].floating.n112 x5[7].floating.n111 0.0120385
R162 x5[7].floating.n67 x5[7].floating.n66 0.00464706
R163 x5[7].floating.n88 x5[7].floating.n87 0.00464706
R164 x5[7].floating.n133 x5[7].floating.n132 0.00464706
R165 x5[7].floating.n162 x5[7].floating.n161 0.00464706
R166 x5[7].floating.n62 x5[7].floating.n61 0.00395588
R167 x5[7].floating.n80 x5[7].floating.n79 0.00395588
R168 x5[7].floating.n128 x5[7].floating.n127 0.00395588
R169 x5[7].floating.n167 x5[7].floating.n166 0.00395588
R170 x5[7].floating.n110 x5[7].floating.n109 0.00359614
R171 x5[7].floating.n25 x5[7].floating.n24 0.00359614
R172 x5[7].floating.n55 x5[7].floating.n54 0.00359614
R173 x5[7].floating.n143 x5[7].floating.n142 0.00359614
R174 x5[7].floating.n94 x5[7].floating.n93 0.0035
R175 x5[7].floating.n58 x5[7].floating.n53 0.0035
R176 x5[7].floating.n48 x5[7].floating.n47 0.0035
R177 x5[7].floating.n28 x5[7].floating.n23 0.0035
R178 x5[7].floating.n18 x5[7].floating.n17 0.0035
R179 x5[7].floating.n147 x5[7].floating.n146 0.0035
R180 x5[7].floating.n153 x5[7].floating.n152 0.0035
R181 x5[7].floating.n113 x5[7].floating.n108 0.0035
R182 x5[7].floating.n99 x5[7].floating.n94 0.003
R183 x5[7].floating.n53 x5[7].floating.n52 0.003
R184 x5[7].floating.n47 x5[7].floating.n46 0.003
R185 x5[7].floating.n23 x5[7].floating.n22 0.003
R186 x5[7].floating.n17 x5[7].floating.n16 0.003
R187 x5[7].floating.n148 x5[7].floating.n147 0.003
R188 x5[7].floating.n158 x5[7].floating.n153 0.003
R189 x5[7].floating.n108 x5[7].floating.n107 0.003
R190 x5[7].floating.n155 x5[7].floating.n154 0.00277942
R191 x5[7].floating.n96 x5[7].floating.n95 0.0023396
R192 x5[7].floating.n43 x5[7].floating.n42 0.0023396
R193 x5[7].floating.n13 x5[7].floating.n12 0.0023396
R194 x5[7].floating.n157 x5[7].floating.n155 0.00233747
R195 x5[7].floating.n98 x5[7].floating.n96 0.00200689
R196 x5[7].floating.n45 x5[7].floating.n43 0.00200689
R197 x5[7].floating.n15 x5[7].floating.n13 0.00200689
R198 x5[7].floating.n27 x5[7].floating.n25 0.0010233
R199 x5[7].floating.n57 x5[7].floating.n55 0.0010233
R200 x5[7].floating.n145 x5[7].floating.n143 0.0010233
R201 x5[7].floating.n112 x5[7].floating.n110 0.0010233
R202 x5[7].floating.n99 x5[7].floating.n98 0.00053972
R203 x5[7].floating.n58 x5[7].floating.n57 0.00053972
R204 x5[7].floating.n46 x5[7].floating.n45 0.00053972
R205 x5[7].floating.n28 x5[7].floating.n27 0.00053972
R206 x5[7].floating.n16 x5[7].floating.n15 0.00053972
R207 x5[7].floating.n146 x5[7].floating.n145 0.00053972
R208 x5[7].floating.n158 x5[7].floating.n157 0.00053972
R209 x5[7].floating.n113 x5[7].floating.n112 0.00053972
R210 VDD.n1742 VDD.n4 426
R211 VDD.n1766 VDD.n2 351
R212 VDD.t11 VDD.n3 258.856
R213 VDD.n717 VDD.n129 198.118
R214 VDD.n540 VDD.n140 198.118
R215 VDD.n363 VDD.n151 198.118
R216 VDD.n1015 VDD.n1014 198.118
R217 VDD.n362 VDD.n152 198.118
R218 VDD.n539 VDD.n141 198.118
R219 VDD.n716 VDD.n130 198.118
R220 VDD.t5 VDD.n1764 188.965
R221 VDD.n902 VDD.n901 185
R222 VDD.n1071 VDD.n889 185
R223 VDD.n932 VDD.n930 185
R224 VDD.n1050 VDD.n928 185
R225 VDD.n1020 VDD.n1018 185
R226 VDD.n1070 VDD.n1069 185
R227 VDD.n1070 VDD.n118 185
R228 VDD.n941 VDD.n940 185
R229 VDD.n941 VDD.n118 185
R230 VDD.n1049 VDD.n1048 185
R231 VDD.n1049 VDD.n118 185
R232 VDD.n1029 VDD.n1028 185
R233 VDD.n1016 VDD.n967 185
R234 VDD.n894 VDD.n893 185
R235 VDD.n189 VDD.n82 185
R236 VDD.n161 VDD.n159 185
R237 VDD.n237 VDD.n236 185
R238 VDD.n1682 VDD.n246 185
R239 VDD.n264 VDD.n247 185
R240 VDD.n1657 VDD.n1656 185
R241 VDD.n1659 VDD.n1658 185
R242 VDD.n1629 VDD.n1628 185
R243 VDD.n1638 VDD.n1637 185
R244 VDD.n1623 VDD.n1622 185
R245 VDD.n1625 VDD.n1624 185
R246 VDD.n1595 VDD.n1594 185
R247 VDD.n1604 VDD.n1603 185
R248 VDD.n1589 VDD.n1588 185
R249 VDD.n1591 VDD.n1590 185
R250 VDD.n361 VDD.n360 185
R251 VDD.n380 VDD.n379 185
R252 VDD.n396 VDD.n395 185
R253 VDD.n412 VDD.n411 185
R254 VDD.n1519 VDD.n427 185
R255 VDD.n441 VDD.n428 185
R256 VDD.n1494 VDD.n1493 185
R257 VDD.n1496 VDD.n1495 185
R258 VDD.n1466 VDD.n1465 185
R259 VDD.n1475 VDD.n1474 185
R260 VDD.n1460 VDD.n1459 185
R261 VDD.n1462 VDD.n1461 185
R262 VDD.n1432 VDD.n1431 185
R263 VDD.n1441 VDD.n1440 185
R264 VDD.n1426 VDD.n1425 185
R265 VDD.n1428 VDD.n1427 185
R266 VDD.n538 VDD.n537 185
R267 VDD.n557 VDD.n556 185
R268 VDD.n573 VDD.n572 185
R269 VDD.n589 VDD.n588 185
R270 VDD.n1356 VDD.n604 185
R271 VDD.n618 VDD.n605 185
R272 VDD.n1331 VDD.n1330 185
R273 VDD.n1333 VDD.n1332 185
R274 VDD.n1303 VDD.n1302 185
R275 VDD.n1312 VDD.n1311 185
R276 VDD.n1297 VDD.n1296 185
R277 VDD.n1299 VDD.n1298 185
R278 VDD.n1269 VDD.n1268 185
R279 VDD.n1278 VDD.n1277 185
R280 VDD.n1263 VDD.n1262 185
R281 VDD.n1265 VDD.n1264 185
R282 VDD.n715 VDD.n714 185
R283 VDD.n734 VDD.n733 185
R284 VDD.n750 VDD.n749 185
R285 VDD.n766 VDD.n765 185
R286 VDD.n1193 VDD.n781 185
R287 VDD.n795 VDD.n782 185
R288 VDD.n1168 VDD.n1167 185
R289 VDD.n1170 VDD.n1169 185
R290 VDD.n1140 VDD.n1139 185
R291 VDD.n1149 VDD.n1148 185
R292 VDD.n1134 VDD.n1133 185
R293 VDD.n1136 VDD.n1135 185
R294 VDD.n1106 VDD.n1105 185
R295 VDD.n1115 VDD.n1114 185
R296 VDD.n1100 VDD.n1099 185
R297 VDD.n1102 VDD.n1101 185
R298 VDD.n768 VDD.n767 185
R299 VDD.n752 VDD.n751 185
R300 VDD.n736 VDD.n735 185
R301 VDD.n721 VDD.n720 185
R302 VDD.n797 VDD.n796 185
R303 VDD.n719 VDD.n718 185
R304 VDD.n591 VDD.n590 185
R305 VDD.n575 VDD.n574 185
R306 VDD.n559 VDD.n558 185
R307 VDD.n544 VDD.n543 185
R308 VDD.n620 VDD.n619 185
R309 VDD.n542 VDD.n541 185
R310 VDD.n414 VDD.n413 185
R311 VDD.n398 VDD.n397 185
R312 VDD.n382 VDD.n381 185
R313 VDD.n367 VDD.n366 185
R314 VDD.n443 VDD.n442 185
R315 VDD.n365 VDD.n364 185
R316 VDD.n245 VDD.n244 185
R317 VDD.n235 VDD.n160 185
R318 VDD.n208 VDD.n207 185
R319 VDD.n266 VDD.n265 185
R320 VDD.n179 VDD.n178 185
R321 VDD.n1760 VDD.n2 185
R322 VDD.n1764 VDD.n2 185
R323 VDD.n1765 VDD 160.49
R324 VDD.n1768 VDD.t6 152.88
R325 VDD.n28 VDD.t12 152.879
R326 VDD.n1734 VDD.n29 121.447
R327 VDD.n1734 VDD.n34 121.447
R328 VDD.n1738 VDD.n29 118.555
R329 VDD.n1011 VDD.n989 117.007
R330 VDD.n1765 VDD.t5 113.897
R331 VDD.n1150 VDD.n1149 111.177
R332 VDD.n1116 VDD.n1115 111.177
R333 VDD.n720 VDD.n128 111.177
R334 VDD.n735 VDD.n110 111.177
R335 VDD.n751 VDD.n126 111.177
R336 VDD.n767 VDD.n112 111.177
R337 VDD.n1313 VDD.n1312 111.177
R338 VDD.n1279 VDD.n1278 111.177
R339 VDD.n543 VDD.n139 111.177
R340 VDD.n558 VDD.n101 111.177
R341 VDD.n574 VDD.n137 111.177
R342 VDD.n590 VDD.n103 111.177
R343 VDD.n1476 VDD.n1475 111.177
R344 VDD.n1442 VDD.n1441 111.177
R345 VDD.n366 VDD.n150 111.177
R346 VDD.n381 VDD.n92 111.177
R347 VDD.n397 VDD.n148 111.177
R348 VDD.n413 VDD.n94 111.177
R349 VDD.n1639 VDD.n1638 111.177
R350 VDD.n1605 VDD.n1604 111.177
R351 VDD.n207 VDD.n206 111.177
R352 VDD.n1705 VDD.n160 111.177
R353 VDD.n244 VDD.n85 111.177
R354 VDD.n1073 VDD.n902 111.177
R355 VDD.n1070 VDD.n903 111.177
R356 VDD.n1052 VDD.n941 111.177
R357 VDD.n1049 VDD.n942 111.177
R358 VDD.n1741 VDD.t11 108.719
R359 VDD.n1006 VDD.n989 106.648
R360 VDD.n1003 VDD.n34 101.276
R361 VDD.n1006 VDD.n1003 101.206
R362 VDD.n1762 VDD.n1761 92.5005
R363 VDD.n1763 VDD.n1762 92.5005
R364 VDD.n1767 VDD.n1766 92.5005
R365 VDD.n1766 VDD.n1765 92.5005
R366 VDD.n1743 VDD.n1742 92.5005
R367 VDD.n1742 VDD.n1741 92.5005
R368 VDD.n890 VDD.n118 85.9427
R369 VDD.n1015 VDD.n118 85.9427
R370 VDD.n1706 VDD.n84 85.9427
R371 VDD.n1706 VDD.n158 85.9427
R372 VDD.n1706 VDD.n86 85.9427
R373 VDD.n1706 VDD.n156 85.9427
R374 VDD.n1706 VDD.n154 85.9427
R375 VDD.n1706 VDD.n152 85.9427
R376 VDD.n1706 VDD.n151 85.9427
R377 VDD.n1706 VDD.n149 85.9427
R378 VDD.n1706 VDD.n93 85.9427
R379 VDD.n1706 VDD.n147 85.9427
R380 VDD.n1706 VDD.n95 85.9427
R381 VDD.n1706 VDD.n145 85.9427
R382 VDD.n1706 VDD.n143 85.9427
R383 VDD.n1706 VDD.n141 85.9427
R384 VDD.n1706 VDD.n140 85.9427
R385 VDD.n1706 VDD.n138 85.9427
R386 VDD.n1706 VDD.n102 85.9427
R387 VDD.n1706 VDD.n136 85.9427
R388 VDD.n1706 VDD.n104 85.9427
R389 VDD.n1706 VDD.n134 85.9427
R390 VDD.n1706 VDD.n132 85.9427
R391 VDD.n1706 VDD.n130 85.9427
R392 VDD.n1706 VDD.n129 85.9427
R393 VDD.n1706 VDD.n127 85.9427
R394 VDD.n1706 VDD.n111 85.9427
R395 VDD.n1706 VDD.n125 85.9427
R396 VDD.n1706 VDD.n113 85.9427
R397 VDD.n1706 VDD.n123 85.9427
R398 VDD.n1706 VDD.n121 85.9427
R399 VDD.n1741 VDD 77.6572
R400 VDD.n52 VDD.t1 70.3649
R401 VDD.n987 VDD.t4 68.0287
R402 VDD.n1707 VDD.n82 67.5405
R403 VDD.n1100 VDD.n119 67.5405
R404 VDD.n795 VDD.n114 67.3307
R405 VDD.n618 VDD.n105 67.3307
R406 VDD.n441 VDD.n96 67.3307
R407 VDD.n264 VDD.n87 67.3307
R408 VDD.n1030 VDD.n1029 67.3307
R409 VDD.n1657 VDD.n89 67.3307
R410 VDD.n1623 VDD.n90 67.3307
R411 VDD.n1589 VDD.n91 67.3307
R412 VDD.n1494 VDD.n98 67.3307
R413 VDD.n1460 VDD.n99 67.3307
R414 VDD.n1426 VDD.n100 67.3307
R415 VDD.n1331 VDD.n107 67.3307
R416 VDD.n1297 VDD.n108 67.3307
R417 VDD.n1263 VDD.n109 67.3307
R418 VDD.n1168 VDD.n116 67.3307
R419 VDD.n1134 VDD.n117 67.3307
R420 VDD VDD.n1740 49.0494
R421 VDD.n45 VDD.t9 47.1434
R422 VDD.n45 VDD.t15 47.1434
R423 VDD.n31 VDD.n30 41.3127
R424 VDD.n1762 VDD.n2 39.0005
R425 VDD.n32 VDD.t0 35.8207
R426 VDD.n363 VDD.n362 33.746
R427 VDD.n540 VDD.n539 33.746
R428 VDD.n717 VDD.n716 33.746
R429 VDD.n1764 VDD.n1763 33.6517
R430 VDD.n1668 VDD.n267 32.9702
R431 VDD.n1505 VDD.n444 32.9702
R432 VDD.n1342 VDD.n621 32.9702
R433 VDD.n1179 VDD.n798 32.9702
R434 VDD.n1169 VDD.n1168 28.2358
R435 VDD.n1135 VDD.n1134 28.2358
R436 VDD.n1101 VDD.n1100 28.2358
R437 VDD.n796 VDD.n795 28.2358
R438 VDD.n1332 VDD.n1331 28.2358
R439 VDD.n1298 VDD.n1297 28.2358
R440 VDD.n1264 VDD.n1263 28.2358
R441 VDD.n619 VDD.n618 28.2358
R442 VDD.n1495 VDD.n1494 28.2358
R443 VDD.n1461 VDD.n1460 28.2358
R444 VDD.n1427 VDD.n1426 28.2358
R445 VDD.n442 VDD.n441 28.2358
R446 VDD.n1658 VDD.n1657 28.2358
R447 VDD.n1624 VDD.n1623 28.2358
R448 VDD.n1590 VDD.n1589 28.2358
R449 VDD.n178 VDD.n82 28.2358
R450 VDD.n265 VDD.n264 28.2358
R451 VDD.n1071 VDD.n1070 28.2358
R452 VDD.n941 VDD.n930 28.2358
R453 VDD.n1050 VDD.n1049 28.2358
R454 VDD.n1029 VDD.n1018 28.2358
R455 VDD.t0 VDD.t2 21.1252
R456 VDD.n1013 VDD.n1012 21.0038
R457 VDD.n993 VDD.n992 20.7428
R458 VDD.n1009 VDD.n996 20.7428
R459 VDD.n1000 VDD.n999 20.7428
R460 VDD.n61 VDD.n35 20.7428
R461 VDD.n1731 VDD.n1730 20.7428
R462 VDD.n1737 VDD.n32 18.2316
R463 VDD.t13 VDD 16.5329
R464 VDD.n1746 VDD.n1745 15.7543
R465 VDD.n1760 VDD.n1 13.7851
R466 VDD.n1013 VDD.n987 13.3673
R467 VDD.n1737 VDD.n1736 13.1567
R468 VDD.n28 VDD 13.1403
R469 VDD.n1769 VDD.n1768 13.1182
R470 VDD.n1139 VDD.n123 13.1177
R471 VDD.n1105 VDD.n121 13.1177
R472 VDD.n733 VDD.n127 13.1177
R473 VDD.n749 VDD.n111 13.1177
R474 VDD.n765 VDD.n125 13.1177
R475 VDD.n1193 VDD.n113 13.1177
R476 VDD.n1302 VDD.n134 13.1177
R477 VDD.n1268 VDD.n132 13.1177
R478 VDD.n714 VDD.n130 13.1177
R479 VDD.n556 VDD.n138 13.1177
R480 VDD.n572 VDD.n102 13.1177
R481 VDD.n588 VDD.n136 13.1177
R482 VDD.n1356 VDD.n104 13.1177
R483 VDD.n1465 VDD.n145 13.1177
R484 VDD.n1431 VDD.n143 13.1177
R485 VDD.n537 VDD.n141 13.1177
R486 VDD.n379 VDD.n149 13.1177
R487 VDD.n395 VDD.n93 13.1177
R488 VDD.n411 VDD.n147 13.1177
R489 VDD.n1519 VDD.n95 13.1177
R490 VDD.n1628 VDD.n156 13.1177
R491 VDD.n1594 VDD.n154 13.1177
R492 VDD.n360 VDD.n152 13.1177
R493 VDD.n159 VDD.n84 13.1177
R494 VDD.n236 VDD.n158 13.1177
R495 VDD.n1682 VDD.n86 13.1177
R496 VDD.n902 VDD.n890 13.1177
R497 VDD.n1016 VDD.n1015 13.1177
R498 VDD.n893 VDD.n890 13.1177
R499 VDD.n1638 VDD.n156 13.1177
R500 VDD.n1604 VDD.n154 13.1177
R501 VDD.n1475 VDD.n145 13.1177
R502 VDD.n1441 VDD.n143 13.1177
R503 VDD.n1312 VDD.n134 13.1177
R504 VDD.n1278 VDD.n132 13.1177
R505 VDD.n1149 VDD.n123 13.1177
R506 VDD.n1115 VDD.n121 13.1177
R507 VDD.n767 VDD.n113 13.1177
R508 VDD.n751 VDD.n125 13.1177
R509 VDD.n735 VDD.n111 13.1177
R510 VDD.n720 VDD.n127 13.1177
R511 VDD.n718 VDD.n129 13.1177
R512 VDD.n590 VDD.n104 13.1177
R513 VDD.n574 VDD.n136 13.1177
R514 VDD.n558 VDD.n102 13.1177
R515 VDD.n543 VDD.n138 13.1177
R516 VDD.n541 VDD.n140 13.1177
R517 VDD.n413 VDD.n95 13.1177
R518 VDD.n397 VDD.n147 13.1177
R519 VDD.n381 VDD.n93 13.1177
R520 VDD.n366 VDD.n149 13.1177
R521 VDD.n364 VDD.n151 13.1177
R522 VDD.n244 VDD.n86 13.1177
R523 VDD.n160 VDD.n158 13.1177
R524 VDD.n207 VDD.n84 13.1177
R525 VDD.n1736 VDD.n1735 12.9547
R526 VDD.n1735 VDD.n33 12.9547
R527 VDD.n1012 VDD.n988 12.4812
R528 VDD.n1762 VDD.n4 12.0005
R529 VDD.n32 VDD.t10 11.7875
R530 VDD.n862 VDD.n119 11.5452
R531 VDD.n1708 VDD.n1707 11.5452
R532 VDD.n1005 VDD.n988 11.3763
R533 VDD.n1004 VDD.n33 10.8033
R534 VDD.n1005 VDD.n1004 10.7957
R535 VDD.n1009 VDD.n1008 10.4098
R536 VDD.n1763 VDD.n3 10.3547
R537 VDD.n1171 VDD.n124 9.38471
R538 VDD.n1181 VDD.n115 9.38471
R539 VDD.n1334 VDD.n135 9.38471
R540 VDD.n1344 VDD.n106 9.38471
R541 VDD.n1497 VDD.n146 9.38471
R542 VDD.n1507 VDD.n97 9.38471
R543 VDD.n1660 VDD.n157 9.38471
R544 VDD.n1670 VDD.n88 9.38471
R545 VDD.n1668 VDD.n1667 9.3005
R546 VDD.n1587 VDD.n1586 9.3005
R547 VDD.n1621 VDD.n1620 9.3005
R548 VDD.n1655 VDD.n1654 9.3005
R549 VDD.n270 VDD.n267 9.3005
R550 VDD.n1636 VDD.n1635 9.3005
R551 VDD.n1602 VDD.n1601 9.3005
R552 VDD.n1505 VDD.n1504 9.3005
R553 VDD.n1424 VDD.n1423 9.3005
R554 VDD.n1458 VDD.n1457 9.3005
R555 VDD.n1492 VDD.n1491 9.3005
R556 VDD.n447 VDD.n444 9.3005
R557 VDD.n1473 VDD.n1472 9.3005
R558 VDD.n1439 VDD.n1438 9.3005
R559 VDD.n1342 VDD.n1341 9.3005
R560 VDD.n1261 VDD.n1260 9.3005
R561 VDD.n1295 VDD.n1294 9.3005
R562 VDD.n1329 VDD.n1328 9.3005
R563 VDD.n624 VDD.n621 9.3005
R564 VDD.n1310 VDD.n1309 9.3005
R565 VDD.n1276 VDD.n1275 9.3005
R566 VDD.n1179 VDD.n1178 9.3005
R567 VDD.n1098 VDD.n1097 9.3005
R568 VDD.n1132 VDD.n1131 9.3005
R569 VDD.n1166 VDD.n1165 9.3005
R570 VDD.n801 VDD.n798 9.3005
R571 VDD.n1147 VDD.n1146 9.3005
R572 VDD.n1113 VDD.n1112 9.3005
R573 VDD.n1191 VDD.n1190 9.3005
R574 VDD.n1205 VDD.n1204 9.3005
R575 VDD.n1217 VDD.n1216 9.3005
R576 VDD.n1229 VDD.n1228 9.3005
R577 VDD.n1241 VDD.n1240 9.3005
R578 VDD.n1354 VDD.n1353 9.3005
R579 VDD.n1368 VDD.n1367 9.3005
R580 VDD.n1380 VDD.n1379 9.3005
R581 VDD.n1392 VDD.n1391 9.3005
R582 VDD.n1404 VDD.n1403 9.3005
R583 VDD.n1517 VDD.n1516 9.3005
R584 VDD.n1531 VDD.n1530 9.3005
R585 VDD.n1543 VDD.n1542 9.3005
R586 VDD.n1555 VDD.n1554 9.3005
R587 VDD.n1567 VDD.n1566 9.3005
R588 VDD.n1680 VDD.n1679 9.3005
R589 VDD.n243 VDD.n242 9.3005
R590 VDD.n234 VDD.n165 9.3005
R591 VDD.n191 VDD.n190 9.3005
R592 VDD.n210 VDD.n209 9.3005
R593 VDD.n900 VDD.n899 9.3005
R594 VDD.n1068 VDD.n1067 9.3005
R595 VDD.n939 VDD.n938 9.3005
R596 VDD.n1047 VDD.n1046 9.3005
R597 VDD.n1027 VDD.n1026 9.3005
R598 VDD.n1075 VDD.n1074 9.3005
R599 VDD.n1074 VDD.n1073 9.3005
R600 VDD.n931 VDD.n906 9.3005
R601 VDD.n931 VDD.n903 9.3005
R602 VDD.n1054 VDD.n1053 9.3005
R603 VDD.n1053 VDD.n1052 9.3005
R604 VDD.n1019 VDD.n945 9.3005
R605 VDD.n1019 VDD.n942 9.3005
R606 VDD.n1033 VDD.n1032 9.3005
R607 VDD.n1032 VDD.n1031 9.3005
R608 VDD.n892 VDD.n891 9.3005
R609 VDD.n892 VDD.n118 9.3005
R610 VDD.n358 VDD.n331 9.3005
R611 VDD.n359 VDD.n358 9.3005
R612 VDD.n1592 VDD.n307 9.3005
R613 VDD.n1593 VDD.n1592 9.3005
R614 VDD.n1626 VDD.n274 9.3005
R615 VDD.n1627 VDD.n1626 9.3005
R616 VDD.n1660 VDD.n271 9.3005
R617 VDD.n1641 VDD.n1640 9.3005
R618 VDD.n1640 VDD.n1639 9.3005
R619 VDD.n1607 VDD.n1606 9.3005
R620 VDD.n1606 VDD.n1605 9.3005
R621 VDD.n535 VDD.n508 9.3005
R622 VDD.n536 VDD.n535 9.3005
R623 VDD.n1429 VDD.n484 9.3005
R624 VDD.n1430 VDD.n1429 9.3005
R625 VDD.n1463 VDD.n451 9.3005
R626 VDD.n1464 VDD.n1463 9.3005
R627 VDD.n1497 VDD.n448 9.3005
R628 VDD.n1478 VDD.n1477 9.3005
R629 VDD.n1477 VDD.n1476 9.3005
R630 VDD.n1444 VDD.n1443 9.3005
R631 VDD.n1443 VDD.n1442 9.3005
R632 VDD.n712 VDD.n685 9.3005
R633 VDD.n713 VDD.n712 9.3005
R634 VDD.n1266 VDD.n661 9.3005
R635 VDD.n1267 VDD.n1266 9.3005
R636 VDD.n1300 VDD.n628 9.3005
R637 VDD.n1301 VDD.n1300 9.3005
R638 VDD.n1334 VDD.n625 9.3005
R639 VDD.n1315 VDD.n1314 9.3005
R640 VDD.n1314 VDD.n1313 9.3005
R641 VDD.n1281 VDD.n1280 9.3005
R642 VDD.n1280 VDD.n1279 9.3005
R643 VDD.n1103 VDD.n838 9.3005
R644 VDD.n1104 VDD.n1103 9.3005
R645 VDD.n1137 VDD.n805 9.3005
R646 VDD.n1138 VDD.n1137 9.3005
R647 VDD.n1171 VDD.n802 9.3005
R648 VDD.n1152 VDD.n1151 9.3005
R649 VDD.n1151 VDD.n1150 9.3005
R650 VDD.n1118 VDD.n1117 9.3005
R651 VDD.n1117 VDD.n1116 9.3005
R652 VDD.n863 VDD.n862 9.3005
R653 VDD.n1196 VDD.n1195 9.3005
R654 VDD.n1195 VDD.n1194 9.3005
R655 VDD.n1208 VDD.n1207 9.3005
R656 VDD.n1207 VDD.n112 9.3005
R657 VDD.n1706 VDD.n112 9.3005
R658 VDD.n1220 VDD.n1219 9.3005
R659 VDD.n1219 VDD.n126 9.3005
R660 VDD.n1706 VDD.n126 9.3005
R661 VDD.n1232 VDD.n1231 9.3005
R662 VDD.n1231 VDD.n110 9.3005
R663 VDD.n1706 VDD.n110 9.3005
R664 VDD.n1182 VDD.n1181 9.3005
R665 VDD.n1244 VDD.n1243 9.3005
R666 VDD.n1243 VDD.n128 9.3005
R667 VDD.n1706 VDD.n128 9.3005
R668 VDD.n1359 VDD.n1358 9.3005
R669 VDD.n1358 VDD.n1357 9.3005
R670 VDD.n1371 VDD.n1370 9.3005
R671 VDD.n1370 VDD.n103 9.3005
R672 VDD.n1706 VDD.n103 9.3005
R673 VDD.n1383 VDD.n1382 9.3005
R674 VDD.n1382 VDD.n137 9.3005
R675 VDD.n1706 VDD.n137 9.3005
R676 VDD.n1395 VDD.n1394 9.3005
R677 VDD.n1394 VDD.n101 9.3005
R678 VDD.n1706 VDD.n101 9.3005
R679 VDD.n1345 VDD.n1344 9.3005
R680 VDD.n1407 VDD.n1406 9.3005
R681 VDD.n1406 VDD.n139 9.3005
R682 VDD.n1706 VDD.n139 9.3005
R683 VDD.n1522 VDD.n1521 9.3005
R684 VDD.n1521 VDD.n1520 9.3005
R685 VDD.n1534 VDD.n1533 9.3005
R686 VDD.n1533 VDD.n94 9.3005
R687 VDD.n1706 VDD.n94 9.3005
R688 VDD.n1546 VDD.n1545 9.3005
R689 VDD.n1545 VDD.n148 9.3005
R690 VDD.n1706 VDD.n148 9.3005
R691 VDD.n1558 VDD.n1557 9.3005
R692 VDD.n1557 VDD.n92 9.3005
R693 VDD.n1706 VDD.n92 9.3005
R694 VDD.n1508 VDD.n1507 9.3005
R695 VDD.n1570 VDD.n1569 9.3005
R696 VDD.n1569 VDD.n150 9.3005
R697 VDD.n1706 VDD.n150 9.3005
R698 VDD.n1685 VDD.n1684 9.3005
R699 VDD.n1684 VDD.n1683 9.3005
R700 VDD.n238 VDD.n167 9.3005
R701 VDD.n238 VDD.n85 9.3005
R702 VDD.n1706 VDD.n85 9.3005
R703 VDD.n1704 VDD.n1703 9.3005
R704 VDD.n1705 VDD.n1704 9.3005
R705 VDD.n1706 VDD.n1705 9.3005
R706 VDD.n1671 VDD.n1670 9.3005
R707 VDD.n1709 VDD.n1708 9.3005
R708 VDD.n205 VDD.n204 9.3005
R709 VDD.n206 VDD.n205 9.3005
R710 VDD.n1745 VDD.n1744 9.3005
R711 VDD.n1759 VDD.n1758 9.3005
R712 VDD.n1759 VDD.n4 9.3005
R713 VDD.n4 VDD.n3 9.3005
R714 VDD.n1767 VDD.n1 9.25588
R715 VDD.n1002 VDD.n1000 9.18516
R716 VDD.n190 VDD.n189 8.92171
R717 VDD.n209 VDD.n208 8.92171
R718 VDD.n235 VDD.n234 8.92171
R719 VDD.n245 VDD.n243 8.92171
R720 VDD.n1680 VDD.n247 8.92171
R721 VDD.n1656 VDD.n1655 8.92171
R722 VDD.n1637 VDD.n1636 8.92171
R723 VDD.n1622 VDD.n1621 8.92171
R724 VDD.n1603 VDD.n1602 8.92171
R725 VDD.n1588 VDD.n1587 8.92171
R726 VDD.n1567 VDD.n367 8.92171
R727 VDD.n1555 VDD.n382 8.92171
R728 VDD.n1543 VDD.n398 8.92171
R729 VDD.n1531 VDD.n414 8.92171
R730 VDD.n1517 VDD.n428 8.92171
R731 VDD.n1493 VDD.n1492 8.92171
R732 VDD.n1474 VDD.n1473 8.92171
R733 VDD.n1459 VDD.n1458 8.92171
R734 VDD.n1440 VDD.n1439 8.92171
R735 VDD.n1425 VDD.n1424 8.92171
R736 VDD.n1404 VDD.n544 8.92171
R737 VDD.n1392 VDD.n559 8.92171
R738 VDD.n1380 VDD.n575 8.92171
R739 VDD.n1368 VDD.n591 8.92171
R740 VDD.n1354 VDD.n605 8.92171
R741 VDD.n1330 VDD.n1329 8.92171
R742 VDD.n1311 VDD.n1310 8.92171
R743 VDD.n1296 VDD.n1295 8.92171
R744 VDD.n1277 VDD.n1276 8.92171
R745 VDD.n1262 VDD.n1261 8.92171
R746 VDD.n1241 VDD.n721 8.92171
R747 VDD.n1229 VDD.n736 8.92171
R748 VDD.n1217 VDD.n752 8.92171
R749 VDD.n1205 VDD.n768 8.92171
R750 VDD.n1191 VDD.n782 8.92171
R751 VDD.n1167 VDD.n1166 8.92171
R752 VDD.n1148 VDD.n1147 8.92171
R753 VDD.n1133 VDD.n1132 8.92171
R754 VDD.n1114 VDD.n1113 8.92171
R755 VDD.n1099 VDD.n1098 8.92171
R756 VDD.n901 VDD.n900 8.92171
R757 VDD.n1069 VDD.n1068 8.92171
R758 VDD.n940 VDD.n939 8.92171
R759 VDD.n1048 VDD.n1047 8.92171
R760 VDD.n1028 VDD.n1027 8.92171
R761 VDD.n1746 VDD.n1743 8.86204
R762 VDD.n1072 VDD.n118 8.77616
R763 VDD.n929 VDD.n118 8.77616
R764 VDD.n1051 VDD.n118 8.77616
R765 VDD.n1017 VDD.n118 8.77616
R766 VDD.n1706 VDD.n157 8.77616
R767 VDD.n1706 VDD.n155 8.77616
R768 VDD.n1706 VDD.n153 8.77616
R769 VDD.n1706 VDD.n146 8.77616
R770 VDD.n1706 VDD.n144 8.77616
R771 VDD.n1706 VDD.n142 8.77616
R772 VDD.n1706 VDD.n135 8.77616
R773 VDD.n1706 VDD.n133 8.77616
R774 VDD.n1706 VDD.n131 8.77616
R775 VDD.n1706 VDD.n124 8.77616
R776 VDD.n1706 VDD.n122 8.77616
R777 VDD.n1706 VDD.n120 8.77616
R778 VDD.n1706 VDD.n115 8.77616
R779 VDD.n1706 VDD.n106 8.77616
R780 VDD.n1706 VDD.n97 8.77616
R781 VDD.n1706 VDD.n88 8.77616
R782 VDD.n1706 VDD.n83 8.77616
R783 VDD.n1008 VDD.t7 8.11362
R784 VDD.t14 VDD.n1732 8.11362
R785 VDD.n1002 VDD.t17 7.19515
R786 VDD.n1733 VDD.n35 6.73592
R787 VDD.n1001 VDD.n35 6.12361
R788 VDD.n1030 VDD.n118 5.63319
R789 VDD.n1706 VDD.n87 5.63319
R790 VDD.n1706 VDD.n91 5.63319
R791 VDD.n1706 VDD.n90 5.63319
R792 VDD.n1706 VDD.n89 5.63319
R793 VDD.n1706 VDD.n96 5.63319
R794 VDD.n1706 VDD.n100 5.63319
R795 VDD.n1706 VDD.n99 5.63319
R796 VDD.n1706 VDD.n98 5.63319
R797 VDD.n1706 VDD.n105 5.63319
R798 VDD.n1706 VDD.n109 5.63319
R799 VDD.n1706 VDD.n108 5.63319
R800 VDD.n1706 VDD.n107 5.63319
R801 VDD.n1706 VDD.n114 5.63319
R802 VDD.n1706 VDD.n117 5.63319
R803 VDD.n1706 VDD.n116 5.63319
R804 VDD.n1707 VDD.n1706 5.1329
R805 VDD.n1706 VDD.n119 5.1329
R806 VDD.n1733 VDD.t14 4.74591
R807 VDD.n7 VDD.n1 4.6505
R808 VDD.n1747 VDD.n1746 4.6505
R809 VDD.n1740 VDD.n1739 4.59283
R810 VDD.n1710 VDD.n1709 4.54027
R811 VDD.n1087 VDD.n863 4.54027
R812 VDD.n47 VDD.n46 4.52882
R813 VDD.n188 VDD.n80 4.5005
R814 VDD.n81 VDD.n80 4.5005
R815 VDD.n193 VDD.n192 4.5005
R816 VDD.n212 VDD.n211 4.5005
R817 VDD.n1666 VDD.n1665 4.5005
R818 VDD.n250 VDD.n248 4.5005
R819 VDD.n356 VDD.n349 4.5005
R820 VDD.n355 VDD.n354 4.5005
R821 VDD.n332 VDD.n330 4.5005
R822 VDD.n1585 VDD.n1584 4.5005
R823 VDD.n1585 VDD.n329 4.5005
R824 VDD.n1597 VDD.n1596 4.5005
R825 VDD.n308 VDD.n306 4.5005
R826 VDD.n1619 VDD.n1618 4.5005
R827 VDD.n1619 VDD.n305 4.5005
R828 VDD.n1631 VDD.n1630 4.5005
R829 VDD.n275 VDD.n273 4.5005
R830 VDD.n1653 VDD.n1652 4.5005
R831 VDD.n1653 VDD.n272 4.5005
R832 VDD.n291 VDD.n290 4.5005
R833 VDD.n1664 VDD.n268 4.5005
R834 VDD.n1663 VDD.n1662 4.5005
R835 VDD.n1662 VDD.n1661 4.5005
R836 VDD.n315 VDD.n303 4.5005
R837 VDD.n1634 VDD.n1633 4.5005
R838 VDD.n302 VDD.n300 4.5005
R839 VDD.n304 VDD.n302 4.5005
R840 VDD.n339 VDD.n327 4.5005
R841 VDD.n1600 VDD.n1599 4.5005
R842 VDD.n326 VDD.n324 4.5005
R843 VDD.n328 VDD.n326 4.5005
R844 VDD.n1503 VDD.n1502 4.5005
R845 VDD.n430 VDD.n429 4.5005
R846 VDD.n533 VDD.n526 4.5005
R847 VDD.n532 VDD.n531 4.5005
R848 VDD.n509 VDD.n507 4.5005
R849 VDD.n1422 VDD.n1421 4.5005
R850 VDD.n1422 VDD.n506 4.5005
R851 VDD.n1434 VDD.n1433 4.5005
R852 VDD.n485 VDD.n483 4.5005
R853 VDD.n1456 VDD.n1455 4.5005
R854 VDD.n1456 VDD.n482 4.5005
R855 VDD.n1468 VDD.n1467 4.5005
R856 VDD.n452 VDD.n450 4.5005
R857 VDD.n1490 VDD.n1489 4.5005
R858 VDD.n1490 VDD.n449 4.5005
R859 VDD.n468 VDD.n467 4.5005
R860 VDD.n1501 VDD.n445 4.5005
R861 VDD.n1500 VDD.n1499 4.5005
R862 VDD.n1499 VDD.n1498 4.5005
R863 VDD.n492 VDD.n480 4.5005
R864 VDD.n1471 VDD.n1470 4.5005
R865 VDD.n479 VDD.n477 4.5005
R866 VDD.n481 VDD.n479 4.5005
R867 VDD.n516 VDD.n504 4.5005
R868 VDD.n1437 VDD.n1436 4.5005
R869 VDD.n503 VDD.n501 4.5005
R870 VDD.n505 VDD.n503 4.5005
R871 VDD.n1340 VDD.n1339 4.5005
R872 VDD.n607 VDD.n606 4.5005
R873 VDD.n710 VDD.n703 4.5005
R874 VDD.n709 VDD.n708 4.5005
R875 VDD.n686 VDD.n684 4.5005
R876 VDD.n1259 VDD.n1258 4.5005
R877 VDD.n1259 VDD.n683 4.5005
R878 VDD.n1271 VDD.n1270 4.5005
R879 VDD.n662 VDD.n660 4.5005
R880 VDD.n1293 VDD.n1292 4.5005
R881 VDD.n1293 VDD.n659 4.5005
R882 VDD.n1305 VDD.n1304 4.5005
R883 VDD.n629 VDD.n627 4.5005
R884 VDD.n1327 VDD.n1326 4.5005
R885 VDD.n1327 VDD.n626 4.5005
R886 VDD.n645 VDD.n644 4.5005
R887 VDD.n1338 VDD.n622 4.5005
R888 VDD.n1337 VDD.n1336 4.5005
R889 VDD.n1336 VDD.n1335 4.5005
R890 VDD.n669 VDD.n657 4.5005
R891 VDD.n1308 VDD.n1307 4.5005
R892 VDD.n656 VDD.n654 4.5005
R893 VDD.n658 VDD.n656 4.5005
R894 VDD.n693 VDD.n681 4.5005
R895 VDD.n1274 VDD.n1273 4.5005
R896 VDD.n680 VDD.n678 4.5005
R897 VDD.n682 VDD.n680 4.5005
R898 VDD.n1177 VDD.n1176 4.5005
R899 VDD.n784 VDD.n783 4.5005
R900 VDD.n864 VDD.n861 4.5005
R901 VDD.n1108 VDD.n1107 4.5005
R902 VDD.n839 VDD.n837 4.5005
R903 VDD.n1130 VDD.n1129 4.5005
R904 VDD.n1130 VDD.n836 4.5005
R905 VDD.n1142 VDD.n1141 4.5005
R906 VDD.n806 VDD.n804 4.5005
R907 VDD.n1164 VDD.n1163 4.5005
R908 VDD.n1164 VDD.n803 4.5005
R909 VDD.n822 VDD.n821 4.5005
R910 VDD.n1175 VDD.n799 4.5005
R911 VDD.n1174 VDD.n1173 4.5005
R912 VDD.n1173 VDD.n1172 4.5005
R913 VDD.n846 VDD.n834 4.5005
R914 VDD.n1145 VDD.n1144 4.5005
R915 VDD.n833 VDD.n831 4.5005
R916 VDD.n835 VDD.n833 4.5005
R917 VDD.n871 VDD.n858 4.5005
R918 VDD.n1111 VDD.n1110 4.5005
R919 VDD.n857 VDD.n855 4.5005
R920 VDD.n859 VDD.n857 4.5005
R921 VDD.n1096 VDD.n1095 4.5005
R922 VDD.n1096 VDD.n860 4.5005
R923 VDD.n723 VDD.n722 4.5005
R924 VDD.n1189 VDD.n1188 4.5005
R925 VDD.n770 VDD.n769 4.5005
R926 VDD.n780 VDD.n778 4.5005
R927 VDD.n1192 VDD.n780 4.5005
R928 VDD.n1203 VDD.n1202 4.5005
R929 VDD.n754 VDD.n753 4.5005
R930 VDD.n764 VDD.n762 4.5005
R931 VDD.n1206 VDD.n764 4.5005
R932 VDD.n1215 VDD.n1214 4.5005
R933 VDD.n738 VDD.n737 4.5005
R934 VDD.n748 VDD.n746 4.5005
R935 VDD.n1218 VDD.n748 4.5005
R936 VDD.n732 VDD.n730 4.5005
R937 VDD.n1230 VDD.n732 4.5005
R938 VDD.n1227 VDD.n1226 4.5005
R939 VDD.n794 VDD.n792 4.5005
R940 VDD.n1180 VDD.n794 4.5005
R941 VDD.n711 VDD.n704 4.5005
R942 VDD.n1242 VDD.n711 4.5005
R943 VDD.n1239 VDD.n1238 4.5005
R944 VDD.n546 VDD.n545 4.5005
R945 VDD.n1352 VDD.n1351 4.5005
R946 VDD.n593 VDD.n592 4.5005
R947 VDD.n603 VDD.n601 4.5005
R948 VDD.n1355 VDD.n603 4.5005
R949 VDD.n1366 VDD.n1365 4.5005
R950 VDD.n577 VDD.n576 4.5005
R951 VDD.n587 VDD.n585 4.5005
R952 VDD.n1369 VDD.n587 4.5005
R953 VDD.n1378 VDD.n1377 4.5005
R954 VDD.n561 VDD.n560 4.5005
R955 VDD.n571 VDD.n569 4.5005
R956 VDD.n1381 VDD.n571 4.5005
R957 VDD.n555 VDD.n553 4.5005
R958 VDD.n1393 VDD.n555 4.5005
R959 VDD.n1390 VDD.n1389 4.5005
R960 VDD.n617 VDD.n615 4.5005
R961 VDD.n1343 VDD.n617 4.5005
R962 VDD.n534 VDD.n527 4.5005
R963 VDD.n1405 VDD.n534 4.5005
R964 VDD.n1402 VDD.n1401 4.5005
R965 VDD.n369 VDD.n368 4.5005
R966 VDD.n1515 VDD.n1514 4.5005
R967 VDD.n416 VDD.n415 4.5005
R968 VDD.n426 VDD.n424 4.5005
R969 VDD.n1518 VDD.n426 4.5005
R970 VDD.n1529 VDD.n1528 4.5005
R971 VDD.n400 VDD.n399 4.5005
R972 VDD.n410 VDD.n408 4.5005
R973 VDD.n1532 VDD.n410 4.5005
R974 VDD.n1541 VDD.n1540 4.5005
R975 VDD.n384 VDD.n383 4.5005
R976 VDD.n394 VDD.n392 4.5005
R977 VDD.n1544 VDD.n394 4.5005
R978 VDD.n378 VDD.n376 4.5005
R979 VDD.n1556 VDD.n378 4.5005
R980 VDD.n1553 VDD.n1552 4.5005
R981 VDD.n440 VDD.n438 4.5005
R982 VDD.n1506 VDD.n440 4.5005
R983 VDD.n357 VDD.n350 4.5005
R984 VDD.n1568 VDD.n357 4.5005
R985 VDD.n1565 VDD.n1564 4.5005
R986 VDD.n214 VDD.n163 4.5005
R987 VDD.n1678 VDD.n1677 4.5005
R988 VDD.n1687 VDD.n1686 4.5005
R989 VDD.n249 VDD.n233 4.5005
R990 VDD.n1681 VDD.n233 4.5005
R991 VDD.n231 VDD.n229 4.5005
R992 VDD.n1698 VDD.n1697 4.5005
R993 VDD.n241 VDD.n240 4.5005
R994 VDD.n241 VDD.n239 4.5005
R995 VDD.n1702 VDD.n1701 4.5005
R996 VDD.n1702 VDD.n162 4.5005
R997 VDD.n1700 VDD.n1699 4.5005
R998 VDD.n263 VDD.n261 4.5005
R999 VDD.n1669 VDD.n263 4.5005
R1000 VDD.n176 VDD.n175 4.5005
R1001 VDD.n177 VDD.n176 4.5005
R1002 VDD.n194 VDD.n180 4.5005
R1003 VDD.n1025 VDD.n1024 4.5005
R1004 VDD.n972 VDD.n965 4.5005
R1005 VDD.n895 VDD.n880 4.5005
R1006 VDD.n914 VDD.n887 4.5005
R1007 VDD.n898 VDD.n897 4.5005
R1008 VDD.n934 VDD.n933 4.5005
R1009 VDD.n907 VDD.n905 4.5005
R1010 VDD.n953 VDD.n926 4.5005
R1011 VDD.n937 VDD.n936 4.5005
R1012 VDD.n1022 VDD.n1021 4.5005
R1013 VDD.n946 VDD.n944 4.5005
R1014 VDD.n964 VDD.n962 4.5005
R1015 VDD.n966 VDD.n964 4.5005
R1016 VDD.n886 VDD.n884 4.5005
R1017 VDD.n888 VDD.n886 4.5005
R1018 VDD.n1066 VDD.n1065 4.5005
R1019 VDD.n1066 VDD.n904 4.5005
R1020 VDD.n925 VDD.n923 4.5005
R1021 VDD.n927 VDD.n925 4.5005
R1022 VDD.n1045 VDD.n1044 4.5005
R1023 VDD.n1045 VDD.n943 4.5005
R1024 VDD.n27 VDD.n26 4.5005
R1025 VDD.n9 VDD.n6 4.5005
R1026 VDD.n10 VDD.n8 4.5005
R1027 VDD.n1732 VDD.n1731 4.43975
R1028 VDD VDD.n118 4.28667
R1029 VDD.n1012 VDD.n1011 4.20505
R1030 VDD.n1011 VDD.n1010 4.20505
R1031 VDD.n1739 VDD.n1738 4.20505
R1032 VDD.n1736 VDD.n29 4.20505
R1033 VDD.n1732 VDD.n29 4.20505
R1034 VDD.n1735 VDD.n1734 4.20505
R1035 VDD.n1734 VDD.n1733 4.20505
R1036 VDD.n34 VDD.n33 4.20505
R1037 VDD.n1001 VDD.n34 4.20505
R1038 VDD.n1004 VDD.n1003 4.20505
R1039 VDD.n1003 VDD.n1002 4.20505
R1040 VDD.n1006 VDD.n1005 4.20505
R1041 VDD.n1007 VDD.n1006 4.20505
R1042 VDD.n989 VDD.n988 4.20505
R1043 VDD.n1008 VDD.n989 4.20505
R1044 VDD.n1738 VDD.n1737 3.56608
R1045 VDD.t17 VDD.n1001 3.52129
R1046 VDD.n1749 VDD.n25 3.46788
R1047 VDD.n20 VDD.n19 3.46651
R1048 VDD.n53 VDD.n52 3.46323
R1049 VDD.n48 VDD.n42 3.46321
R1050 VDD.n1729 VDD.n37 3.45407
R1051 VDD.n63 VDD.n62 3.45407
R1052 VDD.n998 VDD.n67 3.45407
R1053 VDD.n995 VDD.n71 3.45407
R1054 VDD.n991 VDD.n75 3.45407
R1055 VDD.n38 VDD.n36 3.45149
R1056 VDD.n60 VDD.n58 3.45149
R1057 VDD.n997 VDD.n65 3.45149
R1058 VDD.n994 VDD.n69 3.45149
R1059 VDD.n990 VDD.n73 3.45149
R1060 VDD.n1086 VDD.n1085 3.42985
R1061 VDD.n13 VDD.n10 3.4257
R1062 VDD.n984 VDD.n969 3.42443
R1063 VDD.n1711 VDD.n1710 3.42376
R1064 VDD.n1088 VDD.n1087 3.42376
R1065 VDD.n44 VDD.n41 3.41853
R1066 VDD.n26 VDD.n11 3.41388
R1067 VDD.n1089 VDD.n1088 3.41326
R1068 VDD.n1712 VDD.n1711 3.41257
R1069 VDD.n53 VDD.n39 3.41218
R1070 VDD.n1725 VDD.n37 3.41218
R1071 VDD.n63 VDD.n57 3.41218
R1072 VDD.n67 VDD.n64 3.41218
R1073 VDD.n71 VDD.n68 3.41218
R1074 VDD.n75 VDD.n72 3.41218
R1075 VDD.n43 VDD.n40 3.41162
R1076 VDD.n196 VDD.n195 3.4105
R1077 VDD.n203 VDD.n202 3.4105
R1078 VDD.n280 VDD.n269 3.4105
R1079 VDD.n1651 VDD.n1650 3.4105
R1080 VDD.n1643 VDD.n1642 3.4105
R1081 VDD.n1617 VDD.n1616 3.4105
R1082 VDD.n1609 VDD.n1608 3.4105
R1083 VDD.n1583 VDD.n1582 3.4105
R1084 VDD.n352 VDD.n346 3.4105
R1085 VDD.n457 VDD.n446 3.4105
R1086 VDD.n1488 VDD.n1487 3.4105
R1087 VDD.n1480 VDD.n1479 3.4105
R1088 VDD.n1454 VDD.n1453 3.4105
R1089 VDD.n1446 VDD.n1445 3.4105
R1090 VDD.n1420 VDD.n1419 3.4105
R1091 VDD.n529 VDD.n523 3.4105
R1092 VDD.n634 VDD.n623 3.4105
R1093 VDD.n1325 VDD.n1324 3.4105
R1094 VDD.n1317 VDD.n1316 3.4105
R1095 VDD.n1291 VDD.n1290 3.4105
R1096 VDD.n1283 VDD.n1282 3.4105
R1097 VDD.n1257 VDD.n1256 3.4105
R1098 VDD.n706 VDD.n700 3.4105
R1099 VDD.n811 VDD.n800 3.4105
R1100 VDD.n1162 VDD.n1161 3.4105
R1101 VDD.n1154 VDD.n1153 3.4105
R1102 VDD.n1128 VDD.n1127 3.4105
R1103 VDD.n1120 VDD.n1119 3.4105
R1104 VDD.n1094 VDD.n1093 3.4105
R1105 VDD.n873 VDD.n872 3.4105
R1106 VDD.n1109 VDD.n853 3.4105
R1107 VDD.n848 VDD.n847 3.4105
R1108 VDD.n1143 VDD.n829 3.4105
R1109 VDD.n824 VDD.n823 3.4105
R1110 VDD.n1197 VDD.n779 3.4105
R1111 VDD.n1201 VDD.n1200 3.4105
R1112 VDD.n1209 VDD.n763 3.4105
R1113 VDD.n1213 VDD.n1212 3.4105
R1114 VDD.n1221 VDD.n747 3.4105
R1115 VDD.n1225 VDD.n1224 3.4105
R1116 VDD.n1233 VDD.n731 3.4105
R1117 VDD.n1237 VDD.n1236 3.4105
R1118 VDD.n1187 VDD.n1186 3.4105
R1119 VDD.n1183 VDD.n793 3.4105
R1120 VDD.n1245 VDD.n705 3.4105
R1121 VDD.n707 VDD.n699 3.4105
R1122 VDD.n695 VDD.n694 3.4105
R1123 VDD.n1272 VDD.n676 3.4105
R1124 VDD.n671 VDD.n670 3.4105
R1125 VDD.n1306 VDD.n652 3.4105
R1126 VDD.n647 VDD.n646 3.4105
R1127 VDD.n1360 VDD.n602 3.4105
R1128 VDD.n1364 VDD.n1363 3.4105
R1129 VDD.n1372 VDD.n586 3.4105
R1130 VDD.n1376 VDD.n1375 3.4105
R1131 VDD.n1384 VDD.n570 3.4105
R1132 VDD.n1388 VDD.n1387 3.4105
R1133 VDD.n1396 VDD.n554 3.4105
R1134 VDD.n1400 VDD.n1399 3.4105
R1135 VDD.n1350 VDD.n1349 3.4105
R1136 VDD.n1346 VDD.n616 3.4105
R1137 VDD.n1408 VDD.n528 3.4105
R1138 VDD.n530 VDD.n522 3.4105
R1139 VDD.n518 VDD.n517 3.4105
R1140 VDD.n1435 VDD.n499 3.4105
R1141 VDD.n494 VDD.n493 3.4105
R1142 VDD.n1469 VDD.n475 3.4105
R1143 VDD.n470 VDD.n469 3.4105
R1144 VDD.n1523 VDD.n425 3.4105
R1145 VDD.n1527 VDD.n1526 3.4105
R1146 VDD.n1535 VDD.n409 3.4105
R1147 VDD.n1539 VDD.n1538 3.4105
R1148 VDD.n1547 VDD.n393 3.4105
R1149 VDD.n1551 VDD.n1550 3.4105
R1150 VDD.n1559 VDD.n377 3.4105
R1151 VDD.n1563 VDD.n1562 3.4105
R1152 VDD.n1513 VDD.n1512 3.4105
R1153 VDD.n1509 VDD.n439 3.4105
R1154 VDD.n1571 VDD.n351 3.4105
R1155 VDD.n353 VDD.n345 3.4105
R1156 VDD.n341 VDD.n340 3.4105
R1157 VDD.n1598 VDD.n322 3.4105
R1158 VDD.n317 VDD.n316 3.4105
R1159 VDD.n1632 VDD.n298 3.4105
R1160 VDD.n293 VDD.n292 3.4105
R1161 VDD.n256 VDD.n232 3.4105
R1162 VDD.n1689 VDD.n1688 3.4105
R1163 VDD.n227 VDD.n168 3.4105
R1164 VDD.n169 VDD.n166 3.4105
R1165 VDD.n222 VDD.n164 3.4105
R1166 VDD.n216 VDD.n215 3.4105
R1167 VDD.n1676 VDD.n1675 3.4105
R1168 VDD.n1672 VDD.n262 3.4105
R1169 VDD.n186 VDD.n79 3.4105
R1170 VDD.n44 VDD.n43 3.4105
R1171 VDD.n49 VDD.n48 3.4105
R1172 VDD.n1714 VDD.n1713 3.4105
R1173 VDD.n1715 VDD.n1714 3.4105
R1174 VDD.n1717 VDD.n1716 3.4105
R1175 VDD.n1718 VDD.n1717 3.4105
R1176 VDD.n1720 VDD.n1719 3.4105
R1177 VDD.n1721 VDD.n1720 3.4105
R1178 VDD.n1723 VDD.n1722 3.4105
R1179 VDD.n1724 VDD.n1723 3.4105
R1180 VDD.n1727 VDD.n1726 3.4105
R1181 VDD.n1727 VDD.n56 3.4105
R1182 VDD.n55 VDD.n54 3.4105
R1183 VDD.n54 VDD.n50 3.4105
R1184 VDD.n77 VDD.n76 3.4105
R1185 VDD.n187 VDD.n183 3.4105
R1186 VDD.n174 VDD.n173 3.4105
R1187 VDD.n876 VDD.n866 3.4105
R1188 VDD.n1090 VDD.n867 3.4105
R1189 VDD.n875 VDD.n874 3.4105
R1190 VDD.n1121 VDD.n852 3.4105
R1191 VDD.n870 VDD.n869 3.4105
R1192 VDD.n1123 VDD.n1122 3.4105
R1193 VDD.n851 VDD.n841 3.4105
R1194 VDD.n1124 VDD.n842 3.4105
R1195 VDD.n850 VDD.n849 3.4105
R1196 VDD.n1155 VDD.n828 3.4105
R1197 VDD.n845 VDD.n844 3.4105
R1198 VDD.n1157 VDD.n1156 3.4105
R1199 VDD.n827 VDD.n808 3.4105
R1200 VDD.n1158 VDD.n809 3.4105
R1201 VDD.n826 VDD.n825 3.4105
R1202 VDD.n816 VDD.n815 3.4105
R1203 VDD.n819 VDD.n810 3.4105
R1204 VDD.n743 VDD.n742 3.4105
R1205 VDD.n728 VDD.n724 3.4105
R1206 VDD.n1235 VDD.n729 3.4105
R1207 VDD.n759 VDD.n758 3.4105
R1208 VDD.n744 VDD.n739 3.4105
R1209 VDD.n1223 VDD.n745 3.4105
R1210 VDD.n775 VDD.n774 3.4105
R1211 VDD.n760 VDD.n755 3.4105
R1212 VDD.n1211 VDD.n761 3.4105
R1213 VDD.n789 VDD.n788 3.4105
R1214 VDD.n776 VDD.n771 3.4105
R1215 VDD.n1199 VDD.n777 3.4105
R1216 VDD.n814 VDD.n813 3.4105
R1217 VDD.n790 VDD.n785 3.4105
R1218 VDD.n1185 VDD.n791 3.4105
R1219 VDD.n727 VDD.n726 3.4105
R1220 VDD.n1250 VDD.n1249 3.4105
R1221 VDD.n1248 VDD.n1247 3.4105
R1222 VDD.n1252 VDD.n1251 3.4105
R1223 VDD.n698 VDD.n688 3.4105
R1224 VDD.n1253 VDD.n689 3.4105
R1225 VDD.n697 VDD.n696 3.4105
R1226 VDD.n1284 VDD.n675 3.4105
R1227 VDD.n692 VDD.n691 3.4105
R1228 VDD.n1286 VDD.n1285 3.4105
R1229 VDD.n674 VDD.n664 3.4105
R1230 VDD.n1287 VDD.n665 3.4105
R1231 VDD.n673 VDD.n672 3.4105
R1232 VDD.n1318 VDD.n651 3.4105
R1233 VDD.n668 VDD.n667 3.4105
R1234 VDD.n1320 VDD.n1319 3.4105
R1235 VDD.n650 VDD.n631 3.4105
R1236 VDD.n1321 VDD.n632 3.4105
R1237 VDD.n649 VDD.n648 3.4105
R1238 VDD.n639 VDD.n638 3.4105
R1239 VDD.n642 VDD.n633 3.4105
R1240 VDD.n566 VDD.n565 3.4105
R1241 VDD.n551 VDD.n547 3.4105
R1242 VDD.n1398 VDD.n552 3.4105
R1243 VDD.n582 VDD.n581 3.4105
R1244 VDD.n567 VDD.n562 3.4105
R1245 VDD.n1386 VDD.n568 3.4105
R1246 VDD.n598 VDD.n597 3.4105
R1247 VDD.n583 VDD.n578 3.4105
R1248 VDD.n1374 VDD.n584 3.4105
R1249 VDD.n612 VDD.n611 3.4105
R1250 VDD.n599 VDD.n594 3.4105
R1251 VDD.n1362 VDD.n600 3.4105
R1252 VDD.n637 VDD.n636 3.4105
R1253 VDD.n613 VDD.n608 3.4105
R1254 VDD.n1348 VDD.n614 3.4105
R1255 VDD.n550 VDD.n549 3.4105
R1256 VDD.n1413 VDD.n1412 3.4105
R1257 VDD.n1411 VDD.n1410 3.4105
R1258 VDD.n1415 VDD.n1414 3.4105
R1259 VDD.n521 VDD.n511 3.4105
R1260 VDD.n1416 VDD.n512 3.4105
R1261 VDD.n520 VDD.n519 3.4105
R1262 VDD.n1447 VDD.n498 3.4105
R1263 VDD.n515 VDD.n514 3.4105
R1264 VDD.n1449 VDD.n1448 3.4105
R1265 VDD.n497 VDD.n487 3.4105
R1266 VDD.n1450 VDD.n488 3.4105
R1267 VDD.n496 VDD.n495 3.4105
R1268 VDD.n1481 VDD.n474 3.4105
R1269 VDD.n491 VDD.n490 3.4105
R1270 VDD.n1483 VDD.n1482 3.4105
R1271 VDD.n473 VDD.n454 3.4105
R1272 VDD.n1484 VDD.n455 3.4105
R1273 VDD.n472 VDD.n471 3.4105
R1274 VDD.n462 VDD.n461 3.4105
R1275 VDD.n465 VDD.n456 3.4105
R1276 VDD.n389 VDD.n388 3.4105
R1277 VDD.n374 VDD.n370 3.4105
R1278 VDD.n1561 VDD.n375 3.4105
R1279 VDD.n405 VDD.n404 3.4105
R1280 VDD.n390 VDD.n385 3.4105
R1281 VDD.n1549 VDD.n391 3.4105
R1282 VDD.n421 VDD.n420 3.4105
R1283 VDD.n406 VDD.n401 3.4105
R1284 VDD.n1537 VDD.n407 3.4105
R1285 VDD.n435 VDD.n434 3.4105
R1286 VDD.n422 VDD.n417 3.4105
R1287 VDD.n1525 VDD.n423 3.4105
R1288 VDD.n460 VDD.n459 3.4105
R1289 VDD.n436 VDD.n431 3.4105
R1290 VDD.n1511 VDD.n437 3.4105
R1291 VDD.n373 VDD.n372 3.4105
R1292 VDD.n1576 VDD.n1575 3.4105
R1293 VDD.n1574 VDD.n1573 3.4105
R1294 VDD.n1578 VDD.n1577 3.4105
R1295 VDD.n344 VDD.n334 3.4105
R1296 VDD.n1579 VDD.n335 3.4105
R1297 VDD.n343 VDD.n342 3.4105
R1298 VDD.n1610 VDD.n321 3.4105
R1299 VDD.n338 VDD.n337 3.4105
R1300 VDD.n1612 VDD.n1611 3.4105
R1301 VDD.n320 VDD.n310 3.4105
R1302 VDD.n1613 VDD.n311 3.4105
R1303 VDD.n319 VDD.n318 3.4105
R1304 VDD.n1644 VDD.n297 3.4105
R1305 VDD.n314 VDD.n313 3.4105
R1306 VDD.n1646 VDD.n1645 3.4105
R1307 VDD.n296 VDD.n277 3.4105
R1308 VDD.n1647 VDD.n278 3.4105
R1309 VDD.n295 VDD.n294 3.4105
R1310 VDD.n285 VDD.n284 3.4105
R1311 VDD.n288 VDD.n279 3.4105
R1312 VDD.n223 VDD.n171 3.4105
R1313 VDD.n218 VDD.n217 3.4105
R1314 VDD.n219 VDD.n172 3.4105
R1315 VDD.n1692 VDD.n1691 3.4105
R1316 VDD.n225 VDD.n224 3.4105
R1317 VDD.n1695 VDD.n1694 3.4105
R1318 VDD.n258 VDD.n257 3.4105
R1319 VDD.n1690 VDD.n226 3.4105
R1320 VDD.n253 VDD.n228 3.4105
R1321 VDD.n283 VDD.n282 3.4105
R1322 VDD.n259 VDD.n251 3.4105
R1323 VDD.n1674 VDD.n260 3.4105
R1324 VDD.n199 VDD.n182 3.4105
R1325 VDD.n198 VDD.n197 3.4105
R1326 VDD.n979 VDD.n978 3.4105
R1327 VDD.n1036 VDD.n959 3.4105
R1328 VDD.n958 VDD.n948 3.4105
R1329 VDD.n1038 VDD.n1037 3.4105
R1330 VDD.n957 VDD.n956 3.4105
R1331 VDD.n1057 VDD.n920 3.4105
R1332 VDD.n919 VDD.n909 3.4105
R1333 VDD.n1059 VDD.n1058 3.4105
R1334 VDD.n918 VDD.n917 3.4105
R1335 VDD.n1078 VDD.n882 3.4105
R1336 VDD.n1080 VDD.n1079 3.4105
R1337 VDD.n981 VDD.n980 3.4105
R1338 VDD.n970 VDD.n968 3.4105
R1339 VDD.n974 VDD.n973 3.4105
R1340 VDD.n1039 VDD.n949 3.4105
R1341 VDD.n952 VDD.n951 3.4105
R1342 VDD.n1060 VDD.n910 3.4105
R1343 VDD.n913 VDD.n912 3.4105
R1344 VDD.n1085 VDD.n1084 3.4105
R1345 VDD.n896 VDD.n881 3.4105
R1346 VDD.n1023 VDD.n960 3.4105
R1347 VDD.n1043 VDD.n1042 3.4105
R1348 VDD.n955 VDD.n954 3.4105
R1349 VDD.n1056 VDD.n1055 3.4105
R1350 VDD.n935 VDD.n921 3.4105
R1351 VDD.n1064 VDD.n1063 3.4105
R1352 VDD.n916 VDD.n915 3.4105
R1353 VDD.n1077 VDD.n1076 3.4105
R1354 VDD.n1082 VDD.n1081 3.4105
R1355 VDD.n977 VDD.n976 3.4105
R1356 VDD.n1035 VDD.n1034 3.4105
R1357 VDD.n1753 VDD.n1752 3.4105
R1358 VDD.n16 VDD.n15 3.4105
R1359 VDD.n18 VDD.n17 3.4105
R1360 VDD.n1751 VDD.n23 3.4105
R1361 VDD.n22 VDD.n21 3.4105
R1362 VDD.n1755 VDD.n1754 3.4105
R1363 VDD.n24 VDD.n22 3.4105
R1364 VDD.n1138 VDD.n116 3.38568
R1365 VDD.n1104 VDD.n117 3.38568
R1366 VDD.n1301 VDD.n107 3.38568
R1367 VDD.n1267 VDD.n108 3.38568
R1368 VDD.n713 VDD.n109 3.38568
R1369 VDD.n1464 VDD.n98 3.38568
R1370 VDD.n1430 VDD.n99 3.38568
R1371 VDD.n536 VDD.n100 3.38568
R1372 VDD.n1627 VDD.n89 3.38568
R1373 VDD.n1593 VDD.n90 3.38568
R1374 VDD.n359 VDD.n91 3.38568
R1375 VDD.n1031 VDD.n1030 3.38568
R1376 VDD.n1194 VDD.n114 3.38568
R1377 VDD.n1357 VDD.n105 3.38568
R1378 VDD.n1520 VDD.n96 3.38568
R1379 VDD.n1683 VDD.n87 3.38568
R1380 VDD.t7 VDD.n1007 3.21513
R1381 VDD.n190 VDD.n81 3.10353
R1382 VDD.n189 VDD.n179 3.10353
R1383 VDD.n209 VDD.n177 3.10353
R1384 VDD.n208 VDD.n161 3.10353
R1385 VDD.n234 VDD.n162 3.10353
R1386 VDD.n237 VDD.n235 3.10353
R1387 VDD.n243 VDD.n239 3.10353
R1388 VDD.n246 VDD.n245 3.10353
R1389 VDD.n1681 VDD.n1680 3.10353
R1390 VDD.n266 VDD.n247 3.10353
R1391 VDD.n1669 VDD.n1668 3.10353
R1392 VDD.n1661 VDD.n267 3.10353
R1393 VDD.n1659 VDD.n1656 3.10353
R1394 VDD.n1655 VDD.n272 3.10353
R1395 VDD.n1637 VDD.n1629 3.10353
R1396 VDD.n1636 VDD.n304 3.10353
R1397 VDD.n1625 VDD.n1622 3.10353
R1398 VDD.n1621 VDD.n305 3.10353
R1399 VDD.n1603 VDD.n1595 3.10353
R1400 VDD.n1602 VDD.n328 3.10353
R1401 VDD.n1591 VDD.n1588 3.10353
R1402 VDD.n1587 VDD.n329 3.10353
R1403 VDD.n362 VDD.n361 3.10353
R1404 VDD.n365 VDD.n363 3.10353
R1405 VDD.n1568 VDD.n1567 3.10353
R1406 VDD.n380 VDD.n367 3.10353
R1407 VDD.n1556 VDD.n1555 3.10353
R1408 VDD.n396 VDD.n382 3.10353
R1409 VDD.n1544 VDD.n1543 3.10353
R1410 VDD.n412 VDD.n398 3.10353
R1411 VDD.n1532 VDD.n1531 3.10353
R1412 VDD.n427 VDD.n414 3.10353
R1413 VDD.n1518 VDD.n1517 3.10353
R1414 VDD.n443 VDD.n428 3.10353
R1415 VDD.n1506 VDD.n1505 3.10353
R1416 VDD.n1498 VDD.n444 3.10353
R1417 VDD.n1496 VDD.n1493 3.10353
R1418 VDD.n1492 VDD.n449 3.10353
R1419 VDD.n1474 VDD.n1466 3.10353
R1420 VDD.n1473 VDD.n481 3.10353
R1421 VDD.n1462 VDD.n1459 3.10353
R1422 VDD.n1458 VDD.n482 3.10353
R1423 VDD.n1440 VDD.n1432 3.10353
R1424 VDD.n1439 VDD.n505 3.10353
R1425 VDD.n1428 VDD.n1425 3.10353
R1426 VDD.n1424 VDD.n506 3.10353
R1427 VDD.n539 VDD.n538 3.10353
R1428 VDD.n542 VDD.n540 3.10353
R1429 VDD.n1405 VDD.n1404 3.10353
R1430 VDD.n557 VDD.n544 3.10353
R1431 VDD.n1393 VDD.n1392 3.10353
R1432 VDD.n573 VDD.n559 3.10353
R1433 VDD.n1381 VDD.n1380 3.10353
R1434 VDD.n589 VDD.n575 3.10353
R1435 VDD.n1369 VDD.n1368 3.10353
R1436 VDD.n604 VDD.n591 3.10353
R1437 VDD.n1355 VDD.n1354 3.10353
R1438 VDD.n620 VDD.n605 3.10353
R1439 VDD.n1343 VDD.n1342 3.10353
R1440 VDD.n1335 VDD.n621 3.10353
R1441 VDD.n1333 VDD.n1330 3.10353
R1442 VDD.n1329 VDD.n626 3.10353
R1443 VDD.n1311 VDD.n1303 3.10353
R1444 VDD.n1310 VDD.n658 3.10353
R1445 VDD.n1299 VDD.n1296 3.10353
R1446 VDD.n1295 VDD.n659 3.10353
R1447 VDD.n1277 VDD.n1269 3.10353
R1448 VDD.n1276 VDD.n682 3.10353
R1449 VDD.n1265 VDD.n1262 3.10353
R1450 VDD.n1261 VDD.n683 3.10353
R1451 VDD.n716 VDD.n715 3.10353
R1452 VDD.n719 VDD.n717 3.10353
R1453 VDD.n1242 VDD.n1241 3.10353
R1454 VDD.n734 VDD.n721 3.10353
R1455 VDD.n1230 VDD.n1229 3.10353
R1456 VDD.n750 VDD.n736 3.10353
R1457 VDD.n1218 VDD.n1217 3.10353
R1458 VDD.n766 VDD.n752 3.10353
R1459 VDD.n1206 VDD.n1205 3.10353
R1460 VDD.n781 VDD.n768 3.10353
R1461 VDD.n1192 VDD.n1191 3.10353
R1462 VDD.n797 VDD.n782 3.10353
R1463 VDD.n1180 VDD.n1179 3.10353
R1464 VDD.n1172 VDD.n798 3.10353
R1465 VDD.n1170 VDD.n1167 3.10353
R1466 VDD.n1166 VDD.n803 3.10353
R1467 VDD.n1148 VDD.n1140 3.10353
R1468 VDD.n1147 VDD.n835 3.10353
R1469 VDD.n1136 VDD.n1133 3.10353
R1470 VDD.n1132 VDD.n836 3.10353
R1471 VDD.n1114 VDD.n1106 3.10353
R1472 VDD.n1113 VDD.n859 3.10353
R1473 VDD.n1102 VDD.n1099 3.10353
R1474 VDD.n1098 VDD.n860 3.10353
R1475 VDD.n901 VDD.n894 3.10353
R1476 VDD.n900 VDD.n888 3.10353
R1477 VDD.n1069 VDD.n889 3.10353
R1478 VDD.n1068 VDD.n904 3.10353
R1479 VDD.n940 VDD.n932 3.10353
R1480 VDD.n939 VDD.n927 3.10353
R1481 VDD.n1048 VDD.n928 3.10353
R1482 VDD.n1047 VDD.n943 3.10353
R1483 VDD.n1028 VDD.n1020 3.10353
R1484 VDD.n1027 VDD.n966 3.10353
R1485 VDD.n6 VDD.n5 3.03311
R1486 VDD VDD.n993 2.90898
R1487 VDD.n1731 VDD 2.7559
R1488 VDD.n1761 VDD.n1760 2.5605
R1489 VDD.n891 VDD.n879 2.5429
R1490 VDD.n1745 VDD.n5 2.36358
R1491 VDD.n1014 VDD.n967 2.28608
R1492 VDD.n1730 VDD.n36 2.24869
R1493 VDD.n61 VDD.n60 2.24869
R1494 VDD.n999 VDD.n997 2.24869
R1495 VDD.n996 VDD.n994 2.24869
R1496 VDD.n992 VDD.n990 2.24869
R1497 VDD.n1014 VDD.n1013 2.15377
R1498 VDD.n1010 VDD.n1009 1.99051
R1499 VDD.n986 VDD.n985 1.94045
R1500 VDD.n19 VDD.n0 1.94045
R1501 VDD.n1749 VDD.n1748 1.94045
R1502 VDD.n1139 VDD.n1138 1.76521
R1503 VDD.n1105 VDD.n1104 1.76521
R1504 VDD.n718 VDD.n128 1.76521
R1505 VDD.n733 VDD.n110 1.76521
R1506 VDD.n749 VDD.n126 1.76521
R1507 VDD.n765 VDD.n112 1.76521
R1508 VDD.n1194 VDD.n1193 1.76521
R1509 VDD.n1302 VDD.n1301 1.76521
R1510 VDD.n1268 VDD.n1267 1.76521
R1511 VDD.n714 VDD.n713 1.76521
R1512 VDD.n541 VDD.n139 1.76521
R1513 VDD.n556 VDD.n101 1.76521
R1514 VDD.n572 VDD.n137 1.76521
R1515 VDD.n588 VDD.n103 1.76521
R1516 VDD.n1357 VDD.n1356 1.76521
R1517 VDD.n1465 VDD.n1464 1.76521
R1518 VDD.n1431 VDD.n1430 1.76521
R1519 VDD.n537 VDD.n536 1.76521
R1520 VDD.n364 VDD.n150 1.76521
R1521 VDD.n379 VDD.n92 1.76521
R1522 VDD.n395 VDD.n148 1.76521
R1523 VDD.n411 VDD.n94 1.76521
R1524 VDD.n1520 VDD.n1519 1.76521
R1525 VDD.n1628 VDD.n1627 1.76521
R1526 VDD.n1594 VDD.n1593 1.76521
R1527 VDD.n360 VDD.n359 1.76521
R1528 VDD.n1705 VDD.n159 1.76521
R1529 VDD.n236 VDD.n85 1.76521
R1530 VDD.n1683 VDD.n1682 1.76521
R1531 VDD.n893 VDD.n892 1.76521
R1532 VDD.n1031 VDD.n1016 1.76521
R1533 VDD.n993 VDD.t3 1.68435
R1534 VDD.n1072 VDD.n1071 1.66612
R1535 VDD.n930 VDD.n929 1.66612
R1536 VDD.n1051 VDD.n1050 1.66612
R1537 VDD.n1018 VDD.n1017 1.66612
R1538 VDD.n1658 VDD.n157 1.66612
R1539 VDD.n1624 VDD.n155 1.66612
R1540 VDD.n1590 VDD.n153 1.66612
R1541 VDD.n1495 VDD.n146 1.66612
R1542 VDD.n1461 VDD.n144 1.66612
R1543 VDD.n1427 VDD.n142 1.66612
R1544 VDD.n1332 VDD.n135 1.66612
R1545 VDD.n1298 VDD.n133 1.66612
R1546 VDD.n1264 VDD.n131 1.66612
R1547 VDD.n1169 VDD.n124 1.66612
R1548 VDD.n1135 VDD.n122 1.66612
R1549 VDD.n1101 VDD.n120 1.66612
R1550 VDD.n796 VDD.n115 1.66612
R1551 VDD.n619 VDD.n106 1.66612
R1552 VDD.n442 VDD.n97 1.66612
R1553 VDD.n265 VDD.n88 1.66612
R1554 VDD.n178 VDD.n83 1.66612
R1555 VDD.n1007 VDD.n1000 1.53128
R1556 VDD.n1034 VDD.n1033 1.35607
R1557 VDD.n204 VDD.n203 1.35607
R1558 VDD.n271 VDD.n269 1.35607
R1559 VDD.n1651 VDD.n274 1.35607
R1560 VDD.n1642 VDD.n1641 1.35607
R1561 VDD.n1617 VDD.n307 1.35607
R1562 VDD.n1608 VDD.n1607 1.35607
R1563 VDD.n1583 VDD.n331 1.35607
R1564 VDD.n448 VDD.n446 1.35607
R1565 VDD.n1488 VDD.n451 1.35607
R1566 VDD.n1479 VDD.n1478 1.35607
R1567 VDD.n1454 VDD.n484 1.35607
R1568 VDD.n1445 VDD.n1444 1.35607
R1569 VDD.n1420 VDD.n508 1.35607
R1570 VDD.n625 VDD.n623 1.35607
R1571 VDD.n1325 VDD.n628 1.35607
R1572 VDD.n1316 VDD.n1315 1.35607
R1573 VDD.n1291 VDD.n661 1.35607
R1574 VDD.n1282 VDD.n1281 1.35607
R1575 VDD.n1257 VDD.n685 1.35607
R1576 VDD.n802 VDD.n800 1.35607
R1577 VDD.n1162 VDD.n805 1.35607
R1578 VDD.n1153 VDD.n1152 1.35607
R1579 VDD.n1128 VDD.n838 1.35607
R1580 VDD.n1119 VDD.n1118 1.35607
R1581 VDD.n1094 VDD.n863 1.35607
R1582 VDD.n1197 VDD.n1196 1.35607
R1583 VDD.n1209 VDD.n1208 1.35607
R1584 VDD.n1221 VDD.n1220 1.35607
R1585 VDD.n1233 VDD.n1232 1.35607
R1586 VDD.n1183 VDD.n1182 1.35607
R1587 VDD.n1245 VDD.n1244 1.35607
R1588 VDD.n1360 VDD.n1359 1.35607
R1589 VDD.n1372 VDD.n1371 1.35607
R1590 VDD.n1384 VDD.n1383 1.35607
R1591 VDD.n1396 VDD.n1395 1.35607
R1592 VDD.n1346 VDD.n1345 1.35607
R1593 VDD.n1408 VDD.n1407 1.35607
R1594 VDD.n1523 VDD.n1522 1.35607
R1595 VDD.n1535 VDD.n1534 1.35607
R1596 VDD.n1547 VDD.n1546 1.35607
R1597 VDD.n1559 VDD.n1558 1.35607
R1598 VDD.n1509 VDD.n1508 1.35607
R1599 VDD.n1571 VDD.n1570 1.35607
R1600 VDD.n1685 VDD.n232 1.35607
R1601 VDD.n168 VDD.n167 1.35607
R1602 VDD.n1703 VDD.n164 1.35607
R1603 VDD.n1672 VDD.n1671 1.35607
R1604 VDD.n1709 VDD.n79 1.35607
R1605 VDD.n1043 VDD.n945 1.35607
R1606 VDD.n1055 VDD.n1054 1.35607
R1607 VDD.n1064 VDD.n906 1.35607
R1608 VDD.n1076 VDD.n1075 1.35607
R1609 VDD.n1757 VDD.n1756 1.35607
R1610 VDD.n51 VDD.n39 1.13981
R1611 VDD.n1092 VDD.n1091 1.13717
R1612 VDD.n78 VDD.n77 1.13717
R1613 VDD.n867 VDD.n865 1.13717
R1614 VDD.n868 VDD.n854 1.13717
R1615 VDD.n870 VDD.n856 1.13717
R1616 VDD.n1126 VDD.n1125 1.13717
R1617 VDD.n842 VDD.n840 1.13717
R1618 VDD.n843 VDD.n830 1.13717
R1619 VDD.n845 VDD.n832 1.13717
R1620 VDD.n1160 VDD.n1159 1.13717
R1621 VDD.n809 VDD.n807 1.13717
R1622 VDD.n818 VDD.n817 1.13717
R1623 VDD.n820 VDD.n819 1.13717
R1624 VDD.n741 VDD.n725 1.13717
R1625 VDD.n1235 VDD.n1234 1.13717
R1626 VDD.n757 VDD.n740 1.13717
R1627 VDD.n1223 VDD.n1222 1.13717
R1628 VDD.n773 VDD.n756 1.13717
R1629 VDD.n1211 VDD.n1210 1.13717
R1630 VDD.n787 VDD.n772 1.13717
R1631 VDD.n1199 VDD.n1198 1.13717
R1632 VDD.n812 VDD.n786 1.13717
R1633 VDD.n1185 VDD.n1184 1.13717
R1634 VDD.n702 VDD.n701 1.13717
R1635 VDD.n1247 VDD.n1246 1.13717
R1636 VDD.n1255 VDD.n1254 1.13717
R1637 VDD.n689 VDD.n687 1.13717
R1638 VDD.n690 VDD.n677 1.13717
R1639 VDD.n692 VDD.n679 1.13717
R1640 VDD.n1289 VDD.n1288 1.13717
R1641 VDD.n665 VDD.n663 1.13717
R1642 VDD.n666 VDD.n653 1.13717
R1643 VDD.n668 VDD.n655 1.13717
R1644 VDD.n1323 VDD.n1322 1.13717
R1645 VDD.n632 VDD.n630 1.13717
R1646 VDD.n641 VDD.n640 1.13717
R1647 VDD.n643 VDD.n642 1.13717
R1648 VDD.n564 VDD.n548 1.13717
R1649 VDD.n1398 VDD.n1397 1.13717
R1650 VDD.n580 VDD.n563 1.13717
R1651 VDD.n1386 VDD.n1385 1.13717
R1652 VDD.n596 VDD.n579 1.13717
R1653 VDD.n1374 VDD.n1373 1.13717
R1654 VDD.n610 VDD.n595 1.13717
R1655 VDD.n1362 VDD.n1361 1.13717
R1656 VDD.n635 VDD.n609 1.13717
R1657 VDD.n1348 VDD.n1347 1.13717
R1658 VDD.n525 VDD.n524 1.13717
R1659 VDD.n1410 VDD.n1409 1.13717
R1660 VDD.n1418 VDD.n1417 1.13717
R1661 VDD.n512 VDD.n510 1.13717
R1662 VDD.n513 VDD.n500 1.13717
R1663 VDD.n515 VDD.n502 1.13717
R1664 VDD.n1452 VDD.n1451 1.13717
R1665 VDD.n488 VDD.n486 1.13717
R1666 VDD.n489 VDD.n476 1.13717
R1667 VDD.n491 VDD.n478 1.13717
R1668 VDD.n1486 VDD.n1485 1.13717
R1669 VDD.n455 VDD.n453 1.13717
R1670 VDD.n464 VDD.n463 1.13717
R1671 VDD.n466 VDD.n465 1.13717
R1672 VDD.n387 VDD.n371 1.13717
R1673 VDD.n1561 VDD.n1560 1.13717
R1674 VDD.n403 VDD.n386 1.13717
R1675 VDD.n1549 VDD.n1548 1.13717
R1676 VDD.n419 VDD.n402 1.13717
R1677 VDD.n1537 VDD.n1536 1.13717
R1678 VDD.n433 VDD.n418 1.13717
R1679 VDD.n1525 VDD.n1524 1.13717
R1680 VDD.n458 VDD.n432 1.13717
R1681 VDD.n1511 VDD.n1510 1.13717
R1682 VDD.n348 VDD.n347 1.13717
R1683 VDD.n1573 VDD.n1572 1.13717
R1684 VDD.n1581 VDD.n1580 1.13717
R1685 VDD.n335 VDD.n333 1.13717
R1686 VDD.n336 VDD.n323 1.13717
R1687 VDD.n338 VDD.n325 1.13717
R1688 VDD.n1615 VDD.n1614 1.13717
R1689 VDD.n311 VDD.n309 1.13717
R1690 VDD.n312 VDD.n299 1.13717
R1691 VDD.n314 VDD.n301 1.13717
R1692 VDD.n1649 VDD.n1648 1.13717
R1693 VDD.n278 VDD.n276 1.13717
R1694 VDD.n287 VDD.n286 1.13717
R1695 VDD.n289 VDD.n288 1.13717
R1696 VDD.n221 VDD.n220 1.13717
R1697 VDD.n213 VDD.n172 1.13717
R1698 VDD.n1693 VDD.n170 1.13717
R1699 VDD.n1696 VDD.n1695 1.13717
R1700 VDD.n255 VDD.n254 1.13717
R1701 VDD.n230 VDD.n228 1.13717
R1702 VDD.n281 VDD.n252 1.13717
R1703 VDD.n1674 VDD.n1673 1.13717
R1704 VDD.n182 VDD.n181 1.13717
R1705 VDD.n201 VDD.n200 1.13717
R1706 VDD.n185 VDD.n184 1.13717
R1707 VDD.n975 VDD.n961 1.13717
R1708 VDD.n878 VDD.n877 1.13717
R1709 VDD.n911 VDD.n883 1.13717
R1710 VDD.n1062 VDD.n1061 1.13717
R1711 VDD.n950 VDD.n922 1.13717
R1712 VDD.n1041 VDD.n1040 1.13717
R1713 VDD.n949 VDD.n947 1.13717
R1714 VDD.n952 VDD.n924 1.13717
R1715 VDD.n910 VDD.n908 1.13717
R1716 VDD.n913 VDD.n885 1.13717
R1717 VDD.n1083 VDD.n1082 1.13717
R1718 VDD.n976 VDD.n963 1.13717
R1719 VDD.n1755 VDD.n12 1.13717
R1720 VDD.n73 VDD.n72 1.13462
R1721 VDD.n69 VDD.n68 1.13462
R1722 VDD.n65 VDD.n64 1.13462
R1723 VDD.n58 VDD.n57 1.13462
R1724 VDD.n1725 VDD.n38 1.13462
R1725 VDD.n48 VDD.n47 1.13005
R1726 VDD.n1730 VDD.n1729 1.04017
R1727 VDD.n62 VDD.n61 1.04017
R1728 VDD.n999 VDD.n998 1.04017
R1729 VDD.n996 VDD.n995 1.04017
R1730 VDD.n992 VDD.n991 1.04017
R1731 VDD.n30 VDD.t8 1.03618
R1732 VDD.n1759 VDD.n5 0.985115
R1733 VDD.t3 VDD 0.918966
R1734 VDD.n25 VDD.n23 0.870766
R1735 VDD.n20 VDD.n18 0.870578
R1736 VDD.n41 VDD.n40 0.853291
R1737 VDD.n1714 VDD.n74 0.853
R1738 VDD.n1717 VDD.n70 0.853
R1739 VDD.n1720 VDD.n66 0.853
R1740 VDD.n1723 VDD.n59 0.853
R1741 VDD.n1728 VDD.n1727 0.853
R1742 VDD.n983 VDD.n982 0.853
R1743 VDD.n1756 VDD.n1755 0.853
R1744 VDD.n1084 VDD.n879 0.849366
R1745 VDD.n1743 VDD.n28 0.788192
R1746 VDD.n1761 VDD.n1759 0.788192
R1747 VDD.n1740 VDD 0.765888
R1748 VDD.n52 VDD.n51 0.684595
R1749 VDD.n19 VDD.n14 0.682713
R1750 VDD.n1750 VDD.n1749 0.682713
R1751 VDD.n985 VDD.n984 0.682447
R1752 VDD.n1010 VDD.t13 0.612811
R1753 VDD.n1706 VDD.n118 0.459733
R1754 VDD.n1739 VDD.t10 0.459733
R1755 VDD.t8 VDD.t16 0.459733
R1756 VDD.n1768 VDD.n1767 0.394346
R1757 VDD.n50 VDD.n49 0.357419
R1758 VDD.n356 VDD.n355 0.314894
R1759 VDD.n533 VDD.n532 0.314894
R1760 VDD.n710 VDD.n709 0.314894
R1761 VDD.n31 VDD.t16 0.309574
R1762 VDD.n1666 VDD.n268 0.30353
R1763 VDD.n1503 VDD.n445 0.30353
R1764 VDD.n1340 VDD.n622 0.30353
R1765 VDD.n1177 VDD.n799 0.30353
R1766 VDD.n1665 VDD.n1664 0.30353
R1767 VDD.n1502 VDD.n1501 0.30353
R1768 VDD.n1339 VDD.n1338 0.30353
R1769 VDD.n1176 VDD.n1175 0.30353
R1770 VDD.n353 VDD.n352 0.288379
R1771 VDD.n530 VDD.n529 0.288379
R1772 VDD.n707 VDD.n706 0.288379
R1773 VDD.n1708 VDD.n81 0.194439
R1774 VDD.n205 VDD.n179 0.194439
R1775 VDD.n205 VDD.n177 0.194439
R1776 VDD.n1704 VDD.n161 0.194439
R1777 VDD.n1704 VDD.n162 0.194439
R1778 VDD.n238 VDD.n237 0.194439
R1779 VDD.n239 VDD.n238 0.194439
R1780 VDD.n1684 VDD.n246 0.194439
R1781 VDD.n1684 VDD.n1681 0.194439
R1782 VDD.n1670 VDD.n266 0.194439
R1783 VDD.n1670 VDD.n1669 0.194439
R1784 VDD.n1661 VDD.n1660 0.194439
R1785 VDD.n1660 VDD.n1659 0.194439
R1786 VDD.n1626 VDD.n272 0.194439
R1787 VDD.n1629 VDD.n1626 0.194439
R1788 VDD.n1640 VDD.n304 0.194439
R1789 VDD.n1640 VDD.n1625 0.194439
R1790 VDD.n1592 VDD.n305 0.194439
R1791 VDD.n1595 VDD.n1592 0.194439
R1792 VDD.n1606 VDD.n328 0.194439
R1793 VDD.n1606 VDD.n1591 0.194439
R1794 VDD.n358 VDD.n329 0.194439
R1795 VDD.n361 VDD.n358 0.194439
R1796 VDD.n1569 VDD.n365 0.194439
R1797 VDD.n1569 VDD.n1568 0.194439
R1798 VDD.n1557 VDD.n380 0.194439
R1799 VDD.n1557 VDD.n1556 0.194439
R1800 VDD.n1545 VDD.n396 0.194439
R1801 VDD.n1545 VDD.n1544 0.194439
R1802 VDD.n1533 VDD.n412 0.194439
R1803 VDD.n1533 VDD.n1532 0.194439
R1804 VDD.n1521 VDD.n427 0.194439
R1805 VDD.n1521 VDD.n1518 0.194439
R1806 VDD.n1507 VDD.n443 0.194439
R1807 VDD.n1507 VDD.n1506 0.194439
R1808 VDD.n1498 VDD.n1497 0.194439
R1809 VDD.n1497 VDD.n1496 0.194439
R1810 VDD.n1463 VDD.n449 0.194439
R1811 VDD.n1466 VDD.n1463 0.194439
R1812 VDD.n1477 VDD.n481 0.194439
R1813 VDD.n1477 VDD.n1462 0.194439
R1814 VDD.n1429 VDD.n482 0.194439
R1815 VDD.n1432 VDD.n1429 0.194439
R1816 VDD.n1443 VDD.n505 0.194439
R1817 VDD.n1443 VDD.n1428 0.194439
R1818 VDD.n535 VDD.n506 0.194439
R1819 VDD.n538 VDD.n535 0.194439
R1820 VDD.n1406 VDD.n542 0.194439
R1821 VDD.n1406 VDD.n1405 0.194439
R1822 VDD.n1394 VDD.n557 0.194439
R1823 VDD.n1394 VDD.n1393 0.194439
R1824 VDD.n1382 VDD.n573 0.194439
R1825 VDD.n1382 VDD.n1381 0.194439
R1826 VDD.n1370 VDD.n589 0.194439
R1827 VDD.n1370 VDD.n1369 0.194439
R1828 VDD.n1358 VDD.n604 0.194439
R1829 VDD.n1358 VDD.n1355 0.194439
R1830 VDD.n1344 VDD.n620 0.194439
R1831 VDD.n1344 VDD.n1343 0.194439
R1832 VDD.n1335 VDD.n1334 0.194439
R1833 VDD.n1334 VDD.n1333 0.194439
R1834 VDD.n1300 VDD.n626 0.194439
R1835 VDD.n1303 VDD.n1300 0.194439
R1836 VDD.n1314 VDD.n658 0.194439
R1837 VDD.n1314 VDD.n1299 0.194439
R1838 VDD.n1266 VDD.n659 0.194439
R1839 VDD.n1269 VDD.n1266 0.194439
R1840 VDD.n1280 VDD.n682 0.194439
R1841 VDD.n1280 VDD.n1265 0.194439
R1842 VDD.n712 VDD.n683 0.194439
R1843 VDD.n715 VDD.n712 0.194439
R1844 VDD.n1243 VDD.n719 0.194439
R1845 VDD.n1243 VDD.n1242 0.194439
R1846 VDD.n1231 VDD.n734 0.194439
R1847 VDD.n1231 VDD.n1230 0.194439
R1848 VDD.n1219 VDD.n750 0.194439
R1849 VDD.n1219 VDD.n1218 0.194439
R1850 VDD.n1207 VDD.n766 0.194439
R1851 VDD.n1207 VDD.n1206 0.194439
R1852 VDD.n1195 VDD.n781 0.194439
R1853 VDD.n1195 VDD.n1192 0.194439
R1854 VDD.n1181 VDD.n797 0.194439
R1855 VDD.n1181 VDD.n1180 0.194439
R1856 VDD.n1172 VDD.n1171 0.194439
R1857 VDD.n1171 VDD.n1170 0.194439
R1858 VDD.n1137 VDD.n803 0.194439
R1859 VDD.n1140 VDD.n1137 0.194439
R1860 VDD.n1151 VDD.n835 0.194439
R1861 VDD.n1151 VDD.n1136 0.194439
R1862 VDD.n1103 VDD.n836 0.194439
R1863 VDD.n1106 VDD.n1103 0.194439
R1864 VDD.n1117 VDD.n859 0.194439
R1865 VDD.n1117 VDD.n1102 0.194439
R1866 VDD.n862 VDD.n860 0.194439
R1867 VDD.n894 VDD.n891 0.194439
R1868 VDD.n1074 VDD.n888 0.194439
R1869 VDD.n1074 VDD.n889 0.194439
R1870 VDD.n931 VDD.n904 0.194439
R1871 VDD.n932 VDD.n931 0.194439
R1872 VDD.n1053 VDD.n927 0.194439
R1873 VDD.n1053 VDD.n928 0.194439
R1874 VDD.n1019 VDD.n943 0.194439
R1875 VDD.n1020 VDD.n1019 0.194439
R1876 VDD.n1032 VDD.n966 0.194439
R1877 VDD.n1032 VDD.n967 0.194439
R1878 VDD.t2 VDD.n31 0.150466
R1879 VDD.n987 VDD.n986 0.132407
R1880 VDD.n986 VDD.n965 0.127283
R1881 VDD.n1713 VDD 0.103754
R1882 VDD.n284 VDD.n283 0.102103
R1883 VDD.n461 VDD.n460 0.102103
R1884 VDD.n638 VDD.n637 0.102103
R1885 VDD.n815 VDD.n814 0.102103
R1886 VDD.n1577 VDD.n1576 0.100721
R1887 VDD.n1414 VDD.n1413 0.100721
R1888 VDD.n1251 VDD.n1250 0.100721
R1889 VDD VDD.n1086 0.100533
R1890 VDD.n1747 VDD.n27 0.0981562
R1891 VDD.n285 VDD.n282 0.0890769
R1892 VDD.n462 VDD.n459 0.0890769
R1893 VDD.n639 VDD.n636 0.0890769
R1894 VDD.n816 VDD.n813 0.0890769
R1895 VDD.n1150 VDD.n122 0.0847059
R1896 VDD.n1116 VDD.n120 0.0847059
R1897 VDD.n1313 VDD.n133 0.0847059
R1898 VDD.n1279 VDD.n131 0.0847059
R1899 VDD.n1476 VDD.n144 0.0847059
R1900 VDD.n1442 VDD.n142 0.0847059
R1901 VDD.n1639 VDD.n155 0.0847059
R1902 VDD.n1605 VDD.n153 0.0847059
R1903 VDD.n206 VDD.n83 0.0847059
R1904 VDD.n1073 VDD.n1072 0.0847059
R1905 VDD.n929 VDD.n903 0.0847059
R1906 VDD.n1052 VDD.n1051 0.0847059
R1907 VDD.n1017 VDD.n942 0.0847059
R1908 VDD.n973 VDD.n968 0.0796667
R1909 VDD.n898 VDD.n895 0.0705758
R1910 VDD.n905 VDD.n887 0.0705758
R1911 VDD.n937 VDD.n933 0.0705758
R1912 VDD.n944 VDD.n926 0.0705758
R1913 VDD.n1025 VDD.n1021 0.0705758
R1914 VDD.n192 VDD.n180 0.0705758
R1915 VDD.n211 VDD.n163 0.0705758
R1916 VDD.n1699 VDD.n1698 0.0705758
R1917 VDD.n1686 VDD.n231 0.0705758
R1918 VDD.n1678 VDD.n248 0.0705758
R1919 VDD.n290 VDD.n273 0.0705758
R1920 VDD.n1634 VDD.n1630 0.0705758
R1921 VDD.n306 VDD.n303 0.0705758
R1922 VDD.n1600 VDD.n1596 0.0705758
R1923 VDD.n330 VDD.n327 0.0705758
R1924 VDD.n1565 VDD.n368 0.0705758
R1925 VDD.n1553 VDD.n383 0.0705758
R1926 VDD.n1541 VDD.n399 0.0705758
R1927 VDD.n1529 VDD.n415 0.0705758
R1928 VDD.n1515 VDD.n429 0.0705758
R1929 VDD.n467 VDD.n450 0.0705758
R1930 VDD.n1471 VDD.n1467 0.0705758
R1931 VDD.n483 VDD.n480 0.0705758
R1932 VDD.n1437 VDD.n1433 0.0705758
R1933 VDD.n507 VDD.n504 0.0705758
R1934 VDD.n1402 VDD.n545 0.0705758
R1935 VDD.n1390 VDD.n560 0.0705758
R1936 VDD.n1378 VDD.n576 0.0705758
R1937 VDD.n1366 VDD.n592 0.0705758
R1938 VDD.n1352 VDD.n606 0.0705758
R1939 VDD.n644 VDD.n627 0.0705758
R1940 VDD.n1308 VDD.n1304 0.0705758
R1941 VDD.n660 VDD.n657 0.0705758
R1942 VDD.n1274 VDD.n1270 0.0705758
R1943 VDD.n684 VDD.n681 0.0705758
R1944 VDD.n1239 VDD.n722 0.0705758
R1945 VDD.n1227 VDD.n737 0.0705758
R1946 VDD.n1215 VDD.n753 0.0705758
R1947 VDD.n1203 VDD.n769 0.0705758
R1948 VDD.n1189 VDD.n783 0.0705758
R1949 VDD.n821 VDD.n804 0.0705758
R1950 VDD.n1145 VDD.n1141 0.0705758
R1951 VDD.n837 VDD.n834 0.0705758
R1952 VDD.n1111 VDD.n1107 0.0705758
R1953 VDD.n861 VDD.n858 0.0705758
R1954 VDD.n1578 VDD 0.0619615
R1955 VDD.n1415 VDD 0.0619615
R1956 VDD.n1252 VDD 0.0619615
R1957 VDD.n1089 VDD 0.0619615
R1958 VDD.n7 VDD.n0 0.0616979
R1959 VDD VDD.n7 0.0603958
R1960 VDD.n1769 VDD.n0 0.0590938
R1961 VDD.n971 VDD 0.0579444
R1962 VDD.n1748 VDD.n1747 0.0577917
R1963 VDD.n195 VDD.n193 0.0573182
R1964 VDD.n215 VDD.n212 0.0573182
R1965 VDD.n1700 VDD.n166 0.0573182
R1966 VDD.n1688 VDD.n229 0.0573182
R1967 VDD.n1677 VDD.n1676 0.0573182
R1968 VDD.n292 VDD.n275 0.0573182
R1969 VDD.n1633 VDD.n1632 0.0573182
R1970 VDD.n316 VDD.n308 0.0573182
R1971 VDD.n1599 VDD.n1598 0.0573182
R1972 VDD.n340 VDD.n332 0.0573182
R1973 VDD.n1564 VDD.n1563 0.0573182
R1974 VDD.n1552 VDD.n1551 0.0573182
R1975 VDD.n1540 VDD.n1539 0.0573182
R1976 VDD.n1528 VDD.n1527 0.0573182
R1977 VDD.n1514 VDD.n1513 0.0573182
R1978 VDD.n469 VDD.n452 0.0573182
R1979 VDD.n1470 VDD.n1469 0.0573182
R1980 VDD.n493 VDD.n485 0.0573182
R1981 VDD.n1436 VDD.n1435 0.0573182
R1982 VDD.n517 VDD.n509 0.0573182
R1983 VDD.n1401 VDD.n1400 0.0573182
R1984 VDD.n1389 VDD.n1388 0.0573182
R1985 VDD.n1377 VDD.n1376 0.0573182
R1986 VDD.n1365 VDD.n1364 0.0573182
R1987 VDD.n1351 VDD.n1350 0.0573182
R1988 VDD.n646 VDD.n629 0.0573182
R1989 VDD.n1307 VDD.n1306 0.0573182
R1990 VDD.n670 VDD.n662 0.0573182
R1991 VDD.n1273 VDD.n1272 0.0573182
R1992 VDD.n694 VDD.n686 0.0573182
R1993 VDD.n1238 VDD.n1237 0.0573182
R1994 VDD.n1226 VDD.n1225 0.0573182
R1995 VDD.n1214 VDD.n1213 0.0573182
R1996 VDD.n1202 VDD.n1201 0.0573182
R1997 VDD.n1188 VDD.n1187 0.0573182
R1998 VDD.n823 VDD.n806 0.0573182
R1999 VDD.n1144 VDD.n1143 0.0573182
R2000 VDD.n847 VDD.n839 0.0573182
R2001 VDD.n1110 VDD.n1109 0.0573182
R2002 VDD.n872 VDD.n864 0.0573182
R2003 VDD.n897 VDD.n896 0.0573182
R2004 VDD.n915 VDD.n907 0.0573182
R2005 VDD.n936 VDD.n935 0.0573182
R2006 VDD.n954 VDD.n946 0.0573182
R2007 VDD.n1024 VDD.n1023 0.0573182
R2008 VDD.n1753 VDD.n23 0.0517727
R2009 VDD.n985 VDD.n968 0.0455
R2010 VDD.n18 VDD.n15 0.0438377
R2011 VDD.n895 VDD.n879 0.0429036
R2012 VDD.n1752 VDD.n1751 0.041625
R2013 VDD.n1748 VDD 0.0408646
R2014 VDD.n1075 VDD.n887 0.0402727
R2015 VDD.n933 VDD.n906 0.0402727
R2016 VDD.n1054 VDD.n926 0.0402727
R2017 VDD.n1021 VDD.n945 0.0402727
R2018 VDD.n1033 VDD.n965 0.0402727
R2019 VDD.n204 VDD.n180 0.0402727
R2020 VDD.n1703 VDD.n163 0.0402727
R2021 VDD.n1698 VDD.n167 0.0402727
R2022 VDD.n1686 VDD.n1685 0.0402727
R2023 VDD.n1671 VDD.n248 0.0402727
R2024 VDD.n290 VDD.n271 0.0402727
R2025 VDD.n1630 VDD.n274 0.0402727
R2026 VDD.n1641 VDD.n303 0.0402727
R2027 VDD.n1596 VDD.n307 0.0402727
R2028 VDD.n1607 VDD.n327 0.0402727
R2029 VDD.n355 VDD.n331 0.0402727
R2030 VDD.n1570 VDD.n356 0.0402727
R2031 VDD.n1558 VDD.n368 0.0402727
R2032 VDD.n1546 VDD.n383 0.0402727
R2033 VDD.n1534 VDD.n399 0.0402727
R2034 VDD.n1522 VDD.n415 0.0402727
R2035 VDD.n1508 VDD.n429 0.0402727
R2036 VDD.n467 VDD.n448 0.0402727
R2037 VDD.n1467 VDD.n451 0.0402727
R2038 VDD.n1478 VDD.n480 0.0402727
R2039 VDD.n1433 VDD.n484 0.0402727
R2040 VDD.n1444 VDD.n504 0.0402727
R2041 VDD.n532 VDD.n508 0.0402727
R2042 VDD.n1407 VDD.n533 0.0402727
R2043 VDD.n1395 VDD.n545 0.0402727
R2044 VDD.n1383 VDD.n560 0.0402727
R2045 VDD.n1371 VDD.n576 0.0402727
R2046 VDD.n1359 VDD.n592 0.0402727
R2047 VDD.n1345 VDD.n606 0.0402727
R2048 VDD.n644 VDD.n625 0.0402727
R2049 VDD.n1304 VDD.n628 0.0402727
R2050 VDD.n1315 VDD.n657 0.0402727
R2051 VDD.n1270 VDD.n661 0.0402727
R2052 VDD.n1281 VDD.n681 0.0402727
R2053 VDD.n709 VDD.n685 0.0402727
R2054 VDD.n1244 VDD.n710 0.0402727
R2055 VDD.n1232 VDD.n722 0.0402727
R2056 VDD.n1220 VDD.n737 0.0402727
R2057 VDD.n1208 VDD.n753 0.0402727
R2058 VDD.n1196 VDD.n769 0.0402727
R2059 VDD.n1182 VDD.n783 0.0402727
R2060 VDD.n821 VDD.n802 0.0402727
R2061 VDD.n1141 VDD.n805 0.0402727
R2062 VDD.n1152 VDD.n834 0.0402727
R2063 VDD.n1107 VDD.n838 0.0402727
R2064 VDD.n1118 VDD.n858 0.0402727
R2065 VDD.n193 VDD.n188 0.0402727
R2066 VDD.n212 VDD.n175 0.0402727
R2067 VDD.n1701 VDD.n1700 0.0402727
R2068 VDD.n240 VDD.n229 0.0402727
R2069 VDD.n1677 VDD.n249 0.0402727
R2070 VDD.n1665 VDD.n261 0.0402727
R2071 VDD.n1664 VDD.n1663 0.0402727
R2072 VDD.n1652 VDD.n275 0.0402727
R2073 VDD.n1633 VDD.n300 0.0402727
R2074 VDD.n1618 VDD.n308 0.0402727
R2075 VDD.n1599 VDD.n324 0.0402727
R2076 VDD.n1584 VDD.n332 0.0402727
R2077 VDD.n1564 VDD.n350 0.0402727
R2078 VDD.n1552 VDD.n376 0.0402727
R2079 VDD.n1540 VDD.n392 0.0402727
R2080 VDD.n1528 VDD.n408 0.0402727
R2081 VDD.n1514 VDD.n424 0.0402727
R2082 VDD.n1502 VDD.n438 0.0402727
R2083 VDD.n1501 VDD.n1500 0.0402727
R2084 VDD.n1489 VDD.n452 0.0402727
R2085 VDD.n1470 VDD.n477 0.0402727
R2086 VDD.n1455 VDD.n485 0.0402727
R2087 VDD.n1436 VDD.n501 0.0402727
R2088 VDD.n1421 VDD.n509 0.0402727
R2089 VDD.n1401 VDD.n527 0.0402727
R2090 VDD.n1389 VDD.n553 0.0402727
R2091 VDD.n1377 VDD.n569 0.0402727
R2092 VDD.n1365 VDD.n585 0.0402727
R2093 VDD.n1351 VDD.n601 0.0402727
R2094 VDD.n1339 VDD.n615 0.0402727
R2095 VDD.n1338 VDD.n1337 0.0402727
R2096 VDD.n1326 VDD.n629 0.0402727
R2097 VDD.n1307 VDD.n654 0.0402727
R2098 VDD.n1292 VDD.n662 0.0402727
R2099 VDD.n1273 VDD.n678 0.0402727
R2100 VDD.n1258 VDD.n686 0.0402727
R2101 VDD.n1238 VDD.n704 0.0402727
R2102 VDD.n1226 VDD.n730 0.0402727
R2103 VDD.n1214 VDD.n746 0.0402727
R2104 VDD.n1202 VDD.n762 0.0402727
R2105 VDD.n1188 VDD.n778 0.0402727
R2106 VDD.n1176 VDD.n792 0.0402727
R2107 VDD.n1175 VDD.n1174 0.0402727
R2108 VDD.n1163 VDD.n806 0.0402727
R2109 VDD.n1144 VDD.n831 0.0402727
R2110 VDD.n1129 VDD.n839 0.0402727
R2111 VDD.n1110 VDD.n855 0.0402727
R2112 VDD.n1095 VDD.n864 0.0402727
R2113 VDD.n897 VDD.n884 0.0402727
R2114 VDD.n1065 VDD.n907 0.0402727
R2115 VDD.n936 VDD.n923 0.0402727
R2116 VDD.n1044 VDD.n946 0.0402727
R2117 VDD.n1024 VDD.n962 0.0402727
R2118 VDD.n1710 VDD.n78 0.0364848
R2119 VDD.n194 VDD.n181 0.0364848
R2120 VDD.n214 VDD.n213 0.0364848
R2121 VDD.n1697 VDD.n1696 0.0364848
R2122 VDD.n1687 VDD.n230 0.0364848
R2123 VDD.n1673 VDD.n250 0.0364848
R2124 VDD.n291 VDD.n289 0.0364848
R2125 VDD.n1631 VDD.n276 0.0364848
R2126 VDD.n315 VDD.n301 0.0364848
R2127 VDD.n1597 VDD.n309 0.0364848
R2128 VDD.n339 VDD.n325 0.0364848
R2129 VDD.n354 VDD.n333 0.0364848
R2130 VDD.n1572 VDD.n349 0.0364848
R2131 VDD.n1560 VDD.n369 0.0364848
R2132 VDD.n1548 VDD.n384 0.0364848
R2133 VDD.n1536 VDD.n400 0.0364848
R2134 VDD.n1524 VDD.n416 0.0364848
R2135 VDD.n1510 VDD.n430 0.0364848
R2136 VDD.n468 VDD.n466 0.0364848
R2137 VDD.n1468 VDD.n453 0.0364848
R2138 VDD.n492 VDD.n478 0.0364848
R2139 VDD.n1434 VDD.n486 0.0364848
R2140 VDD.n516 VDD.n502 0.0364848
R2141 VDD.n531 VDD.n510 0.0364848
R2142 VDD.n1409 VDD.n526 0.0364848
R2143 VDD.n1397 VDD.n546 0.0364848
R2144 VDD.n1385 VDD.n561 0.0364848
R2145 VDD.n1373 VDD.n577 0.0364848
R2146 VDD.n1361 VDD.n593 0.0364848
R2147 VDD.n1347 VDD.n607 0.0364848
R2148 VDD.n645 VDD.n643 0.0364848
R2149 VDD.n1305 VDD.n630 0.0364848
R2150 VDD.n669 VDD.n655 0.0364848
R2151 VDD.n1271 VDD.n663 0.0364848
R2152 VDD.n693 VDD.n679 0.0364848
R2153 VDD.n708 VDD.n687 0.0364848
R2154 VDD.n1246 VDD.n703 0.0364848
R2155 VDD.n1234 VDD.n723 0.0364848
R2156 VDD.n1222 VDD.n738 0.0364848
R2157 VDD.n1210 VDD.n754 0.0364848
R2158 VDD.n1198 VDD.n770 0.0364848
R2159 VDD.n1184 VDD.n784 0.0364848
R2160 VDD.n822 VDD.n820 0.0364848
R2161 VDD.n1142 VDD.n807 0.0364848
R2162 VDD.n846 VDD.n832 0.0364848
R2163 VDD.n1108 VDD.n840 0.0364848
R2164 VDD.n871 VDD.n856 0.0364848
R2165 VDD.n1087 VDD.n865 0.0364848
R2166 VDD.n1083 VDD.n880 0.0364848
R2167 VDD.n914 VDD.n885 0.0364848
R2168 VDD.n934 VDD.n908 0.0364848
R2169 VDD.n953 VDD.n924 0.0364848
R2170 VDD.n1022 VDD.n947 0.0364848
R2171 VDD.n972 VDD.n963 0.0364848
R2172 VDD.n17 VDD.n16 0.0351948
R2173 VDD.n1756 VDD.n10 0.0309054
R2174 VDD.n899 VDD.n886 0.030803
R2175 VDD.n1067 VDD.n1066 0.030803
R2176 VDD.n938 VDD.n925 0.030803
R2177 VDD.n1046 VDD.n1045 0.030803
R2178 VDD.n1026 VDD.n964 0.030803
R2179 VDD.n191 VDD.n80 0.030803
R2180 VDD.n210 VDD.n176 0.030803
R2181 VDD.n1702 VDD.n165 0.030803
R2182 VDD.n242 VDD.n241 0.030803
R2183 VDD.n1679 VDD.n233 0.030803
R2184 VDD.n1667 VDD.n263 0.030803
R2185 VDD.n1662 VDD.n270 0.030803
R2186 VDD.n1654 VDD.n1653 0.030803
R2187 VDD.n1635 VDD.n302 0.030803
R2188 VDD.n1620 VDD.n1619 0.030803
R2189 VDD.n1601 VDD.n326 0.030803
R2190 VDD.n1586 VDD.n1585 0.030803
R2191 VDD.n1566 VDD.n357 0.030803
R2192 VDD.n1554 VDD.n378 0.030803
R2193 VDD.n1542 VDD.n394 0.030803
R2194 VDD.n1530 VDD.n410 0.030803
R2195 VDD.n1516 VDD.n426 0.030803
R2196 VDD.n1504 VDD.n440 0.030803
R2197 VDD.n1499 VDD.n447 0.030803
R2198 VDD.n1491 VDD.n1490 0.030803
R2199 VDD.n1472 VDD.n479 0.030803
R2200 VDD.n1457 VDD.n1456 0.030803
R2201 VDD.n1438 VDD.n503 0.030803
R2202 VDD.n1423 VDD.n1422 0.030803
R2203 VDD.n1403 VDD.n534 0.030803
R2204 VDD.n1391 VDD.n555 0.030803
R2205 VDD.n1379 VDD.n571 0.030803
R2206 VDD.n1367 VDD.n587 0.030803
R2207 VDD.n1353 VDD.n603 0.030803
R2208 VDD.n1341 VDD.n617 0.030803
R2209 VDD.n1336 VDD.n624 0.030803
R2210 VDD.n1328 VDD.n1327 0.030803
R2211 VDD.n1309 VDD.n656 0.030803
R2212 VDD.n1294 VDD.n1293 0.030803
R2213 VDD.n1275 VDD.n680 0.030803
R2214 VDD.n1260 VDD.n1259 0.030803
R2215 VDD.n1240 VDD.n711 0.030803
R2216 VDD.n1228 VDD.n732 0.030803
R2217 VDD.n1216 VDD.n748 0.030803
R2218 VDD.n1204 VDD.n764 0.030803
R2219 VDD.n1190 VDD.n780 0.030803
R2220 VDD.n1178 VDD.n794 0.030803
R2221 VDD.n1173 VDD.n801 0.030803
R2222 VDD.n1165 VDD.n1164 0.030803
R2223 VDD.n1146 VDD.n833 0.030803
R2224 VDD.n1131 VDD.n1130 0.030803
R2225 VDD.n1112 VDD.n857 0.030803
R2226 VDD.n1097 VDD.n1096 0.030803
R2227 VDD.n26 VDD.n9 0.0292162
R2228 VDD.n56 VDD.n55 0.0273994
R2229 VDD.n30 VDD 0.0271814
R2230 VDD.n8 VDD 0.0265417
R2231 VDD.n1728 VDD.n36 0.0242893
R2232 VDD.n60 VDD.n59 0.0242893
R2233 VDD.n997 VDD.n66 0.0242893
R2234 VDD.n994 VDD.n70 0.0242893
R2235 VDD.n990 VDD.n74 0.0242893
R2236 VDD.n1757 VDD.n8 0.0239375
R2237 VDD.n46 VDD.n45 0.0234759
R2238 VDD VDD.n1769 0.0226354
R2239 VDD.n980 VDD.n979 0.0206084
R2240 VDD.n187 VDD.n186 0.0205441
R2241 VDD.n202 VDD.n174 0.0205441
R2242 VDD.n223 VDD.n222 0.0205441
R2243 VDD.n1691 VDD.n227 0.0205441
R2244 VDD.n257 VDD.n256 0.0205441
R2245 VDD.n283 VDD.n262 0.0205441
R2246 VDD.n372 VDD.n351 0.0205441
R2247 VDD.n388 VDD.n377 0.0205441
R2248 VDD.n404 VDD.n393 0.0205441
R2249 VDD.n420 VDD.n409 0.0205441
R2250 VDD.n434 VDD.n425 0.0205441
R2251 VDD.n460 VDD.n439 0.0205441
R2252 VDD.n549 VDD.n528 0.0205441
R2253 VDD.n565 VDD.n554 0.0205441
R2254 VDD.n581 VDD.n570 0.0205441
R2255 VDD.n597 VDD.n586 0.0205441
R2256 VDD.n611 VDD.n602 0.0205441
R2257 VDD.n637 VDD.n616 0.0205441
R2258 VDD.n726 VDD.n705 0.0205441
R2259 VDD.n742 VDD.n731 0.0205441
R2260 VDD.n758 VDD.n747 0.0205441
R2261 VDD.n774 VDD.n763 0.0205441
R2262 VDD.n788 VDD.n779 0.0205441
R2263 VDD.n814 VDD.n793 0.0205441
R2264 VDD.n284 VDD.n280 0.0198529
R2265 VDD.n1650 VDD.n277 0.0198529
R2266 VDD.n1644 VDD.n1643 0.0198529
R2267 VDD.n1616 VDD.n310 0.0198529
R2268 VDD.n1610 VDD.n1609 0.0198529
R2269 VDD.n1582 VDD.n334 0.0198529
R2270 VDD.n461 VDD.n457 0.0198529
R2271 VDD.n1487 VDD.n454 0.0198529
R2272 VDD.n1481 VDD.n1480 0.0198529
R2273 VDD.n1453 VDD.n487 0.0198529
R2274 VDD.n1447 VDD.n1446 0.0198529
R2275 VDD.n1419 VDD.n511 0.0198529
R2276 VDD.n638 VDD.n634 0.0198529
R2277 VDD.n1324 VDD.n631 0.0198529
R2278 VDD.n1318 VDD.n1317 0.0198529
R2279 VDD.n1290 VDD.n664 0.0198529
R2280 VDD.n1284 VDD.n1283 0.0198529
R2281 VDD.n1256 VDD.n688 0.0198529
R2282 VDD.n815 VDD.n811 0.0198529
R2283 VDD.n1161 VDD.n808 0.0198529
R2284 VDD.n1155 VDD.n1154 0.0198529
R2285 VDD.n1127 VDD.n841 0.0198529
R2286 VDD.n1121 VDD.n1120 0.0198529
R2287 VDD.n1093 VDD.n866 0.0198529
R2288 VDD.n1078 VDD.n1077 0.0198529
R2289 VDD.n1063 VDD.n909 0.0198529
R2290 VDD.n1057 VDD.n1056 0.0198529
R2291 VDD.n1042 VDD.n948 0.0198529
R2292 VDD.n1036 VDD.n1035 0.0198529
R2293 VDD.n1753 VDD.n12 0.0188117
R2294 VDD.n15 VDD.n12 0.0188117
R2295 VDD.n184 VDD.n183 0.0185769
R2296 VDD.n200 VDD.n173 0.0185769
R2297 VDD.n220 VDD.n171 0.0185769
R2298 VDD.n1693 VDD.n1692 0.0185769
R2299 VDD.n258 VDD.n254 0.0185769
R2300 VDD.n282 VDD.n281 0.0185769
R2301 VDD.n295 VDD.n279 0.0185769
R2302 VDD.n1647 VDD.n1646 0.0185769
R2303 VDD.n319 VDD.n313 0.0185769
R2304 VDD.n1613 VDD.n1612 0.0185769
R2305 VDD.n343 VDD.n337 0.0185769
R2306 VDD.n1579 VDD.n1578 0.0185769
R2307 VDD.n373 VDD.n347 0.0185769
R2308 VDD.n389 VDD.n387 0.0185769
R2309 VDD.n405 VDD.n403 0.0185769
R2310 VDD.n421 VDD.n419 0.0185769
R2311 VDD.n435 VDD.n433 0.0185769
R2312 VDD.n459 VDD.n458 0.0185769
R2313 VDD.n472 VDD.n456 0.0185769
R2314 VDD.n1484 VDD.n1483 0.0185769
R2315 VDD.n496 VDD.n490 0.0185769
R2316 VDD.n1450 VDD.n1449 0.0185769
R2317 VDD.n520 VDD.n514 0.0185769
R2318 VDD.n1416 VDD.n1415 0.0185769
R2319 VDD.n550 VDD.n524 0.0185769
R2320 VDD.n566 VDD.n564 0.0185769
R2321 VDD.n582 VDD.n580 0.0185769
R2322 VDD.n598 VDD.n596 0.0185769
R2323 VDD.n612 VDD.n610 0.0185769
R2324 VDD.n636 VDD.n635 0.0185769
R2325 VDD.n649 VDD.n633 0.0185769
R2326 VDD.n1321 VDD.n1320 0.0185769
R2327 VDD.n673 VDD.n667 0.0185769
R2328 VDD.n1287 VDD.n1286 0.0185769
R2329 VDD.n697 VDD.n691 0.0185769
R2330 VDD.n1253 VDD.n1252 0.0185769
R2331 VDD.n727 VDD.n701 0.0185769
R2332 VDD.n743 VDD.n741 0.0185769
R2333 VDD.n759 VDD.n757 0.0185769
R2334 VDD.n775 VDD.n773 0.0185769
R2335 VDD.n789 VDD.n787 0.0185769
R2336 VDD.n813 VDD.n812 0.0185769
R2337 VDD.n826 VDD.n810 0.0185769
R2338 VDD.n1158 VDD.n1157 0.0185769
R2339 VDD.n850 VDD.n844 0.0185769
R2340 VDD.n1124 VDD.n1123 0.0185769
R2341 VDD.n875 VDD.n869 0.0185769
R2342 VDD.n1090 VDD.n1089 0.0185769
R2343 VDD.n981 VDD.n971 0.0185349
R2344 VDD.n1711 VDD.n77 0.0184706
R2345 VDD.n196 VDD.n182 0.0184706
R2346 VDD.n216 VDD.n172 0.0184706
R2347 VDD.n1695 VDD.n169 0.0184706
R2348 VDD.n1689 VDD.n228 0.0184706
R2349 VDD.n1675 VDD.n1674 0.0184706
R2350 VDD.n293 VDD.n288 0.0184706
R2351 VDD.n298 VDD.n278 0.0184706
R2352 VDD.n317 VDD.n314 0.0184706
R2353 VDD.n322 VDD.n311 0.0184706
R2354 VDD.n341 VDD.n338 0.0184706
R2355 VDD.n345 VDD.n335 0.0184706
R2356 VDD.n1573 VDD.n346 0.0184706
R2357 VDD.n1562 VDD.n1561 0.0184706
R2358 VDD.n1550 VDD.n1549 0.0184706
R2359 VDD.n1538 VDD.n1537 0.0184706
R2360 VDD.n1526 VDD.n1525 0.0184706
R2361 VDD.n1512 VDD.n1511 0.0184706
R2362 VDD.n470 VDD.n465 0.0184706
R2363 VDD.n475 VDD.n455 0.0184706
R2364 VDD.n494 VDD.n491 0.0184706
R2365 VDD.n499 VDD.n488 0.0184706
R2366 VDD.n518 VDD.n515 0.0184706
R2367 VDD.n522 VDD.n512 0.0184706
R2368 VDD.n1410 VDD.n523 0.0184706
R2369 VDD.n1399 VDD.n1398 0.0184706
R2370 VDD.n1387 VDD.n1386 0.0184706
R2371 VDD.n1375 VDD.n1374 0.0184706
R2372 VDD.n1363 VDD.n1362 0.0184706
R2373 VDD.n1349 VDD.n1348 0.0184706
R2374 VDD.n647 VDD.n642 0.0184706
R2375 VDD.n652 VDD.n632 0.0184706
R2376 VDD.n671 VDD.n668 0.0184706
R2377 VDD.n676 VDD.n665 0.0184706
R2378 VDD.n695 VDD.n692 0.0184706
R2379 VDD.n699 VDD.n689 0.0184706
R2380 VDD.n1247 VDD.n700 0.0184706
R2381 VDD.n1236 VDD.n1235 0.0184706
R2382 VDD.n1224 VDD.n1223 0.0184706
R2383 VDD.n1212 VDD.n1211 0.0184706
R2384 VDD.n1200 VDD.n1199 0.0184706
R2385 VDD.n1186 VDD.n1185 0.0184706
R2386 VDD.n824 VDD.n819 0.0184706
R2387 VDD.n829 VDD.n809 0.0184706
R2388 VDD.n848 VDD.n845 0.0184706
R2389 VDD.n853 VDD.n842 0.0184706
R2390 VDD.n873 VDD.n870 0.0184706
R2391 VDD.n1088 VDD.n867 0.0184706
R2392 VDD.n1082 VDD.n881 0.0184706
R2393 VDD.n916 VDD.n913 0.0184706
R2394 VDD.n921 VDD.n910 0.0184706
R2395 VDD.n955 VDD.n952 0.0184706
R2396 VDD.n960 VDD.n949 0.0184706
R2397 VDD.n976 VDD.n974 0.0184706
R2398 VDD.n1712 VDD.n76 0.0179744
R2399 VDD.n199 VDD.n198 0.0179744
R2400 VDD.n219 VDD.n218 0.0179744
R2401 VDD.n1694 VDD.n225 0.0179744
R2402 VDD.n253 VDD.n226 0.0179744
R2403 VDD.n260 VDD.n259 0.0179744
R2404 VDD.n286 VDD.n285 0.0179744
R2405 VDD.n1648 VDD.n296 0.0179744
R2406 VDD.n312 VDD.n297 0.0179744
R2407 VDD.n1614 VDD.n320 0.0179744
R2408 VDD.n336 VDD.n321 0.0179744
R2409 VDD.n1580 VDD.n344 0.0179744
R2410 VDD.n1575 VDD.n1574 0.0179744
R2411 VDD.n375 VDD.n374 0.0179744
R2412 VDD.n391 VDD.n390 0.0179744
R2413 VDD.n407 VDD.n406 0.0179744
R2414 VDD.n423 VDD.n422 0.0179744
R2415 VDD.n437 VDD.n436 0.0179744
R2416 VDD.n463 VDD.n462 0.0179744
R2417 VDD.n1485 VDD.n473 0.0179744
R2418 VDD.n489 VDD.n474 0.0179744
R2419 VDD.n1451 VDD.n497 0.0179744
R2420 VDD.n513 VDD.n498 0.0179744
R2421 VDD.n1417 VDD.n521 0.0179744
R2422 VDD.n1412 VDD.n1411 0.0179744
R2423 VDD.n552 VDD.n551 0.0179744
R2424 VDD.n568 VDD.n567 0.0179744
R2425 VDD.n584 VDD.n583 0.0179744
R2426 VDD.n600 VDD.n599 0.0179744
R2427 VDD.n614 VDD.n613 0.0179744
R2428 VDD.n640 VDD.n639 0.0179744
R2429 VDD.n1322 VDD.n650 0.0179744
R2430 VDD.n666 VDD.n651 0.0179744
R2431 VDD.n1288 VDD.n674 0.0179744
R2432 VDD.n690 VDD.n675 0.0179744
R2433 VDD.n1254 VDD.n698 0.0179744
R2434 VDD.n1249 VDD.n1248 0.0179744
R2435 VDD.n729 VDD.n728 0.0179744
R2436 VDD.n745 VDD.n744 0.0179744
R2437 VDD.n761 VDD.n760 0.0179744
R2438 VDD.n777 VDD.n776 0.0179744
R2439 VDD.n791 VDD.n790 0.0179744
R2440 VDD.n817 VDD.n816 0.0179744
R2441 VDD.n1159 VDD.n827 0.0179744
R2442 VDD.n843 VDD.n828 0.0179744
R2443 VDD.n1125 VDD.n851 0.0179744
R2444 VDD.n868 VDD.n852 0.0179744
R2445 VDD.n1091 VDD.n876 0.0179744
R2446 VDD.n1081 VDD.n1080 0.0179074
R2447 VDD.n918 VDD.n912 0.0179074
R2448 VDD.n1060 VDD.n1059 0.0179074
R2449 VDD.n957 VDD.n951 0.0179074
R2450 VDD.n1039 VDD.n1038 0.0179074
R2451 VDD.n978 VDD.n977 0.0179074
R2452 VDD.n1086 VDD.n877 0.0173272
R2453 VDD.n911 VDD.n882 0.0173272
R2454 VDD.n1061 VDD.n919 0.0173272
R2455 VDD.n950 VDD.n920 0.0173272
R2456 VDD.n1040 VDD.n958 0.0173272
R2457 VDD.n975 VDD.n959 0.0173272
R2458 VDD.n49 VDD.n40 0.0172857
R2459 VDD.n982 VDD.n981 0.0168953
R2460 VDD.n982 VDD.n969 0.0168953
R2461 VDD.n1722 VDD.n1721 0.0167579
R2462 VDD.n1744 VDD.n6 0.016125
R2463 VDD.n54 VDD.n53 0.0156071
R2464 VDD.n1727 VDD.n37 0.0156071
R2465 VDD.n1723 VDD.n63 0.0156071
R2466 VDD.n1720 VDD.n67 0.0156071
R2467 VDD.n1717 VDD.n71 0.0156071
R2468 VDD.n1714 VDD.n75 0.0156071
R2469 VDD.n983 VDD.n970 0.0152558
R2470 VDD.n47 VDD.n44 0.0148621
R2471 VDD.n1726 VDD.n1724 0.0148365
R2472 VDD.n197 VDD.n187 0.0143235
R2473 VDD.n217 VDD.n174 0.0143235
R2474 VDD.n224 VDD.n223 0.0143235
R2475 VDD.n1691 VDD.n1690 0.0143235
R2476 VDD.n257 VDD.n251 0.0143235
R2477 VDD.n294 VDD.n277 0.0143235
R2478 VDD.n1645 VDD.n1644 0.0143235
R2479 VDD.n318 VDD.n310 0.0143235
R2480 VDD.n1611 VDD.n1610 0.0143235
R2481 VDD.n342 VDD.n334 0.0143235
R2482 VDD.n372 VDD.n370 0.0143235
R2483 VDD.n388 VDD.n385 0.0143235
R2484 VDD.n404 VDD.n401 0.0143235
R2485 VDD.n420 VDD.n417 0.0143235
R2486 VDD.n434 VDD.n431 0.0143235
R2487 VDD.n471 VDD.n454 0.0143235
R2488 VDD.n1482 VDD.n1481 0.0143235
R2489 VDD.n495 VDD.n487 0.0143235
R2490 VDD.n1448 VDD.n1447 0.0143235
R2491 VDD.n519 VDD.n511 0.0143235
R2492 VDD.n549 VDD.n547 0.0143235
R2493 VDD.n565 VDD.n562 0.0143235
R2494 VDD.n581 VDD.n578 0.0143235
R2495 VDD.n597 VDD.n594 0.0143235
R2496 VDD.n611 VDD.n608 0.0143235
R2497 VDD.n648 VDD.n631 0.0143235
R2498 VDD.n1319 VDD.n1318 0.0143235
R2499 VDD.n672 VDD.n664 0.0143235
R2500 VDD.n1285 VDD.n1284 0.0143235
R2501 VDD.n696 VDD.n688 0.0143235
R2502 VDD.n726 VDD.n724 0.0143235
R2503 VDD.n742 VDD.n739 0.0143235
R2504 VDD.n758 VDD.n755 0.0143235
R2505 VDD.n774 VDD.n771 0.0143235
R2506 VDD.n788 VDD.n785 0.0143235
R2507 VDD.n825 VDD.n808 0.0143235
R2508 VDD.n1156 VDD.n1155 0.0143235
R2509 VDD.n849 VDD.n841 0.0143235
R2510 VDD.n1122 VDD.n1121 0.0143235
R2511 VDD.n874 VDD.n866 0.0143235
R2512 VDD.n1079 VDD.n1078 0.0143235
R2513 VDD.n917 VDD.n909 0.0143235
R2514 VDD.n1058 VDD.n1057 0.0143235
R2515 VDD.n956 VDD.n948 0.0143235
R2516 VDD.n1037 VDD.n1036 0.0143235
R2517 VDD.n1719 VDD.n1718 0.0140975
R2518 VDD.n1756 VDD.n9 0.0140135
R2519 VDD.n195 VDD.n194 0.0137576
R2520 VDD.n215 VDD.n214 0.0137576
R2521 VDD.n1697 VDD.n166 0.0137576
R2522 VDD.n1688 VDD.n1687 0.0137576
R2523 VDD.n1676 VDD.n250 0.0137576
R2524 VDD.n292 VDD.n291 0.0137576
R2525 VDD.n1632 VDD.n1631 0.0137576
R2526 VDD.n316 VDD.n315 0.0137576
R2527 VDD.n1598 VDD.n1597 0.0137576
R2528 VDD.n340 VDD.n339 0.0137576
R2529 VDD.n354 VDD.n353 0.0137576
R2530 VDD.n352 VDD.n349 0.0137576
R2531 VDD.n1563 VDD.n369 0.0137576
R2532 VDD.n1551 VDD.n384 0.0137576
R2533 VDD.n1539 VDD.n400 0.0137576
R2534 VDD.n1527 VDD.n416 0.0137576
R2535 VDD.n1513 VDD.n430 0.0137576
R2536 VDD.n469 VDD.n468 0.0137576
R2537 VDD.n1469 VDD.n1468 0.0137576
R2538 VDD.n493 VDD.n492 0.0137576
R2539 VDD.n1435 VDD.n1434 0.0137576
R2540 VDD.n517 VDD.n516 0.0137576
R2541 VDD.n531 VDD.n530 0.0137576
R2542 VDD.n529 VDD.n526 0.0137576
R2543 VDD.n1400 VDD.n546 0.0137576
R2544 VDD.n1388 VDD.n561 0.0137576
R2545 VDD.n1376 VDD.n577 0.0137576
R2546 VDD.n1364 VDD.n593 0.0137576
R2547 VDD.n1350 VDD.n607 0.0137576
R2548 VDD.n646 VDD.n645 0.0137576
R2549 VDD.n1306 VDD.n1305 0.0137576
R2550 VDD.n670 VDD.n669 0.0137576
R2551 VDD.n1272 VDD.n1271 0.0137576
R2552 VDD.n694 VDD.n693 0.0137576
R2553 VDD.n708 VDD.n707 0.0137576
R2554 VDD.n706 VDD.n703 0.0137576
R2555 VDD.n1237 VDD.n723 0.0137576
R2556 VDD.n1225 VDD.n738 0.0137576
R2557 VDD.n1213 VDD.n754 0.0137576
R2558 VDD.n1201 VDD.n770 0.0137576
R2559 VDD.n1187 VDD.n784 0.0137576
R2560 VDD.n823 VDD.n822 0.0137576
R2561 VDD.n1143 VDD.n1142 0.0137576
R2562 VDD.n847 VDD.n846 0.0137576
R2563 VDD.n1109 VDD.n1108 0.0137576
R2564 VDD.n872 VDD.n871 0.0137576
R2565 VDD.n896 VDD.n880 0.0137576
R2566 VDD.n915 VDD.n914 0.0137576
R2567 VDD.n935 VDD.n934 0.0137576
R2568 VDD.n954 VDD.n953 0.0137576
R2569 VDD.n1023 VDD.n1022 0.0137576
R2570 VDD.n973 VDD.n972 0.0137576
R2571 VDD.n46 VDD.n42 0.0137243
R2572 VDD.n1755 VDD.n11 0.0137188
R2573 VDD.n1755 VDD.n13 0.0137188
R2574 VDD.n1751 VDD.n1750 0.0130393
R2575 VDD.n17 VDD.n14 0.0130393
R2576 VDD.n1716 VDD.n1715 0.0129151
R2577 VDD.n198 VDD.n183 0.0125513
R2578 VDD.n218 VDD.n173 0.0125513
R2579 VDD.n225 VDD.n171 0.0125513
R2580 VDD.n1692 VDD.n226 0.0125513
R2581 VDD.n259 VDD.n258 0.0125513
R2582 VDD.n296 VDD.n295 0.0125513
R2583 VDD.n1646 VDD.n297 0.0125513
R2584 VDD.n320 VDD.n319 0.0125513
R2585 VDD.n1612 VDD.n321 0.0125513
R2586 VDD.n344 VDD.n343 0.0125513
R2587 VDD.n374 VDD.n373 0.0125513
R2588 VDD.n390 VDD.n389 0.0125513
R2589 VDD.n406 VDD.n405 0.0125513
R2590 VDD.n422 VDD.n421 0.0125513
R2591 VDD.n436 VDD.n435 0.0125513
R2592 VDD.n473 VDD.n472 0.0125513
R2593 VDD.n1483 VDD.n474 0.0125513
R2594 VDD.n497 VDD.n496 0.0125513
R2595 VDD.n1449 VDD.n498 0.0125513
R2596 VDD.n521 VDD.n520 0.0125513
R2597 VDD.n551 VDD.n550 0.0125513
R2598 VDD.n567 VDD.n566 0.0125513
R2599 VDD.n583 VDD.n582 0.0125513
R2600 VDD.n599 VDD.n598 0.0125513
R2601 VDD.n613 VDD.n612 0.0125513
R2602 VDD.n650 VDD.n649 0.0125513
R2603 VDD.n1320 VDD.n651 0.0125513
R2604 VDD.n674 VDD.n673 0.0125513
R2605 VDD.n1286 VDD.n675 0.0125513
R2606 VDD.n698 VDD.n697 0.0125513
R2607 VDD.n728 VDD.n727 0.0125513
R2608 VDD.n744 VDD.n743 0.0125513
R2609 VDD.n760 VDD.n759 0.0125513
R2610 VDD.n776 VDD.n775 0.0125513
R2611 VDD.n790 VDD.n789 0.0125513
R2612 VDD.n827 VDD.n826 0.0125513
R2613 VDD.n1157 VDD.n828 0.0125513
R2614 VDD.n851 VDD.n850 0.0125513
R2615 VDD.n1123 VDD.n852 0.0125513
R2616 VDD.n876 VDD.n875 0.0125513
R2617 VDD.n1080 VDD.n882 0.0121049
R2618 VDD.n919 VDD.n918 0.0121049
R2619 VDD.n1059 VDD.n920 0.0121049
R2620 VDD.n958 VDD.n957 0.0121049
R2621 VDD.n1038 VDD.n959 0.0121049
R2622 VDD.n48 VDD.n43 0.0105714
R2623 VDD.n1729 VDD.n1728 0.0103794
R2624 VDD.n62 VDD.n59 0.0103794
R2625 VDD.n998 VDD.n66 0.0103794
R2626 VDD.n995 VDD.n70 0.0103794
R2627 VDD.n991 VDD.n74 0.0103794
R2628 VDD.n899 VDD.n898 0.0099697
R2629 VDD.n1067 VDD.n905 0.0099697
R2630 VDD.n938 VDD.n937 0.0099697
R2631 VDD.n1046 VDD.n944 0.0099697
R2632 VDD.n1026 VDD.n1025 0.0099697
R2633 VDD.n192 VDD.n191 0.0099697
R2634 VDD.n211 VDD.n210 0.0099697
R2635 VDD.n1699 VDD.n165 0.0099697
R2636 VDD.n242 VDD.n231 0.0099697
R2637 VDD.n1679 VDD.n1678 0.0099697
R2638 VDD.n1667 VDD.n1666 0.0099697
R2639 VDD.n270 VDD.n268 0.0099697
R2640 VDD.n1654 VDD.n273 0.0099697
R2641 VDD.n1635 VDD.n1634 0.0099697
R2642 VDD.n1620 VDD.n306 0.0099697
R2643 VDD.n1601 VDD.n1600 0.0099697
R2644 VDD.n1586 VDD.n330 0.0099697
R2645 VDD.n1566 VDD.n1565 0.0099697
R2646 VDD.n1554 VDD.n1553 0.0099697
R2647 VDD.n1542 VDD.n1541 0.0099697
R2648 VDD.n1530 VDD.n1529 0.0099697
R2649 VDD.n1516 VDD.n1515 0.0099697
R2650 VDD.n1504 VDD.n1503 0.0099697
R2651 VDD.n447 VDD.n445 0.0099697
R2652 VDD.n1491 VDD.n450 0.0099697
R2653 VDD.n1472 VDD.n1471 0.0099697
R2654 VDD.n1457 VDD.n483 0.0099697
R2655 VDD.n1438 VDD.n1437 0.0099697
R2656 VDD.n1423 VDD.n507 0.0099697
R2657 VDD.n1403 VDD.n1402 0.0099697
R2658 VDD.n1391 VDD.n1390 0.0099697
R2659 VDD.n1379 VDD.n1378 0.0099697
R2660 VDD.n1367 VDD.n1366 0.0099697
R2661 VDD.n1353 VDD.n1352 0.0099697
R2662 VDD.n1341 VDD.n1340 0.0099697
R2663 VDD.n624 VDD.n622 0.0099697
R2664 VDD.n1328 VDD.n627 0.0099697
R2665 VDD.n1309 VDD.n1308 0.0099697
R2666 VDD.n1294 VDD.n660 0.0099697
R2667 VDD.n1275 VDD.n1274 0.0099697
R2668 VDD.n1260 VDD.n684 0.0099697
R2669 VDD.n1240 VDD.n1239 0.0099697
R2670 VDD.n1228 VDD.n1227 0.0099697
R2671 VDD.n1216 VDD.n1215 0.0099697
R2672 VDD.n1204 VDD.n1203 0.0099697
R2673 VDD.n1190 VDD.n1189 0.0099697
R2674 VDD.n1178 VDD.n1177 0.0099697
R2675 VDD.n801 VDD.n799 0.0099697
R2676 VDD.n1165 VDD.n804 0.0099697
R2677 VDD.n1146 VDD.n1145 0.0099697
R2678 VDD.n1131 VDD.n837 0.0099697
R2679 VDD.n1112 VDD.n1111 0.0099697
R2680 VDD.n1097 VDD.n861 0.0099697
R2681 VDD.n1744 VDD.n27 0.00701042
R2682 VDD.n1758 VDD.n6 0.00701042
R2683 VDD.n1727 VDD.n38 0.00635126
R2684 VDD.n1723 VDD.n58 0.00635126
R2685 VDD.n1720 VDD.n65 0.00635126
R2686 VDD.n1717 VDD.n69 0.00635126
R2687 VDD.n1714 VDD.n73 0.00635126
R2688 VDD.n1713 VDD.n72 0.00493396
R2689 VDD.n1715 VDD.n72 0.00493396
R2690 VDD.n1716 VDD.n68 0.00493396
R2691 VDD.n1718 VDD.n68 0.00493396
R2692 VDD.n1719 VDD.n64 0.00493396
R2693 VDD.n1721 VDD.n64 0.00493396
R2694 VDD.n1722 VDD.n57 0.00493396
R2695 VDD.n1724 VDD.n57 0.00493396
R2696 VDD.n1726 VDD.n1725 0.00493396
R2697 VDD.n1725 VDD.n56 0.00493396
R2698 VDD.n55 VDD.n39 0.00493396
R2699 VDD.n50 VDD.n39 0.00493396
R2700 VDD.n25 VDD.n24 0.00490305
R2701 VDD.n1758 VDD.n1757 0.00440625
R2702 VDD.n79 VDD.n78 0.00428788
R2703 VDD.n203 VDD.n181 0.00428788
R2704 VDD.n213 VDD.n164 0.00428788
R2705 VDD.n1696 VDD.n168 0.00428788
R2706 VDD.n232 VDD.n230 0.00428788
R2707 VDD.n1673 VDD.n1672 0.00428788
R2708 VDD.n289 VDD.n269 0.00428788
R2709 VDD.n1651 VDD.n276 0.00428788
R2710 VDD.n1642 VDD.n301 0.00428788
R2711 VDD.n1617 VDD.n309 0.00428788
R2712 VDD.n1608 VDD.n325 0.00428788
R2713 VDD.n1583 VDD.n333 0.00428788
R2714 VDD.n1572 VDD.n1571 0.00428788
R2715 VDD.n1560 VDD.n1559 0.00428788
R2716 VDD.n1548 VDD.n1547 0.00428788
R2717 VDD.n1536 VDD.n1535 0.00428788
R2718 VDD.n1524 VDD.n1523 0.00428788
R2719 VDD.n1510 VDD.n1509 0.00428788
R2720 VDD.n466 VDD.n446 0.00428788
R2721 VDD.n1488 VDD.n453 0.00428788
R2722 VDD.n1479 VDD.n478 0.00428788
R2723 VDD.n1454 VDD.n486 0.00428788
R2724 VDD.n1445 VDD.n502 0.00428788
R2725 VDD.n1420 VDD.n510 0.00428788
R2726 VDD.n1409 VDD.n1408 0.00428788
R2727 VDD.n1397 VDD.n1396 0.00428788
R2728 VDD.n1385 VDD.n1384 0.00428788
R2729 VDD.n1373 VDD.n1372 0.00428788
R2730 VDD.n1361 VDD.n1360 0.00428788
R2731 VDD.n1347 VDD.n1346 0.00428788
R2732 VDD.n643 VDD.n623 0.00428788
R2733 VDD.n1325 VDD.n630 0.00428788
R2734 VDD.n1316 VDD.n655 0.00428788
R2735 VDD.n1291 VDD.n663 0.00428788
R2736 VDD.n1282 VDD.n679 0.00428788
R2737 VDD.n1257 VDD.n687 0.00428788
R2738 VDD.n1246 VDD.n1245 0.00428788
R2739 VDD.n1234 VDD.n1233 0.00428788
R2740 VDD.n1222 VDD.n1221 0.00428788
R2741 VDD.n1210 VDD.n1209 0.00428788
R2742 VDD.n1198 VDD.n1197 0.00428788
R2743 VDD.n1184 VDD.n1183 0.00428788
R2744 VDD.n820 VDD.n800 0.00428788
R2745 VDD.n1162 VDD.n807 0.00428788
R2746 VDD.n1153 VDD.n832 0.00428788
R2747 VDD.n1128 VDD.n840 0.00428788
R2748 VDD.n1119 VDD.n856 0.00428788
R2749 VDD.n1094 VDD.n865 0.00428788
R2750 VDD.n1084 VDD.n1083 0.00428788
R2751 VDD.n1076 VDD.n885 0.00428788
R2752 VDD.n1064 VDD.n908 0.00428788
R2753 VDD.n1055 VDD.n924 0.00428788
R2754 VDD.n1043 VDD.n947 0.00428788
R2755 VDD.n1034 VDD.n963 0.00428788
R2756 VDD.n21 VDD.n20 0.00428087
R2757 VDD.n984 VDD.n983 0.00391036
R2758 VDD.n969 VDD 0.00377907
R2759 VDD.n1750 VDD.n24 0.00360776
R2760 VDD.n21 VDD.n14 0.00360776
R2761 VDD.n48 VDD.n41 0.00351641
R2762 VDD.n294 VDD.n293 0.00326471
R2763 VDD.n1645 VDD.n298 0.00326471
R2764 VDD.n318 VDD.n317 0.00326471
R2765 VDD.n1611 VDD.n322 0.00326471
R2766 VDD.n342 VDD.n341 0.00326471
R2767 VDD.n1577 VDD.n345 0.00326471
R2768 VDD.n471 VDD.n470 0.00326471
R2769 VDD.n1482 VDD.n475 0.00326471
R2770 VDD.n495 VDD.n494 0.00326471
R2771 VDD.n1448 VDD.n499 0.00326471
R2772 VDD.n519 VDD.n518 0.00326471
R2773 VDD.n1414 VDD.n522 0.00326471
R2774 VDD.n648 VDD.n647 0.00326471
R2775 VDD.n1319 VDD.n652 0.00326471
R2776 VDD.n672 VDD.n671 0.00326471
R2777 VDD.n1285 VDD.n676 0.00326471
R2778 VDD.n696 VDD.n695 0.00326471
R2779 VDD.n1251 VDD.n699 0.00326471
R2780 VDD.n825 VDD.n824 0.00326471
R2781 VDD.n1156 VDD.n829 0.00326471
R2782 VDD.n849 VDD.n848 0.00326471
R2783 VDD.n1122 VDD.n853 0.00326471
R2784 VDD.n874 VDD.n873 0.00326471
R2785 VDD.n1079 VDD.n881 0.00326471
R2786 VDD.n917 VDD.n916 0.00326471
R2787 VDD.n1058 VDD.n921 0.00326471
R2788 VDD.n956 VDD.n955 0.00326471
R2789 VDD.n1037 VDD.n960 0.00326471
R2790 VDD.n979 VDD.n974 0.00326471
R2791 VDD.n197 VDD.n196 0.00257353
R2792 VDD.n217 VDD.n216 0.00257353
R2793 VDD.n224 VDD.n169 0.00257353
R2794 VDD.n1690 VDD.n1689 0.00257353
R2795 VDD.n1675 VDD.n251 0.00257353
R2796 VDD.n1576 VDD.n346 0.00257353
R2797 VDD.n1562 VDD.n370 0.00257353
R2798 VDD.n1550 VDD.n385 0.00257353
R2799 VDD.n1538 VDD.n401 0.00257353
R2800 VDD.n1526 VDD.n417 0.00257353
R2801 VDD.n1512 VDD.n431 0.00257353
R2802 VDD.n1413 VDD.n523 0.00257353
R2803 VDD.n1399 VDD.n547 0.00257353
R2804 VDD.n1387 VDD.n562 0.00257353
R2805 VDD.n1375 VDD.n578 0.00257353
R2806 VDD.n1363 VDD.n594 0.00257353
R2807 VDD.n1349 VDD.n608 0.00257353
R2808 VDD.n1250 VDD.n700 0.00257353
R2809 VDD.n1236 VDD.n724 0.00257353
R2810 VDD.n1224 VDD.n739 0.00257353
R2811 VDD.n1212 VDD.n755 0.00257353
R2812 VDD.n1200 VDD.n771 0.00257353
R2813 VDD.n1186 VDD.n785 0.00257353
R2814 VDD.n1075 VDD.n886 0.00239394
R2815 VDD.n1066 VDD.n906 0.00239394
R2816 VDD.n1054 VDD.n925 0.00239394
R2817 VDD.n1045 VDD.n945 0.00239394
R2818 VDD.n1033 VDD.n964 0.00239394
R2819 VDD.n1709 VDD.n80 0.00239394
R2820 VDD.n204 VDD.n176 0.00239394
R2821 VDD.n1703 VDD.n1702 0.00239394
R2822 VDD.n241 VDD.n167 0.00239394
R2823 VDD.n1685 VDD.n233 0.00239394
R2824 VDD.n1671 VDD.n263 0.00239394
R2825 VDD.n1662 VDD.n271 0.00239394
R2826 VDD.n1653 VDD.n274 0.00239394
R2827 VDD.n1641 VDD.n302 0.00239394
R2828 VDD.n1619 VDD.n307 0.00239394
R2829 VDD.n1607 VDD.n326 0.00239394
R2830 VDD.n1585 VDD.n331 0.00239394
R2831 VDD.n1570 VDD.n357 0.00239394
R2832 VDD.n1558 VDD.n378 0.00239394
R2833 VDD.n1546 VDD.n394 0.00239394
R2834 VDD.n1534 VDD.n410 0.00239394
R2835 VDD.n1522 VDD.n426 0.00239394
R2836 VDD.n1508 VDD.n440 0.00239394
R2837 VDD.n1499 VDD.n448 0.00239394
R2838 VDD.n1490 VDD.n451 0.00239394
R2839 VDD.n1478 VDD.n479 0.00239394
R2840 VDD.n1456 VDD.n484 0.00239394
R2841 VDD.n1444 VDD.n503 0.00239394
R2842 VDD.n1422 VDD.n508 0.00239394
R2843 VDD.n1407 VDD.n534 0.00239394
R2844 VDD.n1395 VDD.n555 0.00239394
R2845 VDD.n1383 VDD.n571 0.00239394
R2846 VDD.n1371 VDD.n587 0.00239394
R2847 VDD.n1359 VDD.n603 0.00239394
R2848 VDD.n1345 VDD.n617 0.00239394
R2849 VDD.n1336 VDD.n625 0.00239394
R2850 VDD.n1327 VDD.n628 0.00239394
R2851 VDD.n1315 VDD.n656 0.00239394
R2852 VDD.n1293 VDD.n661 0.00239394
R2853 VDD.n1281 VDD.n680 0.00239394
R2854 VDD.n1259 VDD.n685 0.00239394
R2855 VDD.n1244 VDD.n711 0.00239394
R2856 VDD.n1232 VDD.n732 0.00239394
R2857 VDD.n1220 VDD.n748 0.00239394
R2858 VDD.n1208 VDD.n764 0.00239394
R2859 VDD.n1196 VDD.n780 0.00239394
R2860 VDD.n1182 VDD.n794 0.00239394
R2861 VDD.n1173 VDD.n802 0.00239394
R2862 VDD.n1164 VDD.n805 0.00239394
R2863 VDD.n1152 VDD.n833 0.00239394
R2864 VDD.n1130 VDD.n838 0.00239394
R2865 VDD.n1118 VDD.n857 0.00239394
R2866 VDD.n1096 VDD.n863 0.00239394
R2867 VDD.n188 VDD.n79 0.00239394
R2868 VDD.n203 VDD.n175 0.00239394
R2869 VDD.n1701 VDD.n164 0.00239394
R2870 VDD.n240 VDD.n168 0.00239394
R2871 VDD.n249 VDD.n232 0.00239394
R2872 VDD.n1672 VDD.n261 0.00239394
R2873 VDD.n1663 VDD.n269 0.00239394
R2874 VDD.n1652 VDD.n1651 0.00239394
R2875 VDD.n1642 VDD.n300 0.00239394
R2876 VDD.n1618 VDD.n1617 0.00239394
R2877 VDD.n1608 VDD.n324 0.00239394
R2878 VDD.n1584 VDD.n1583 0.00239394
R2879 VDD.n1571 VDD.n350 0.00239394
R2880 VDD.n1559 VDD.n376 0.00239394
R2881 VDD.n1547 VDD.n392 0.00239394
R2882 VDD.n1535 VDD.n408 0.00239394
R2883 VDD.n1523 VDD.n424 0.00239394
R2884 VDD.n1509 VDD.n438 0.00239394
R2885 VDD.n1500 VDD.n446 0.00239394
R2886 VDD.n1489 VDD.n1488 0.00239394
R2887 VDD.n1479 VDD.n477 0.00239394
R2888 VDD.n1455 VDD.n1454 0.00239394
R2889 VDD.n1445 VDD.n501 0.00239394
R2890 VDD.n1421 VDD.n1420 0.00239394
R2891 VDD.n1408 VDD.n527 0.00239394
R2892 VDD.n1396 VDD.n553 0.00239394
R2893 VDD.n1384 VDD.n569 0.00239394
R2894 VDD.n1372 VDD.n585 0.00239394
R2895 VDD.n1360 VDD.n601 0.00239394
R2896 VDD.n1346 VDD.n615 0.00239394
R2897 VDD.n1337 VDD.n623 0.00239394
R2898 VDD.n1326 VDD.n1325 0.00239394
R2899 VDD.n1316 VDD.n654 0.00239394
R2900 VDD.n1292 VDD.n1291 0.00239394
R2901 VDD.n1282 VDD.n678 0.00239394
R2902 VDD.n1258 VDD.n1257 0.00239394
R2903 VDD.n1245 VDD.n704 0.00239394
R2904 VDD.n1233 VDD.n730 0.00239394
R2905 VDD.n1221 VDD.n746 0.00239394
R2906 VDD.n1209 VDD.n762 0.00239394
R2907 VDD.n1197 VDD.n778 0.00239394
R2908 VDD.n1183 VDD.n792 0.00239394
R2909 VDD.n1174 VDD.n800 0.00239394
R2910 VDD.n1163 VDD.n1162 0.00239394
R2911 VDD.n1153 VDD.n831 0.00239394
R2912 VDD.n1129 VDD.n1128 0.00239394
R2913 VDD.n1119 VDD.n855 0.00239394
R2914 VDD.n1095 VDD.n1094 0.00239394
R2915 VDD.n1076 VDD.n884 0.00239394
R2916 VDD.n1065 VDD.n1064 0.00239394
R2917 VDD.n1055 VDD.n923 0.00239394
R2918 VDD.n1044 VDD.n1043 0.00239394
R2919 VDD.n1034 VDD.n962 0.00239394
R2920 VDD.n978 VDD.n971 0.00224074
R2921 VDD.n54 VDD.n51 0.0021514
R2922 VDD.n980 VDD.n970 0.00213953
R2923 VDD.n1752 VDD.n11 0.00196875
R2924 VDD.n16 VDD.n13 0.00196875
R2925 VDD VDD.n1712 0.00170513
R2926 VDD.n1575 VDD 0.00170513
R2927 VDD.n1412 VDD 0.00170513
R2928 VDD.n1249 VDD 0.00170513
R2929 VDD.n185 VDD.n77 0.00119118
R2930 VDD.n186 VDD.n185 0.00119118
R2931 VDD.n201 VDD.n182 0.00119118
R2932 VDD.n202 VDD.n201 0.00119118
R2933 VDD.n221 VDD.n172 0.00119118
R2934 VDD.n222 VDD.n221 0.00119118
R2935 VDD.n1695 VDD.n170 0.00119118
R2936 VDD.n227 VDD.n170 0.00119118
R2937 VDD.n255 VDD.n228 0.00119118
R2938 VDD.n256 VDD.n255 0.00119118
R2939 VDD.n1674 VDD.n252 0.00119118
R2940 VDD.n262 VDD.n252 0.00119118
R2941 VDD.n287 VDD.n280 0.00119118
R2942 VDD.n288 VDD.n287 0.00119118
R2943 VDD.n1650 VDD.n1649 0.00119118
R2944 VDD.n1649 VDD.n278 0.00119118
R2945 VDD.n1643 VDD.n299 0.00119118
R2946 VDD.n314 VDD.n299 0.00119118
R2947 VDD.n1616 VDD.n1615 0.00119118
R2948 VDD.n1615 VDD.n311 0.00119118
R2949 VDD.n1609 VDD.n323 0.00119118
R2950 VDD.n338 VDD.n323 0.00119118
R2951 VDD.n1582 VDD.n1581 0.00119118
R2952 VDD.n1581 VDD.n335 0.00119118
R2953 VDD.n1573 VDD.n348 0.00119118
R2954 VDD.n351 VDD.n348 0.00119118
R2955 VDD.n1561 VDD.n371 0.00119118
R2956 VDD.n377 VDD.n371 0.00119118
R2957 VDD.n1549 VDD.n386 0.00119118
R2958 VDD.n393 VDD.n386 0.00119118
R2959 VDD.n1537 VDD.n402 0.00119118
R2960 VDD.n409 VDD.n402 0.00119118
R2961 VDD.n1525 VDD.n418 0.00119118
R2962 VDD.n425 VDD.n418 0.00119118
R2963 VDD.n1511 VDD.n432 0.00119118
R2964 VDD.n439 VDD.n432 0.00119118
R2965 VDD.n464 VDD.n457 0.00119118
R2966 VDD.n465 VDD.n464 0.00119118
R2967 VDD.n1487 VDD.n1486 0.00119118
R2968 VDD.n1486 VDD.n455 0.00119118
R2969 VDD.n1480 VDD.n476 0.00119118
R2970 VDD.n491 VDD.n476 0.00119118
R2971 VDD.n1453 VDD.n1452 0.00119118
R2972 VDD.n1452 VDD.n488 0.00119118
R2973 VDD.n1446 VDD.n500 0.00119118
R2974 VDD.n515 VDD.n500 0.00119118
R2975 VDD.n1419 VDD.n1418 0.00119118
R2976 VDD.n1418 VDD.n512 0.00119118
R2977 VDD.n1410 VDD.n525 0.00119118
R2978 VDD.n528 VDD.n525 0.00119118
R2979 VDD.n1398 VDD.n548 0.00119118
R2980 VDD.n554 VDD.n548 0.00119118
R2981 VDD.n1386 VDD.n563 0.00119118
R2982 VDD.n570 VDD.n563 0.00119118
R2983 VDD.n1374 VDD.n579 0.00119118
R2984 VDD.n586 VDD.n579 0.00119118
R2985 VDD.n1362 VDD.n595 0.00119118
R2986 VDD.n602 VDD.n595 0.00119118
R2987 VDD.n1348 VDD.n609 0.00119118
R2988 VDD.n616 VDD.n609 0.00119118
R2989 VDD.n641 VDD.n634 0.00119118
R2990 VDD.n642 VDD.n641 0.00119118
R2991 VDD.n1324 VDD.n1323 0.00119118
R2992 VDD.n1323 VDD.n632 0.00119118
R2993 VDD.n1317 VDD.n653 0.00119118
R2994 VDD.n668 VDD.n653 0.00119118
R2995 VDD.n1290 VDD.n1289 0.00119118
R2996 VDD.n1289 VDD.n665 0.00119118
R2997 VDD.n1283 VDD.n677 0.00119118
R2998 VDD.n692 VDD.n677 0.00119118
R2999 VDD.n1256 VDD.n1255 0.00119118
R3000 VDD.n1255 VDD.n689 0.00119118
R3001 VDD.n1247 VDD.n702 0.00119118
R3002 VDD.n705 VDD.n702 0.00119118
R3003 VDD.n1235 VDD.n725 0.00119118
R3004 VDD.n731 VDD.n725 0.00119118
R3005 VDD.n1223 VDD.n740 0.00119118
R3006 VDD.n747 VDD.n740 0.00119118
R3007 VDD.n1211 VDD.n756 0.00119118
R3008 VDD.n763 VDD.n756 0.00119118
R3009 VDD.n1199 VDD.n772 0.00119118
R3010 VDD.n779 VDD.n772 0.00119118
R3011 VDD.n1185 VDD.n786 0.00119118
R3012 VDD.n793 VDD.n786 0.00119118
R3013 VDD.n818 VDD.n811 0.00119118
R3014 VDD.n819 VDD.n818 0.00119118
R3015 VDD.n1161 VDD.n1160 0.00119118
R3016 VDD.n1160 VDD.n809 0.00119118
R3017 VDD.n1154 VDD.n830 0.00119118
R3018 VDD.n845 VDD.n830 0.00119118
R3019 VDD.n1127 VDD.n1126 0.00119118
R3020 VDD.n1126 VDD.n842 0.00119118
R3021 VDD.n1120 VDD.n854 0.00119118
R3022 VDD.n870 VDD.n854 0.00119118
R3023 VDD.n1093 VDD.n1092 0.00119118
R3024 VDD.n1092 VDD.n867 0.00119118
R3025 VDD.n1085 VDD.n878 0.00119118
R3026 VDD.n1082 VDD.n878 0.00119118
R3027 VDD.n1077 VDD.n883 0.00119118
R3028 VDD.n913 VDD.n883 0.00119118
R3029 VDD.n1063 VDD.n1062 0.00119118
R3030 VDD.n1062 VDD.n910 0.00119118
R3031 VDD.n1056 VDD.n922 0.00119118
R3032 VDD.n952 VDD.n922 0.00119118
R3033 VDD.n1042 VDD.n1041 0.00119118
R3034 VDD.n1041 VDD.n949 0.00119118
R3035 VDD.n1035 VDD.n961 0.00119118
R3036 VDD.n976 VDD.n961 0.00119118
R3037 VDD.n44 VDD.n42 0.0011215
R3038 VDD.n184 VDD.n76 0.00110256
R3039 VDD.n200 VDD.n199 0.00110256
R3040 VDD.n220 VDD.n219 0.00110256
R3041 VDD.n1694 VDD.n1693 0.00110256
R3042 VDD.n254 VDD.n253 0.00110256
R3043 VDD.n281 VDD.n260 0.00110256
R3044 VDD.n286 VDD.n279 0.00110256
R3045 VDD.n1648 VDD.n1647 0.00110256
R3046 VDD.n313 VDD.n312 0.00110256
R3047 VDD.n1614 VDD.n1613 0.00110256
R3048 VDD.n337 VDD.n336 0.00110256
R3049 VDD.n1580 VDD.n1579 0.00110256
R3050 VDD.n1574 VDD.n347 0.00110256
R3051 VDD.n387 VDD.n375 0.00110256
R3052 VDD.n403 VDD.n391 0.00110256
R3053 VDD.n419 VDD.n407 0.00110256
R3054 VDD.n433 VDD.n423 0.00110256
R3055 VDD.n458 VDD.n437 0.00110256
R3056 VDD.n463 VDD.n456 0.00110256
R3057 VDD.n1485 VDD.n1484 0.00110256
R3058 VDD.n490 VDD.n489 0.00110256
R3059 VDD.n1451 VDD.n1450 0.00110256
R3060 VDD.n514 VDD.n513 0.00110256
R3061 VDD.n1417 VDD.n1416 0.00110256
R3062 VDD.n1411 VDD.n524 0.00110256
R3063 VDD.n564 VDD.n552 0.00110256
R3064 VDD.n580 VDD.n568 0.00110256
R3065 VDD.n596 VDD.n584 0.00110256
R3066 VDD.n610 VDD.n600 0.00110256
R3067 VDD.n635 VDD.n614 0.00110256
R3068 VDD.n640 VDD.n633 0.00110256
R3069 VDD.n1322 VDD.n1321 0.00110256
R3070 VDD.n667 VDD.n666 0.00110256
R3071 VDD.n1288 VDD.n1287 0.00110256
R3072 VDD.n691 VDD.n690 0.00110256
R3073 VDD.n1254 VDD.n1253 0.00110256
R3074 VDD.n1248 VDD.n701 0.00110256
R3075 VDD.n741 VDD.n729 0.00110256
R3076 VDD.n757 VDD.n745 0.00110256
R3077 VDD.n773 VDD.n761 0.00110256
R3078 VDD.n787 VDD.n777 0.00110256
R3079 VDD.n812 VDD.n791 0.00110256
R3080 VDD.n817 VDD.n810 0.00110256
R3081 VDD.n1159 VDD.n1158 0.00110256
R3082 VDD.n844 VDD.n843 0.00110256
R3083 VDD.n1125 VDD.n1124 0.00110256
R3084 VDD.n869 VDD.n868 0.00110256
R3085 VDD.n1091 VDD.n1090 0.00110256
R3086 VDD.n1081 VDD.n877 0.00108025
R3087 VDD.n912 VDD.n911 0.00108025
R3088 VDD.n1061 VDD.n1060 0.00108025
R3089 VDD.n951 VDD.n950 0.00108025
R3090 VDD.n1040 VDD.n1039 0.00108025
R3091 VDD.n977 VDD.n975 0.00108025
R3092 VDD.n1754 VDD.n1753 0.000837321
R3093 VDD VDD.n22 0.00072488
R3094 VDD.n1754 VDD.n22 0.00061244
R3095 code[2] code[2].t1 140.387
R3096 code[2].n1 code[2].t2 140.34
R3097 code[2].n0 code[2].t0 140.34
R3098 code[2].n2 code[2].t3 140.34
R3099 code[2].n2 code[2] 2.82659
R3100 code[2].n1 code[2] 0.285826
R3101 code[2].n2 code[2].n0 0.264087
R3102 code[2].n0 code[2] 0.0466957
R3103 code[2] code[2].n1 0.0466957
R3104 code[2] code[2].n2 0.0371379
R3105 VSS.n617 VSS.n616 1265.93
R3106 VSS.n684 VSS 1043.16
R3107 VSS.n710 VSS.t9 641.946
R3108 VSS.n623 VSS.t4 569.832
R3109 VSS.n637 VSS.n636 362.961
R3110 VSS.n567 VSS.t1 359.05
R3111 VSS.n710 VSS 320.974
R3112 VSS.n626 VSS.n625 292.5
R3113 VSS.n628 VSS.n627 292.5
R3114 VSS.n630 VSS.n629 292.5
R3115 VSS.n633 VSS.n632 292.5
R3116 VSS.n635 VSS.n634 292.5
R3117 VSS.n712 VSS.n711 292.5
R3118 VSS.n711 VSS.n710 292.5
R3119 VSS.n622 VSS 255.776
R3120 VSS.t4 VSS.t3 233.113
R3121 VSS.n662 VSS.n661 200.608
R3122 VSS.n624 VSS.n623 197.27
R3123 VSS.n686 VSS.n685 173.861
R3124 VSS.n686 VSS.t6 147.113
R3125 VSS.t3 VSS.n622 132.745
R3126 VSS.n568 VSS.n567 126.269
R3127 VSS.t1 VSS.t8 112.822
R3128 VSS.n679 VSS.t7 107.867
R3129 VSS.n712 VSS.t10 107.195
R3130 VSS.n663 VSS.n659 93.0283
R3131 VSS.n624 VSS.n9 92.1828
R3132 VSS.n626 VSS.n624 81.7271
R3133 VSS.n531 VSS.t12 77.3934
R3134 VSS.n531 VSS.t11 77.3934
R3135 VSS.n687 VSS.n683 71.1394
R3136 VSS.n632 VSS.n631 69.3633
R3137 VSS.n685 VSS.n684 53.4959
R3138 VSS.n542 VSS.t2 43.7547
R3139 VSS.n638 VSS.n637 41.5854
R3140 VSS.n638 VSS.t5 41.4448
R3141 VSS.n630 VSS.n628 36.9236
R3142 VSS.n661 VSS.n660 26.7482
R3143 VSS.n620 VSS.n619 25.9019
R3144 VSS.n683 VSS.n682 21.8894
R3145 VSS.n46 VSS.n45 17.6402
R3146 VSS.n257 VSS.n60 17.6402
R3147 VSS.n90 VSS.n89 17.6402
R3148 VSS.n330 VSS.n329 17.6402
R3149 VSS.n199 VSS.n53 17.6397
R3150 VSS.n75 VSS.n74 17.6397
R3151 VSS.n290 VSS.n289 17.6397
R3152 VSS.n430 VSS.n429 17.6397
R3153 VSS.n558 VSS.n557 17.6348
R3154 VSS.n482 VSS.n455 17.6348
R3155 VSS.n400 VSS.n315 17.6348
R3156 VSS.n623 VSS.n621 12.9512
R3157 VSS.n637 VSS.n635 12.062
R3158 VSS.n628 VSS.n626 11.8159
R3159 VSS.n633 VSS.n630 11.8159
R3160 VSS.n635 VSS.n633 11.8159
R3161 VSS.n688 VSS.n687 9.3005
R3162 VSS.n687 VSS.n686 9.3005
R3163 VSS.n562 VSS.n561 9.15497
R3164 VSS.n52 VSS.n51 9.15497
R3165 VSS.n37 VSS.n36 9.15497
R3166 VSS.n66 VSS.n65 9.15497
R3167 VSS.n59 VSS.n58 9.15497
R3168 VSS.n96 VSS.n95 9.15497
R3169 VSS.n81 VSS.n80 9.15497
R3170 VSS.n30 VSS.n29 9.15497
R3171 VSS.n304 VSS.n303 9.15497
R3172 VSS.n559 VSS.n304 9.15497
R3173 VSS.n314 VSS.n313 9.15497
R3174 VSS.n336 VSS.n335 9.15497
R3175 VSS.n321 VSS.n320 9.15497
R3176 VSS.n23 VSS.n22 9.15497
R3177 VSS.n444 VSS.n443 9.15497
R3178 VSS.n559 VSS.n444 9.15497
R3179 VSS.n454 VSS.n453 9.15497
R3180 VSS.n16 VSS.n15 9.15497
R3181 VSS.n502 VSS.n501 9.15497
R3182 VSS.n559 VSS.n502 9.15497
R3183 VSS.n512 VSS.n511 9.15497
R3184 VSS.n570 VSS.n569 9.15497
R3185 VSS.n569 VSS.n568 9.15497
R3186 VSS.n615 VSS.n614 9.15497
R3187 VSS.n616 VSS.n615 9.15497
R3188 VSS.n664 VSS.n663 9.01392
R3189 VSS.n663 VSS.n662 9.01392
R3190 VSS.n315 VSS.n314 8.61509
R3191 VSS.n455 VSS.n454 8.61509
R3192 VSS.n558 VSS.n512 8.61509
R3193 VSS.n53 VSS.n52 8.48617
R3194 VSS.n75 VSS.n66 8.48617
R3195 VSS.n290 VSS.n96 8.48617
R3196 VSS.n430 VSS.n336 8.48617
R3197 VSS.n46 VSS.n37 8.48574
R3198 VSS.n60 VSS.n59 8.48574
R3199 VSS.n90 VSS.n81 8.48574
R3200 VSS.n330 VSS.n321 8.48574
R3201 VSS.n561 VSS.n560 8.48521
R3202 VSS VSS.n712 7.60922
R3203 VSS.n559 VSS.n31 6.48513
R3204 VSS.n559 VSS.n24 6.48513
R3205 VSS.n559 VSS.n17 6.48513
R3206 VSS.n618 VSS.n617 6.47585
R3207 VSS.n619 VSS.n618 6.47585
R3208 VSS.n621 VSS.n620 6.47585
R3209 VSS.n654 VSS.n653 4.6505
R3210 VSS.n690 VSS.n689 4.5005
R3211 VSS.n680 VSS.n679 3.72317
R3212 VSS.n664 VSS.n658 3.34819
R3213 VSS.n665 VSS.n657 3.15127
R3214 VSS.n401 VSS.n400 3.03311
R3215 VSS.n95 VSS.n94 3.03311
R3216 VSS.n65 VSS.n64 3.03311
R3217 VSS.n51 VSS.n50 3.03311
R3218 VSS.n483 VSS.n482 3.03311
R3219 VSS.n335 VSS.n334 3.03311
R3220 VSS.n557 VSS.n556 3.03311
R3221 VSS.n157 VSS.n154 3.03311
R3222 VSS.n563 VSS.n562 3.03311
R3223 VSS.n36 VSS.n35 3.03311
R3224 VSS.n45 VSS.n44 3.03311
R3225 VSS.n200 VSS.n199 3.03311
R3226 VSS.n58 VSS.n57 3.03311
R3227 VSS.n258 VSS.n257 3.03311
R3228 VSS.n74 VSS.n73 3.03311
R3229 VSS.n80 VSS.n79 3.03311
R3230 VSS.n89 VSS.n88 3.03311
R3231 VSS.n289 VSS.n288 3.03311
R3232 VSS.n29 VSS.n28 3.03311
R3233 VSS.n303 VSS.n302 3.03311
R3234 VSS.n313 VSS.n312 3.03311
R3235 VSS.n320 VSS.n319 3.03311
R3236 VSS.n329 VSS.n328 3.03311
R3237 VSS.n429 VSS.n428 3.03311
R3238 VSS.n22 VSS.n21 3.03311
R3239 VSS.n443 VSS.n442 3.03311
R3240 VSS.n453 VSS.n452 3.03311
R3241 VSS.n15 VSS.n14 3.03311
R3242 VSS.n501 VSS.n500 3.03311
R3243 VSS.n511 VSS.n510 3.03311
R3244 VSS.n571 VSS.n570 3.03311
R3245 VSS.n614 VSS.n613 3.03311
R3246 VSS.n666 VSS.n665 3.03311
R3247 VSS.n17 VSS.n16 2.56987
R3248 VSS.n24 VSS.n23 2.56987
R3249 VSS.n31 VSS.n30 2.56987
R3250 VSS.n688 VSS.n681 2.5605
R3251 VSS.n641 VSS.n640 2.24031
R3252 VSS.n689 VSS.n678 1.96973
R3253 VSS.n642 VSS 1.94963
R3254 VSS.n671 VSS.n670 1.35607
R3255 VSS.n695 VSS.n694 1.35607
R3256 VSS.n43 VSS.n42 1.35607
R3257 VSS.n72 VSS.n71 1.35607
R3258 VSS.n87 VSS.n86 1.35607
R3259 VSS.n311 VSS.n310 1.35607
R3260 VSS.n405 VSS.n404 1.35607
R3261 VSS.n327 VSS.n326 1.35607
R3262 VSS.n451 VSS.n450 1.35607
R3263 VSS.n487 VSS.n486 1.35607
R3264 VSS.n509 VSS.n508 1.35607
R3265 VSS.n555 VSS.n554 1.35607
R3266 VSS.n612 VSS.n611 1.35607
R3267 VSS.n709 VSS.n708 1.35607
R3268 VSS.n544 VSS.n543 1.13981
R3269 VSS.n302 VSS.n301 1.04008
R3270 VSS.n259 VSS.n258 1.04008
R3271 VSS.n442 VSS.n441 1.04008
R3272 VSS.n500 VSS.n499 1.04008
R3273 VSS.n158 VSS.n157 1.03985
R3274 VSS.n288 VSS.n286 1.03985
R3275 VSS.n201 VSS.n200 1.03985
R3276 VSS.n428 VSS.n426 1.03985
R3277 VSS.n498 VSS.n497 0.853
R3278 VSS.n536 VSS.n534 0.853
R3279 VSS.n497 VSS.n496 0.853
R3280 VSS.n554 VSS.n553 0.853
R3281 VSS.n553 VSS.n552 0.853
R3282 VSS.n492 VSS.n487 0.853
R3283 VSS.n424 VSS.n423 0.853
R3284 VSS.n425 VSS.n424 0.853
R3285 VSS.n389 VSS.n388 0.853
R3286 VSS.n493 VSS.n492 0.853
R3287 VSS.n410 VSS.n405 0.853
R3288 VSS.n219 VSS.n218 0.853
R3289 VSS.n218 VSS.n217 0.853
R3290 VSS.n262 VSS.n261 0.853
R3291 VSS.n261 VSS.n260 0.853
R3292 VSS.n284 VSS.n283 0.853
R3293 VSS.n285 VSS.n284 0.853
R3294 VSS.n150 VSS.n149 0.853
R3295 VSS.n411 VSS.n410 0.853
R3296 VSS.n644 VSS.n642 0.853
R3297 VSS.n645 VSS.n644 0.853
R3298 VSS.n610 VSS.n609 0.853
R3299 VSS.n167 VSS.n166 0.853
R3300 VSS.n168 VSS.n167 0.853
R3301 VSS.n611 VSS.n610 0.853
R3302 VSS.n697 VSS.n695 0.853
R3303 VSS.n708 VSS.n707 0.853
R3304 VSS.t8 VSS.t0 0.824007
R3305 VSS.n677 VSS.n676 0.788192
R3306 VSS.n689 VSS.n688 0.788192
R3307 VSS.n681 VSS.n680 0.788192
R3308 VSS.n650 VSS.n649 0.699777
R3309 VSS.n538 VSS.n537 0.698382
R3310 VSS.n543 VSS.n542 0.684595
R3311 VSS.n678 VSS.n677 0.591269
R3312 VSS.n539 VSS.n538 0.352759
R3313 VSS.n559 VSS.n315 0.341248
R3314 VSS.n559 VSS.n455 0.341248
R3315 VSS.n559 VSS.n558 0.341248
R3316 VSS.n559 VSS.n46 0.33661
R3317 VSS.n559 VSS.n60 0.33661
R3318 VSS.n559 VSS.n90 0.33661
R3319 VSS.n559 VSS.n330 0.33661
R3320 VSS.n560 VSS.n559 0.336142
R3321 VSS.n559 VSS.n53 0.336142
R3322 VSS.n559 VSS.n75 0.336142
R3323 VSS.n559 VSS.n290 0.336142
R3324 VSS.n559 VSS.n430 0.336142
R3325 VSS.n546 VSS.n545 0.280638
R3326 VSS.n147 VSS.n146 0.212
R3327 VSS.n386 VSS.n385 0.212
R3328 VSS.n665 VSS.n664 0.197423
R3329 VSS VSS.n6 0.177439
R3330 VSS.n648 VSS.n647 0.17525
R3331 VSS VSS.n494 0.148517
R3332 VSS VSS.n412 0.147312
R3333 VSS VSS.n169 0.147312
R3334 VSS.n647 VSS.n646 0.129277
R3335 VSS.n495 VSS 0.111158
R3336 VSS VSS.n390 0.111158
R3337 VSS.n413 VSS 0.111158
R3338 VSS VSS.n151 0.111158
R3339 VSS.n273 VSS 0.111158
R3340 VSS.n221 VSS 0.111158
R3341 VSS.n170 VSS 0.111158
R3342 VSS.n608 VSS 0.111158
R3343 VSS.n639 VSS 0.104812
R3344 VSS.n655 VSS.n654 0.0929479
R3345 VSS.n693 VSS.n692 0.0734167
R3346 VSS.n391 VSS 0.0718924
R3347 VSS.n152 VSS 0.0718924
R3348 VSS VSS.n272 0.0718924
R3349 VSS VSS.n220 0.0718924
R3350 VSS.n403 VSS.n402 0.0685147
R3351 VSS.n306 VSS.n305 0.0685147
R3352 VSS.n26 VSS.n25 0.0685147
R3353 VSS.n485 VSS.n484 0.0685147
R3354 VSS.n446 VSS.n445 0.0685147
R3355 VSS.n19 VSS.n18 0.0685147
R3356 VSS.n514 VSS.n513 0.0685147
R3357 VSS.n504 VSS.n503 0.0685147
R3358 VSS.n12 VSS.n11 0.0685147
R3359 VSS.n156 VSS.n155 0.0685147
R3360 VSS.n565 VSS.n564 0.0685147
R3361 VSS.n573 VSS.n572 0.0685147
R3362 VSS.n654 VSS.n0 0.0643021
R3363 VSS.n673 VSS 0.0512812
R3364 VSS.n649 VSS.n648 0.0498797
R3365 VSS.n163 VSS.n162 0.0482941
R3366 VSS.n576 VSS.n575 0.0482941
R3367 VSS.n582 VSS.n581 0.0482941
R3368 VSS.n398 VSS.n397 0.0482941
R3369 VSS.n297 VSS.n296 0.0482941
R3370 VSS.n109 VSS.n108 0.0482941
R3371 VSS.n103 VSS.n102 0.0482941
R3372 VSS.n247 VSS.n246 0.0482941
R3373 VSS.n253 VSS.n252 0.0482941
R3374 VSS.n214 VSS.n213 0.0482941
R3375 VSS.n208 VSS.n207 0.0482941
R3376 VSS.n480 VSS.n479 0.0482941
R3377 VSS.n437 VSS.n436 0.0482941
R3378 VSS.n349 VSS.n348 0.0482941
R3379 VSS.n343 VSS.n342 0.0482941
R3380 VSS.n518 VSS.n517 0.0482941
R3381 VSS.n462 VSS.n461 0.0482941
R3382 VSS.n708 VSS.n1 0.0427297
R3383 VSS.n534 VSS.n530 0.0415156
R3384 VSS.n642 VSS.n8 0.0415156
R3385 VSS.n705 VSS.n704 0.0411354
R3386 VSS.n165 VSS.n164 0.0391029
R3387 VSS.n161 VSS.n160 0.0391029
R3388 VSS.n578 VSS.n577 0.0391029
R3389 VSS.n580 VSS.n579 0.0391029
R3390 VSS.n611 VSS.n583 0.0391029
R3391 VSS.n404 VSS.n403 0.0391029
R3392 VSS.n311 VSS.n306 0.0391029
R3393 VSS.n27 VSS.n26 0.0391029
R3394 VSS.n405 VSS.n399 0.0391029
R3395 VSS.n310 VSS.n309 0.0391029
R3396 VSS.n293 VSS.n292 0.0391029
R3397 VSS.n295 VSS.n294 0.0391029
R3398 VSS.n299 VSS.n298 0.0391029
R3399 VSS.n288 VSS.n287 0.0391029
R3400 VSS.n92 VSS.n91 0.0391029
R3401 VSS.n94 VSS.n93 0.0391029
R3402 VSS.n77 VSS.n76 0.0391029
R3403 VSS.n79 VSS.n78 0.0391029
R3404 VSS.n87 VSS.n82 0.0391029
R3405 VSS.n111 VSS.n110 0.0391029
R3406 VSS.n107 VSS.n106 0.0391029
R3407 VSS.n105 VSS.n104 0.0391029
R3408 VSS.n101 VSS.n100 0.0391029
R3409 VSS.n99 VSS.n98 0.0391029
R3410 VSS.n86 VSS.n84 0.0391029
R3411 VSS.n72 VSS.n67 0.0391029
R3412 VSS.n64 VSS.n61 0.0391029
R3413 VSS.n63 VSS.n62 0.0391029
R3414 VSS.n57 VSS.n54 0.0391029
R3415 VSS.n56 VSS.n55 0.0391029
R3416 VSS.n258 VSS.n256 0.0391029
R3417 VSS.n71 VSS.n70 0.0391029
R3418 VSS.n243 VSS.n242 0.0391029
R3419 VSS.n245 VSS.n244 0.0391029
R3420 VSS.n249 VSS.n248 0.0391029
R3421 VSS.n251 VSS.n250 0.0391029
R3422 VSS.n255 VSS.n254 0.0391029
R3423 VSS.n200 VSS.n198 0.0391029
R3424 VSS.n48 VSS.n47 0.0391029
R3425 VSS.n50 VSS.n49 0.0391029
R3426 VSS.n33 VSS.n32 0.0391029
R3427 VSS.n35 VSS.n34 0.0391029
R3428 VSS.n43 VSS.n38 0.0391029
R3429 VSS.n216 VSS.n215 0.0391029
R3430 VSS.n212 VSS.n211 0.0391029
R3431 VSS.n210 VSS.n209 0.0391029
R3432 VSS.n206 VSS.n205 0.0391029
R3433 VSS.n204 VSS.n203 0.0391029
R3434 VSS.n42 VSS.n40 0.0391029
R3435 VSS.n486 VSS.n485 0.0391029
R3436 VSS.n451 VSS.n446 0.0391029
R3437 VSS.n20 VSS.n19 0.0391029
R3438 VSS.n487 VSS.n481 0.0391029
R3439 VSS.n450 VSS.n449 0.0391029
R3440 VSS.n433 VSS.n432 0.0391029
R3441 VSS.n435 VSS.n434 0.0391029
R3442 VSS.n439 VSS.n438 0.0391029
R3443 VSS.n428 VSS.n427 0.0391029
R3444 VSS.n332 VSS.n331 0.0391029
R3445 VSS.n334 VSS.n333 0.0391029
R3446 VSS.n317 VSS.n316 0.0391029
R3447 VSS.n319 VSS.n318 0.0391029
R3448 VSS.n327 VSS.n322 0.0391029
R3449 VSS.n351 VSS.n350 0.0391029
R3450 VSS.n347 VSS.n346 0.0391029
R3451 VSS.n345 VSS.n344 0.0391029
R3452 VSS.n341 VSS.n340 0.0391029
R3453 VSS.n339 VSS.n338 0.0391029
R3454 VSS.n326 VSS.n324 0.0391029
R3455 VSS.n555 VSS.n514 0.0391029
R3456 VSS.n509 VSS.n504 0.0391029
R3457 VSS.n13 VSS.n12 0.0391029
R3458 VSS.n554 VSS.n519 0.0391029
R3459 VSS.n508 VSS.n507 0.0391029
R3460 VSS.n458 VSS.n457 0.0391029
R3461 VSS.n460 VSS.n459 0.0391029
R3462 VSS.n464 VSS.n463 0.0391029
R3463 VSS.n157 VSS.n156 0.0391029
R3464 VSS.n155 VSS.n10 0.0391029
R3465 VSS.n564 VSS.n563 0.0391029
R3466 VSS.n566 VSS.n565 0.0391029
R3467 VSS.n572 VSS.n571 0.0391029
R3468 VSS.n612 VSS.n573 0.0391029
R3469 VSS.n4 VSS.n3 0.0361962
R3470 VSS.n668 VSS.n667 0.035973
R3471 VSS.n670 VSS.n669 0.035973
R3472 VSS VSS.n709 0.0330521
R3473 VSS.n695 VSS.n651 0.0325946
R3474 VSS VSS.n672 0.03175
R3475 VSS.n700 VSS.n699 0.029875
R3476 VSS.n672 VSS.n671 0.0278438
R3477 VSS.n640 VSS.n639 0.0257686
R3478 VSS.n532 VSS.n531 0.024008
R3479 VSS.n692 VSS 0.0226354
R3480 VSS.n642 VSS.n641 0.0223823
R3481 VSS.n611 VSS.n584 0.0219755
R3482 VSS.n405 VSS.n395 0.0219755
R3483 VSS.n86 VSS.n85 0.0219755
R3484 VSS.n71 VSS.n68 0.0219755
R3485 VSS.n42 VSS.n41 0.0219755
R3486 VSS.n487 VSS.n477 0.0219755
R3487 VSS.n326 VSS.n325 0.0219755
R3488 VSS.n554 VSS.n515 0.0219755
R3489 VSS.n666 VSS.n656 0.0213333
R3490 VSS.n694 VSS.n691 0.0200312
R3491 VSS.n410 VSS.n394 0.0191618
R3492 VSS.n410 VSS.n409 0.0191618
R3493 VSS.n137 VSS.n136 0.0191618
R3494 VSS.n141 VSS.n140 0.0191618
R3495 VSS.n142 VSS.n141 0.0191618
R3496 VSS.n149 VSS.n145 0.0191618
R3497 VSS.n149 VSS.n148 0.0191618
R3498 VSS.n284 VSS.n112 0.0191618
R3499 VSS.n284 VSS.n129 0.0191618
R3500 VSS.n126 VSS.n125 0.0191618
R3501 VSS.n125 VSS.n124 0.0191618
R3502 VSS.n121 VSS.n120 0.0191618
R3503 VSS.n120 VSS.n119 0.0191618
R3504 VSS.n116 VSS.n115 0.0191618
R3505 VSS.n115 VSS.n114 0.0191618
R3506 VSS.n224 VSS.n223 0.0191618
R3507 VSS.n225 VSS.n224 0.0191618
R3508 VSS.n229 VSS.n228 0.0191618
R3509 VSS.n230 VSS.n229 0.0191618
R3510 VSS.n234 VSS.n233 0.0191618
R3511 VSS.n235 VSS.n234 0.0191618
R3512 VSS.n261 VSS.n238 0.0191618
R3513 VSS.n261 VSS.n240 0.0191618
R3514 VSS.n218 VSS.n181 0.0191618
R3515 VSS.n218 VSS.n197 0.0191618
R3516 VSS.n194 VSS.n193 0.0191618
R3517 VSS.n193 VSS.n192 0.0191618
R3518 VSS.n189 VSS.n188 0.0191618
R3519 VSS.n188 VSS.n187 0.0191618
R3520 VSS.n184 VSS.n183 0.0191618
R3521 VSS.n183 VSS.n182 0.0191618
R3522 VSS.n492 VSS.n476 0.0191618
R3523 VSS.n492 VSS.n491 0.0191618
R3524 VSS.n376 VSS.n375 0.0191618
R3525 VSS.n380 VSS.n379 0.0191618
R3526 VSS.n381 VSS.n380 0.0191618
R3527 VSS.n388 VSS.n384 0.0191618
R3528 VSS.n388 VSS.n387 0.0191618
R3529 VSS.n424 VSS.n352 0.0191618
R3530 VSS.n424 VSS.n368 0.0191618
R3531 VSS.n365 VSS.n364 0.0191618
R3532 VSS.n364 VSS.n363 0.0191618
R3533 VSS.n360 VSS.n359 0.0191618
R3534 VSS.n359 VSS.n358 0.0191618
R3535 VSS.n355 VSS.n354 0.0191618
R3536 VSS.n354 VSS.n353 0.0191618
R3537 VSS.n553 VSS.n520 0.0191618
R3538 VSS.n553 VSS.n529 0.0191618
R3539 VSS.n526 VSS.n525 0.0191618
R3540 VSS.n525 VSS.n524 0.0191618
R3541 VSS.n466 VSS.n465 0.0191618
R3542 VSS.n497 VSS.n469 0.0191618
R3543 VSS.n497 VSS.n470 0.0191618
R3544 VSS.n167 VSS.n153 0.0191618
R3545 VSS.n589 VSS.n588 0.0191618
R3546 VSS.n590 VSS.n589 0.0191618
R3547 VSS.n594 VSS.n593 0.0191618
R3548 VSS.n595 VSS.n594 0.0191618
R3549 VSS.n610 VSS.n598 0.0191618
R3550 VSS.n610 VSS.n599 0.0191618
R3551 VSS.n552 VSS.n546 0.0183481
R3552 VSS.n552 VSS.n551 0.0183481
R3553 VSS.n550 VSS.n549 0.0183481
R3554 VSS.n549 VSS.n548 0.0183481
R3555 VSS.n472 VSS.n471 0.0183481
R3556 VSS.n496 VSS.n473 0.0183481
R3557 VSS.n496 VSS.n495 0.0183481
R3558 VSS.n494 VSS.n493 0.0183481
R3559 VSS.n493 VSS.n475 0.0183481
R3560 VSS.n370 VSS.n369 0.0183481
R3561 VSS.n372 VSS.n371 0.0183481
R3562 VSS.n373 VSS.n372 0.0183481
R3563 VSS.n389 VSS.n374 0.0183481
R3564 VSS.n390 VSS.n389 0.0183481
R3565 VSS.n423 VSS.n391 0.0183481
R3566 VSS.n423 VSS.n422 0.0183481
R3567 VSS.n421 VSS.n420 0.0183481
R3568 VSS.n420 VSS.n419 0.0183481
R3569 VSS.n418 VSS.n417 0.0183481
R3570 VSS.n417 VSS.n416 0.0183481
R3571 VSS.n415 VSS.n414 0.0183481
R3572 VSS.n414 VSS.n413 0.0183481
R3573 VSS.n412 VSS.n411 0.0183481
R3574 VSS.n411 VSS.n393 0.0183481
R3575 VSS.n131 VSS.n130 0.0183481
R3576 VSS.n133 VSS.n132 0.0183481
R3577 VSS.n134 VSS.n133 0.0183481
R3578 VSS.n150 VSS.n135 0.0183481
R3579 VSS.n151 VSS.n150 0.0183481
R3580 VSS.n283 VSS.n152 0.0183481
R3581 VSS.n283 VSS.n282 0.0183481
R3582 VSS.n281 VSS.n280 0.0183481
R3583 VSS.n280 VSS.n279 0.0183481
R3584 VSS.n278 VSS.n277 0.0183481
R3585 VSS.n277 VSS.n276 0.0183481
R3586 VSS.n275 VSS.n274 0.0183481
R3587 VSS.n274 VSS.n273 0.0183481
R3588 VSS.n272 VSS.n271 0.0183481
R3589 VSS.n271 VSS.n270 0.0183481
R3590 VSS.n269 VSS.n268 0.0183481
R3591 VSS.n268 VSS.n267 0.0183481
R3592 VSS.n266 VSS.n265 0.0183481
R3593 VSS.n265 VSS.n264 0.0183481
R3594 VSS.n263 VSS.n262 0.0183481
R3595 VSS.n262 VSS.n221 0.0183481
R3596 VSS.n220 VSS.n219 0.0183481
R3597 VSS.n219 VSS.n179 0.0183481
R3598 VSS.n178 VSS.n177 0.0183481
R3599 VSS.n177 VSS.n176 0.0183481
R3600 VSS.n175 VSS.n174 0.0183481
R3601 VSS.n174 VSS.n173 0.0183481
R3602 VSS.n172 VSS.n171 0.0183481
R3603 VSS.n171 VSS.n170 0.0183481
R3604 VSS.n169 VSS.n168 0.0183481
R3605 VSS.n602 VSS.n601 0.0183481
R3606 VSS.n603 VSS.n602 0.0183481
R3607 VSS.n605 VSS.n604 0.0183481
R3608 VSS.n606 VSS.n605 0.0183481
R3609 VSS.n609 VSS.n607 0.0183481
R3610 VSS.n609 VSS.n608 0.0183481
R3611 VSS.n648 VSS.n5 0.0183481
R3612 VSS.n5 VSS.n4 0.0183481
R3613 VSS.n645 VSS.n6 0.0172857
R3614 VSS.n646 VSS.n645 0.0172857
R3615 VSS.n541 VSS.n540 0.0156071
R3616 VSS.n536 VSS.n535 0.0156071
R3617 VSS.n644 VSS.n7 0.0156071
R3618 VSS.n644 VSS.n643 0.0156071
R3619 VSS.n408 VSS.n407 0.0143235
R3620 VSS.n139 VSS.n138 0.0143235
R3621 VSS.n144 VSS.n143 0.0143235
R3622 VSS.n128 VSS.n127 0.0143235
R3623 VSS.n123 VSS.n122 0.0143235
R3624 VSS.n118 VSS.n117 0.0143235
R3625 VSS.n227 VSS.n226 0.0143235
R3626 VSS.n232 VSS.n231 0.0143235
R3627 VSS.n237 VSS.n236 0.0143235
R3628 VSS.n196 VSS.n195 0.0143235
R3629 VSS.n191 VSS.n190 0.0143235
R3630 VSS.n186 VSS.n185 0.0143235
R3631 VSS.n490 VSS.n489 0.0143235
R3632 VSS.n378 VSS.n377 0.0143235
R3633 VSS.n383 VSS.n382 0.0143235
R3634 VSS.n367 VSS.n366 0.0143235
R3635 VSS.n362 VSS.n361 0.0143235
R3636 VSS.n357 VSS.n356 0.0143235
R3637 VSS.n528 VSS.n527 0.0143235
R3638 VSS.n523 VSS.n522 0.0143235
R3639 VSS.n468 VSS.n467 0.0143235
R3640 VSS.n587 VSS.n586 0.0143235
R3641 VSS.n592 VSS.n591 0.0143235
R3642 VSS.n597 VSS.n596 0.0143235
R3643 VSS.n639 VSS.n638 0.0142993
R3644 VSS.n533 VSS.n532 0.0137243
R3645 VSS.n707 VSS.n706 0.0137188
R3646 VSS.n703 VSS.n702 0.0137188
R3647 VSS.n702 VSS.n701 0.0137188
R3648 VSS.n698 VSS.n697 0.0137188
R3649 VSS.n690 VSS.n675 0.0135208
R3650 VSS.n551 VSS.n550 0.0123987
R3651 VSS.n548 VSS.n547 0.0123987
R3652 VSS.n473 VSS.n472 0.0123987
R3653 VSS.n475 VSS.n474 0.0123987
R3654 VSS.n371 VSS.n370 0.0123987
R3655 VSS.n374 VSS.n373 0.0123987
R3656 VSS.n422 VSS.n421 0.0123987
R3657 VSS.n419 VSS.n418 0.0123987
R3658 VSS.n416 VSS.n415 0.0123987
R3659 VSS.n393 VSS.n392 0.0123987
R3660 VSS.n132 VSS.n131 0.0123987
R3661 VSS.n135 VSS.n134 0.0123987
R3662 VSS.n282 VSS.n281 0.0123987
R3663 VSS.n279 VSS.n278 0.0123987
R3664 VSS.n276 VSS.n275 0.0123987
R3665 VSS.n270 VSS.n269 0.0123987
R3666 VSS.n267 VSS.n266 0.0123987
R3667 VSS.n264 VSS.n263 0.0123987
R3668 VSS.n179 VSS.n178 0.0123987
R3669 VSS.n176 VSS.n175 0.0123987
R3670 VSS.n173 VSS.n172 0.0123987
R3671 VSS.n601 VSS.n600 0.0123987
R3672 VSS.n604 VSS.n603 0.0123987
R3673 VSS.n607 VSS.n606 0.0123987
R3674 VSS.n695 VSS.n652 0.0123243
R3675 VSS.n640 VSS 0.0121822
R3676 VSS.n162 VSS.n161 0.0115294
R3677 VSS.n577 VSS.n576 0.0115294
R3678 VSS.n583 VSS.n582 0.0115294
R3679 VSS.n399 VSS.n398 0.0115294
R3680 VSS.n309 VSS.n308 0.0115294
R3681 VSS.n296 VSS.n295 0.0115294
R3682 VSS.n108 VSS.n107 0.0115294
R3683 VSS.n102 VSS.n101 0.0115294
R3684 VSS.n84 VSS.n83 0.0115294
R3685 VSS.n70 VSS.n69 0.0115294
R3686 VSS.n246 VSS.n245 0.0115294
R3687 VSS.n252 VSS.n251 0.0115294
R3688 VSS.n213 VSS.n212 0.0115294
R3689 VSS.n207 VSS.n206 0.0115294
R3690 VSS.n40 VSS.n39 0.0115294
R3691 VSS.n481 VSS.n480 0.0115294
R3692 VSS.n449 VSS.n448 0.0115294
R3693 VSS.n436 VSS.n435 0.0115294
R3694 VSS.n348 VSS.n347 0.0115294
R3695 VSS.n342 VSS.n341 0.0115294
R3696 VSS.n324 VSS.n323 0.0115294
R3697 VSS.n519 VSS.n518 0.0115294
R3698 VSS.n507 VSS.n506 0.0115294
R3699 VSS.n461 VSS.n460 0.0115294
R3700 VSS.n301 VSS.n300 0.0104679
R3701 VSS.n260 VSS.n259 0.0104679
R3702 VSS.n441 VSS.n440 0.0104679
R3703 VSS.n499 VSS.n498 0.0104679
R3704 VSS.n166 VSS.n158 0.0098203
R3705 VSS.n217 VSS.n201 0.0098203
R3706 VSS.n286 VSS.n285 0.0098203
R3707 VSS.n426 VSS.n425 0.0098203
R3708 VSS.n164 VSS.n163 0.00969118
R3709 VSS.n575 VSS.n574 0.00969118
R3710 VSS.n581 VSS.n580 0.00969118
R3711 VSS.n397 VSS.n396 0.00969118
R3712 VSS.n292 VSS.n291 0.00969118
R3713 VSS.n298 VSS.n297 0.00969118
R3714 VSS.n110 VSS.n109 0.00969118
R3715 VSS.n104 VSS.n103 0.00969118
R3716 VSS.n98 VSS.n97 0.00969118
R3717 VSS.n242 VSS.n241 0.00969118
R3718 VSS.n248 VSS.n247 0.00969118
R3719 VSS.n254 VSS.n253 0.00969118
R3720 VSS.n215 VSS.n214 0.00969118
R3721 VSS.n209 VSS.n208 0.00969118
R3722 VSS.n203 VSS.n202 0.00969118
R3723 VSS.n479 VSS.n478 0.00969118
R3724 VSS.n432 VSS.n431 0.00969118
R3725 VSS.n438 VSS.n437 0.00969118
R3726 VSS.n350 VSS.n349 0.00969118
R3727 VSS.n344 VSS.n343 0.00969118
R3728 VSS.n338 VSS.n337 0.00969118
R3729 VSS.n517 VSS.n516 0.00969118
R3730 VSS.n457 VSS.n456 0.00969118
R3731 VSS.n463 VSS.n462 0.00969118
R3732 VSS.n694 VSS.n693 0.00961458
R3733 VSS.n656 VSS.n655 0.00701042
R3734 VSS.n674 VSS.n673 0.00570833
R3735 VSS.n691 VSS.n690 0.00570833
R3736 VSS.n647 VSS 0.005375
R3737 VSS.n544 VSS.n539 0.00493396
R3738 VSS.n545 VSS.n544 0.00493396
R3739 VSS.n537 VSS.n536 0.00489326
R3740 VSS.n707 VSS.n650 0.00451955
R3741 VSS.n675 VSS.n674 0.00440625
R3742 VSS.n697 VSS.n696 0.00362372
R3743 VSS.n409 VSS.n408 0.00257353
R3744 VSS.n407 VSS.n406 0.00257353
R3745 VSS.n138 VSS.n137 0.00257353
R3746 VSS.n140 VSS.n139 0.00257353
R3747 VSS.n143 VSS.n142 0.00257353
R3748 VSS.n145 VSS.n144 0.00257353
R3749 VSS.n148 VSS.n147 0.00257353
R3750 VSS.n146 VSS.n112 0.00257353
R3751 VSS.n129 VSS.n128 0.00257353
R3752 VSS.n127 VSS.n126 0.00257353
R3753 VSS.n124 VSS.n123 0.00257353
R3754 VSS.n122 VSS.n121 0.00257353
R3755 VSS.n119 VSS.n118 0.00257353
R3756 VSS.n117 VSS.n116 0.00257353
R3757 VSS.n114 VSS.n113 0.00257353
R3758 VSS.n223 VSS.n222 0.00257353
R3759 VSS.n226 VSS.n225 0.00257353
R3760 VSS.n228 VSS.n227 0.00257353
R3761 VSS.n231 VSS.n230 0.00257353
R3762 VSS.n233 VSS.n232 0.00257353
R3763 VSS.n236 VSS.n235 0.00257353
R3764 VSS.n238 VSS.n237 0.00257353
R3765 VSS.n240 VSS.n239 0.00257353
R3766 VSS.n181 VSS.n180 0.00257353
R3767 VSS.n197 VSS.n196 0.00257353
R3768 VSS.n195 VSS.n194 0.00257353
R3769 VSS.n192 VSS.n191 0.00257353
R3770 VSS.n190 VSS.n189 0.00257353
R3771 VSS.n187 VSS.n186 0.00257353
R3772 VSS.n185 VSS.n184 0.00257353
R3773 VSS.n491 VSS.n490 0.00257353
R3774 VSS.n489 VSS.n488 0.00257353
R3775 VSS.n377 VSS.n376 0.00257353
R3776 VSS.n379 VSS.n378 0.00257353
R3777 VSS.n382 VSS.n381 0.00257353
R3778 VSS.n384 VSS.n383 0.00257353
R3779 VSS.n387 VSS.n386 0.00257353
R3780 VSS.n385 VSS.n352 0.00257353
R3781 VSS.n368 VSS.n367 0.00257353
R3782 VSS.n366 VSS.n365 0.00257353
R3783 VSS.n363 VSS.n362 0.00257353
R3784 VSS.n361 VSS.n360 0.00257353
R3785 VSS.n358 VSS.n357 0.00257353
R3786 VSS.n356 VSS.n355 0.00257353
R3787 VSS.n529 VSS.n528 0.00257353
R3788 VSS.n527 VSS.n526 0.00257353
R3789 VSS.n524 VSS.n523 0.00257353
R3790 VSS.n522 VSS.n521 0.00257353
R3791 VSS.n467 VSS.n466 0.00257353
R3792 VSS.n469 VSS.n468 0.00257353
R3793 VSS.n586 VSS.n585 0.00257353
R3794 VSS.n588 VSS.n587 0.00257353
R3795 VSS.n591 VSS.n590 0.00257353
R3796 VSS.n593 VSS.n592 0.00257353
R3797 VSS.n596 VSS.n595 0.00257353
R3798 VSS.n598 VSS.n597 0.00257353
R3799 VSS.n166 VSS.n165 0.00233824
R3800 VSS.n160 VSS.n159 0.00233824
R3801 VSS.n579 VSS.n578 0.00233824
R3802 VSS.n404 VSS.n401 0.00233824
R3803 VSS.n312 VSS.n311 0.00233824
R3804 VSS.n28 VSS.n27 0.00233824
R3805 VSS.n310 VSS.n307 0.00233824
R3806 VSS.n294 VSS.n293 0.00233824
R3807 VSS.n300 VSS.n299 0.00233824
R3808 VSS.n94 VSS.n92 0.00233824
R3809 VSS.n79 VSS.n77 0.00233824
R3810 VSS.n88 VSS.n87 0.00233824
R3811 VSS.n285 VSS.n111 0.00233824
R3812 VSS.n106 VSS.n105 0.00233824
R3813 VSS.n100 VSS.n99 0.00233824
R3814 VSS.n73 VSS.n72 0.00233824
R3815 VSS.n64 VSS.n63 0.00233824
R3816 VSS.n57 VSS.n56 0.00233824
R3817 VSS.n244 VSS.n243 0.00233824
R3818 VSS.n250 VSS.n249 0.00233824
R3819 VSS.n260 VSS.n255 0.00233824
R3820 VSS.n50 VSS.n48 0.00233824
R3821 VSS.n35 VSS.n33 0.00233824
R3822 VSS.n44 VSS.n43 0.00233824
R3823 VSS.n217 VSS.n216 0.00233824
R3824 VSS.n211 VSS.n210 0.00233824
R3825 VSS.n205 VSS.n204 0.00233824
R3826 VSS.n486 VSS.n483 0.00233824
R3827 VSS.n452 VSS.n451 0.00233824
R3828 VSS.n21 VSS.n20 0.00233824
R3829 VSS.n450 VSS.n447 0.00233824
R3830 VSS.n434 VSS.n433 0.00233824
R3831 VSS.n440 VSS.n439 0.00233824
R3832 VSS.n334 VSS.n332 0.00233824
R3833 VSS.n319 VSS.n317 0.00233824
R3834 VSS.n328 VSS.n327 0.00233824
R3835 VSS.n425 VSS.n351 0.00233824
R3836 VSS.n346 VSS.n345 0.00233824
R3837 VSS.n340 VSS.n339 0.00233824
R3838 VSS.n556 VSS.n555 0.00233824
R3839 VSS.n510 VSS.n509 0.00233824
R3840 VSS.n14 VSS.n13 0.00233824
R3841 VSS.n508 VSS.n505 0.00233824
R3842 VSS.n459 VSS.n458 0.00233824
R3843 VSS.n498 VSS.n464 0.00233824
R3844 VSS.n563 VSS.n10 0.00233824
R3845 VSS.n571 VSS.n566 0.00233824
R3846 VSS.n613 VSS.n612 0.00233824
R3847 VSS.n670 VSS.n668 0.00218919
R3848 VSS.n708 VSS.n2 0.00218919
R3849 VSS.n543 VSS.n541 0.0021514
R3850 VSS.n706 VSS.n705 0.00196875
R3851 VSS.n704 VSS.n703 0.00196875
R3852 VSS.n701 VSS.n700 0.00196875
R3853 VSS.n699 VSS.n698 0.00196875
R3854 VSS.n709 VSS.n0 0.00180208
R3855 VSS.n671 VSS.n666 0.00180208
R3856 VSS.n534 VSS.n533 0.0011215
R3857 code_offset.n2 code_offset.t1 230.016
R3858 code_offset.n1 code_offset.t2 153.665
R3859 code_offset.n2 code_offset 153.601
R3860 code_offset code_offset.t0 140.379
R3861 code_offset.n3 code_offset.n2 9.3005
R3862 code_offset.n2 code_offset.n1 4.91671
R3863 code_offset.n5 code_offset.n3 4.9013
R3864 code_offset.n4 code_offset 4.22092
R3865 code_offset code_offset.n0 2.4005
R3866 code_offset.n4 code_offset 1.01229
R3867 code_offset.n5 code_offset.n4 0.726043
R3868 code_offset.n3 code_offset.n0 0.533833
R3869 code_offset.n6 code_offset.n5 0.421696
R3870 code_offset code_offset.n6 0.0195217
R3871 code_offset.n6 code_offset 0.0170094
R3872 OUT.n2 OUT.t5 107.647
R3873 OUT.n1 OUT.t4 107.647
R3874 OUT.n2 OUT.t3 91.5805
R3875 OUT.n1 OUT.t2 91.5805
R3876 OUT.n0 OUT.t0 68.3658
R3877 OUT.n2 OUT.n1 58.5727
R3878 OUT.n0 OUT.t1 41.7552
R3879 OUT OUT.n2 13.4931
R3880 OUT OUT.n0 0.422914
R3881 code[1] code[1].t0 140.387
R3882 code[1].n0 code[1].t1 140.34
R3883 code[1].n0 code[1] 0.201587
R3884 code[1] code[1].n0 0.0371379
R3885 IN.t4 IN.t17 221.72
R3886 IN.t7 IN.t4 221.72
R3887 IN.t14 IN.t7 221.72
R3888 IN.t2 IN.t14 221.72
R3889 IN.t12 IN.t2 221.72
R3890 IN.t5 IN.t9 221.72
R3891 IN.t18 IN.t5 221.72
R3892 IN.t11 IN.t18 221.72
R3893 IN.t0 IN.t11 221.72
R3894 IN.t21 IN.t0 221.72
R3895 IN.t16 IN.t21 221.72
R3896 IN.t10 IN.t16 221.72
R3897 IN.t1 IN.t6 221.72
R3898 IN.t13 IN.t1 221.72
R3899 IN.t8 IN.t13 221.72
R3900 IN.t20 IN.t8 221.72
R3901 IN.t3 IN.t20 221.72
R3902 IN.t19 IN.t3 221.72
R3903 IN.t15 IN.t19 221.72
R3904 IN.n5 IN.t12 154.8
R3905 IN.n0 IN 89.9738
R3906 IN.n1 IN.t10 78.7272
R3907 IN.n0 IN.t15 74.6592
R3908 IN.n2 IN 40.1672
R3909 IN.n3 IN.n1 32.1338
R3910 IN IN.n1 21.4227
R3911 IN.n4 IN.n0 21.3547
R3912 IN.n4 IN.n3 17.8279
R3913 IN.n5 IN.n4 13.4163
R3914 IN.n2 IN 11.8854
R3915 IN.n3 IN.n2 3.96214
R3916 IN.n6 IN 1.64944
R3917 IN.n6 IN 0.10169
R3918 IN IN.n6 0.00215441
R3919 IN.n6 IN.n5 0.00197059
R3920 code[3].n0 code[3].t0 229.971
R3921 code[3].n0 code[3].t1 158.35
R3922 code[3].n1 code[3].n0 8.50845
R3923 code[3].n1 code[3] 3.95275
R3924 code[3].n2 code[3].n1 1.73287
R3925 code[3].n3 code[3] 0.474765
R3926 code[3] code[3].n3 0.366977
R3927 code[3].n2 code[3] 0.339042
R3928 code[3].n3 code[3].n2 0.00334091
R3929 code[0] code[0].t0 140.376
C0 nstack_lab5 x4[3].floating 1.17e-19
C1 a_9893_1017# x7.floating 8.52e-19
C2 OUT VDD 0.239f
C3 pstack_lab5 x5[7].floating 2.76e-19
C4 x6.SW x6.floating 0.13f
C5 nstack_lab1 a_9893_465# 0.00227f
C6 nstack_lab5 nstack_lab7 0.0316f
C7 OUT x10.Y 1.13e-19
C8 VDD a_15703_1681# 0.211f
C9 a_9893_1293# IN 0.00196f
C10 code_offset VDD 0.199f
C11 a_15703_1681# x10.Y 0.00127f
C12 code_offset x10.Y 0.0402f
C13 a_9893_1293# x7.floating 8.52e-19
C14 nstack_lab7 x4[3].floating 1.17e-19
C15 pstack_lab4 VDD 0.127f
C16 pstack_lab3 x5[7].floating 2.76e-19
C17 pstack_lab4 x10.Y 4.2e-19
C18 nstack_lab4 Uc 1.74e-19
C19 nstack_lab6 x6.floating 0.00278f
C20 nstack_lab5 a_9893_1017# 0.00227f
C21 x6.floating IN 0.0293f
C22 code[3] code_offset 0.0293f
C23 x3[1].floating x5[7].floating 0.8f
C24 Uc VDD 0.641f
C25 x7.floating x6.floating 0.202f
C26 IN pstack_lab2 0.00847f
C27 nstack_lab3 code_offset 5.57e-19
C28 Uc x10.Y 1.01f
C29 code_offset nstack_lab1 2.98e-19
C30 x6.SW x5[7].floating 0.00138f
C31 nstack_lab1 a_9893_327# 0.0022f
C32 VDD code[0] 0.00321f
C33 code[0] x10.Y 0.0124f
C34 pstack_lab5 VDD 0.106f
C35 x2.floating a_15703_1340# 0.0104f
C36 nstack_lab7 a_9893_1293# 0.00227f
C37 pstack_lab5 x10.Y 0.039f
C38 nstack_lab2 x6.floating 0.00109f
C39 code[1] x4[3].floating 0.00929f
C40 code[2] code_offset 0.00739f
C41 nstack_lab4 a_9893_741# 0.00227f
C42 code[1] x2.floating 0.0027f
C43 pstack_lab3 VDD 0.0324f
C44 x5[7].floating IN 0.00113f
C45 pstack_lab3 x10.Y 2.35e-19
C46 a_9893_879# IN 5.05e-19
C47 x7.floating x5[7].floating 0.182f
C48 code[3] pstack_lab5 2.69e-19
C49 code_offset a_9893_465# 2.1e-19
C50 a_9893_879# x7.floating 8.52e-19
C51 nstack_lab4 x6.SW 1.28e-19
C52 VDD x3[1].floating 0.0301f
C53 code[2] Uc 0.322f
C54 x3[1].floating x10.Y 0.00302f
C55 x6.SW VDD 0.423f
C56 x6.SW x10.Y 0.788f
C57 nstack_lab3 a_9893_741# 0.00227f
C58 code[1] a_15703_1340# 3.4e-20
C59 OUT a_15703_1681# 0.137f
C60 nstack_lab4 nstack_lab6 0.0316f
C61 a_9893_879# nstack_lab5 0.00227f
C62 x6.floating pstack_lab1 0.00578f
C63 nstack_lab4 IN 0.0135f
C64 x4[3].floating x5[7].floating 1.55f
C65 code_offset a_9893_327# 1.6e-19
C66 x6.SW code[3] 0.00466f
C67 x2.floating x5[7].floating 0.441f
C68 pstack_lab1 pstack_lab2 0.0704f
C69 nstack_lab4 x7.floating 0.0089f
C70 code_offset a_9893_1155# 7.9e-19
C71 VDD IN 0.335f
C72 nstack_lab3 x6.SW 4.74e-20
C73 code_offset pstack_lab4 3.64e-19
C74 x6.SW nstack_lab1 3.1e-20
C75 x10.Y IN 0.0967f
C76 VDD x7.floating 0.0282f
C77 x7.floating x10.Y 0.00345f
C78 code[2] x3[1].floating 0.00115f
C79 OUT Uc 0.127f
C80 nstack_lab3 a_9893_603# 0.00227f
C81 nstack_lab4 nstack_lab2 0.0316f
C82 Uc a_15703_1681# 0.00887f
C83 Uc code_offset 0.255f
C84 OUT code[0] 8.53e-20
C85 code[3] IN 0.00346f
C86 nstack_lab4 nstack_lab5 0.0388f
C87 x5[7].floating pstack_lab1 2.14e-19
C88 x6.floating pstack_lab2 0.0187f
C89 Uc pstack_lab4 0.032f
C90 nstack_lab3 IN 0.0136f
C91 nstack_lab1 IN 0.0127f
C92 nstack_lab3 x7.floating 0.00409f
C93 nstack_lab4 x4[3].floating 6.66e-19
C94 nstack_lab1 x7.floating 0.00218f
C95 nstack_lab5 x10.Y 6.65e-20
C96 code_offset pstack_lab5 0.00273f
C97 code[1] x5[7].floating 0.0022f
C98 pstack_lab4 pstack_lab5 0.0704f
C99 VDD x4[3].floating 0.0565f
C100 VDD x2.floating 0.0334f
C101 VDD nstack_lab7 0.00115f
C102 x4[3].floating x10.Y 0.00668f
C103 x2.floating x10.Y 0.00202f
C104 nstack_lab7 x10.Y 1.69e-19
C105 code_offset pstack_lab3 6.38e-19
C106 nstack_lab3 nstack_lab2 0.0388f
C107 code[2] x7.floating 0.0056f
C108 code_offset a_9893_741# 3.54e-19
C109 nstack_lab1 nstack_lab2 0.0388f
C110 Uc code[0] 0.0232f
C111 pstack_lab3 pstack_lab4 0.0704f
C112 x6.floating x5[7].floating 1.18f
C113 nstack_lab3 nstack_lab5 0.0316f
C114 x5[7].floating pstack_lab2 0.00138f
C115 Uc pstack_lab5 0.0702f
C116 a_9893_465# IN 1.8e-19
C117 nstack_lab3 x4[3].floating 1.17e-19
C118 a_9893_465# x7.floating 8.52e-19
C119 nstack_lab1 x4[3].floating 7.17e-20
C120 VDD pstack_lab1 0.109f
C121 x6.SW code_offset 0.19f
C122 x10.Y pstack_lab1 1.02e-19
C123 VDD a_15703_1340# 0.235f
C124 VDD a_9893_1293# 1.29e-19
C125 code[1] VDD 0.0181f
C126 code_offset a_9893_603# 2.7e-19
C127 code[2] x4[3].floating 0.518f
C128 a_9893_465# nstack_lab2 0.00227f
C129 code[1] x10.Y 6.64e-19
C130 pstack_lab3 pstack_lab5 0.0316f
C131 Uc x3[1].floating 0.341f
C132 nstack_lab4 x6.floating 0.00167f
C133 nstack_lab6 code_offset 0.00297f
C134 x6.SW Uc 0.164f
C135 code_offset IN 0.239f
C136 nstack_lab6 a_9893_1155# 0.00227f
C137 a_9893_327# IN 1.34e-19
C138 x3[1].floating code[0] 0.0326f
C139 VDD x6.floating 5.75f
C140 a_9893_1155# IN 0.0013f
C141 pstack_lab4 IN 0.00921f
C142 code_offset x7.floating 0.17f
C143 x6.floating x10.Y 0.087f
C144 VDD pstack_lab2 0.157f
C145 a_9893_1155# x7.floating 8.52e-19
C146 x10.Y pstack_lab2 1.49e-19
C147 x6.SW pstack_lab5 0.00707f
C148 nstack_lab6 Uc 0.032f
C149 code_offset nstack_lab2 3.98e-19
C150 Uc IN 0.37f
C151 code[3] x6.floating 0.00519f
C152 x6.SW pstack_lab3 9.98e-20
C153 Uc x7.floating 0.185f
C154 nstack_lab5 code_offset 0.0014f
C155 code[2] code[1] 0.00401f
C156 a_9893_879# nstack_lab4 0.00227f
C157 OUT x2.floating 0.0191f
C158 VDD x5[7].floating 43.9f
C159 pstack_lab5 IN 0.0175f
C160 code_offset x4[3].floating 0.00402f
C161 x5[7].floating x10.Y 1.01f
C162 code_offset nstack_lab7 0.0165f
C163 nstack_lab7 a_9893_1155# 0.00227f
C164 Uc nstack_lab2 8.05e-20
C165 pstack_lab3 IN 0.00866f
C166 a_9893_741# IN 3.4e-19
C167 a_9893_741# x7.floating 8.52e-19
C168 Uc x4[3].floating 0.636f
C169 a_9893_1017# code_offset 6.22e-19
C170 Uc x2.floating 0.193f
C171 Uc nstack_lab7 0.0388f
C172 OUT a_15703_1340# 0.141f
C173 code_offset pstack_lab1 3.28e-19
C174 code[0] x4[3].floating 2.28e-21
C175 nstack_lab6 x6.SW 2.44e-19
C176 x2.floating code[0] 0.161f
C177 x6.SW IN 0.0928f
C178 a_15703_1340# a_15703_1681# 0.0158f
C179 OUT code[1] 5.47e-22
C180 code_offset a_9893_1293# 9.08e-19
C181 x6.SW x7.floating 9.72e-19
C182 code[2] x5[7].floating 0.0056f
C183 VDD x10.Y 2.71f
C184 a_9893_603# IN 2.42e-19
C185 a_9893_603# x7.floating 8.52e-19
C186 nstack_lab6 IN 0.0135f
C187 x6.SW nstack_lab2 7.9e-20
C188 code_offset x6.floating 0.0624f
C189 nstack_lab4 nstack_lab3 0.0388f
C190 Uc a_15703_1340# 0.00892f
C191 Uc a_9893_1293# 0.00227f
C192 nstack_lab6 x7.floating 0.0089f
C193 pstack_lab4 x6.floating 0.0187f
C194 code[3] VDD 0.127f
C195 x7.floating IN 0.0241f
C196 code_offset pstack_lab2 1.9e-19
C197 nstack_lab5 x6.SW 8.11e-20
C198 code[1] Uc 0.0622f
C199 a_15703_1340# code[0] 0.00169f
C200 x3[1].floating x4[3].floating 1.19f
C201 code[3] x10.Y 0.0519f
C202 pstack_lab4 pstack_lab2 0.0316f
C203 a_9893_603# nstack_lab2 0.00227f
C204 x3[1].floating x2.floating 1.17f
C205 nstack_lab3 x10.Y 4.07e-20
C206 code[1] code[0] 0.0619f
C207 nstack_lab1 x10.Y 2.2e-20
C208 x6.SW nstack_lab7 0.00179f
C209 nstack_lab2 IN 0.0135f
C210 pstack_lab3 pstack_lab1 0.0316f
C211 Uc x6.floating 0.229f
C212 OUT x5[7].floating 0.0199f
C213 code[2] VDD 0.0372f
C214 nstack_lab6 nstack_lab5 0.0388f
C215 nstack_lab2 x7.floating 0.0089f
C216 Uc pstack_lab2 1.5e-19
C217 nstack_lab5 IN 0.0136f
C218 code[2] x10.Y 0.00201f
C219 a_15703_1681# x5[7].floating 0.0132f
C220 code_offset x5[7].floating 0.00308f
C221 a_9893_879# code_offset 4.7e-19
C222 nstack_lab5 x7.floating 0.00409f
C223 nstack_lab6 x4[3].floating 6.66e-19
C224 nstack_lab3 nstack_lab1 0.0316f
C225 pstack_lab5 x6.floating 0.00996f
C226 pstack_lab4 x5[7].floating 0.00138f
C227 x4[3].floating IN 6.65e-19
C228 nstack_lab6 nstack_lab7 0.0388f
C229 nstack_lab7 IN 0.0217f
C230 x6.SW pstack_lab1 5.11e-20
C231 x7.floating x4[3].floating 1.18f
C232 x3[1].floating a_15703_1340# 3.09e-19
C233 nstack_lab7 x7.floating 0.00409f
C234 pstack_lab3 x6.floating 0.00996f
C235 code[1] x3[1].floating 0.219f
C236 Uc x5[7].floating 1.19f
C237 pstack_lab3 pstack_lab2 0.0704f
C238 nstack_lab6 a_9893_1017# 0.00227f
C239 nstack_lab2 x4[3].floating 6.66e-19
C240 code[0] x5[7].floating 0.00119f
C241 a_9893_1017# IN 7.93e-19
C242 nstack_lab4 code_offset 8.34e-19
C243 IN pstack_lab1 0.00832f
C244 OUT VSS 0.422f
C245 a_9893_327# VSS 0.00426f
C246 a_9893_465# VSS 9.21e-19
C247 nstack_lab1 VSS 0.177f
C248 nstack_lab2 VSS 0.177f
C249 a_9893_603# VSS 8.65e-19
C250 a_9893_741# VSS 8.09e-19
C251 nstack_lab3 VSS 0.114f
C252 nstack_lab4 VSS 0.138f
C253 a_9893_879# VSS 7.57e-19
C254 a_9893_1017# VSS 7.1e-19
C255 nstack_lab5 VSS 0.114f
C256 nstack_lab6 VSS 0.143f
C257 a_9893_1155# VSS 6.69e-19
C258 a_9893_1293# VSS 6.32e-19
C259 nstack_lab7 VSS 0.119f
C260 a_15703_1340# VSS 0.293f
C261 x2.floating VSS 6.42f
C262 x3[1].floating VSS 10.9f
C263 x4[3].floating VSS 21.7f
C264 x7.floating VSS 5.93f
C265 code[0] VSS 0.761f
C266 code[1] VSS 0.911f
C267 code[2] VSS 1.61f
C268 x5[7].floating VSS 0.107p
C269 x6.floating VSS 0.414f
C270 a_15703_1681# VSS 0.32f
C271 Uc VSS 1.55f
C272 x6.SW VSS 0.299f
C273 x10.Y VSS 2.76f
C274 code_offset VSS 1.12f
C275 code[3] VSS 0.267f
C276 pstack_lab5 VSS 0.0143f
C277 pstack_lab4 VSS 0.0172f
C278 pstack_lab3 VSS 0.0815f
C279 pstack_lab2 VSS 0.0204f
C280 pstack_lab1 VSS 0.0953f
C281 IN VSS 1.44f
C282 VDD VSS 38.5f
C283 VDD.n0 VSS 0.024f
C284 VDD.t6 VSS 0.0579f
C285 VDD.n1 VSS 0.0207f
C286 VDD.n2 VSS 0.0142f
C287 VDD.n3 VSS 0.104f
C288 VDD.n4 VSS 0.0159f
C289 VDD.n5 VSS 0.00301f
C290 VDD.n6 VSS 0.00444f
C291 VDD.n7 VSS 0.0243f
C292 VDD.n8 VSS 0.00993f
C293 VDD.n9 VSS 0.00504f
C294 VDD.n10 VSS 0.00765f
C295 VDD.n11 VSS 0.00784f
C296 VDD.n12 VSS 0.0126f
C297 VDD.n13 VSS 0.00785f
C298 VDD.n14 VSS 9.27e-19
C299 VDD.n15 VSS 0.0212f
C300 VDD.n16 VSS 0.0194f
C301 VDD.n17 VSS 0.0264f
C302 VDD.n18 VSS 0.0466f
C303 VDD.n19 VSS 0.0225f
C304 VDD.n20 VSS 0.0181f
C305 VDD.n21 VSS 0.0141f
C306 VDD.n22 VSS 0.00341f
C307 VDD.n23 VSS 0.0689f
C308 VDD.n24 VSS 0.0141f
C309 VDD.n25 VSS 0.0312f
C310 VDD.n26 VSS 0.00463f
C311 VDD.n27 VSS 0.0209f
C312 VDD.t12 VSS 0.0579f
C313 VDD.n28 VSS 0.0677f
C314 VDD.t10 VSS 1.35f
C315 VDD.n29 VSS 0.0375f
C316 VDD.t16 VSS 0.487f
C317 VDD.t8 VSS 0.154f
C318 VDD.n30 VSS 0.464f
C319 VDD.n31 VSS 0.032f
C320 VDD.t2 VSS 2.48f
C321 VDD.t0 VSS 6.29f
C322 VDD.n32 VSS 5.3f
C323 VDD.n33 VSS 0.0348f
C324 VDD.n34 VSS 0.0348f
C325 VDD.n35 VSS 1.45f
C326 VDD.n36 VSS 0.00945f
C327 VDD.n37 VSS 0.0227f
C328 VDD.n38 VSS 0.0226f
C329 VDD.n39 VSS 0.0521f
C330 VDD.n40 VSS 0.0219f
C331 VDD.n41 VSS 0.0195f
C332 VDD.n42 VSS 0.00894f
C333 VDD.n43 VSS 0.0191f
C334 VDD.n44 VSS 0.00754f
C335 VDD.t9 VSS 0.00755f
C336 VDD.t15 VSS 0.00755f
C337 VDD.n45 VSS 0.0185f
C338 VDD.n46 VSS 0.0548f
C339 VDD.n47 VSS 0.00916f
C340 VDD.n48 VSS 0.0187f
C341 VDD.n49 VSS 0.114f
C342 VDD.n50 VSS 0.128f
C343 VDD.n51 VSS 0.0226f
C344 VDD.t1 VSS 0.0107f
C345 VDD.n52 VSS 0.155f
C346 VDD.n53 VSS 0.0228f
C347 VDD.n54 VSS 0.0123f
C348 VDD.n55 VSS 0.184f
C349 VDD.n56 VSS 0.184f
C350 VDD.n57 VSS 0.052f
C351 VDD.n58 VSS 0.0226f
C352 VDD.n59 VSS 0.00721f
C353 VDD.n60 VSS 0.00945f
C354 VDD.n61 VSS 0.0925f
C355 VDD.n62 VSS 0.0093f
C356 VDD.n63 VSS 0.0227f
C357 VDD.n64 VSS 0.052f
C358 VDD.n65 VSS 0.0226f
C359 VDD.n66 VSS 0.00721f
C360 VDD.n67 VSS 0.0227f
C361 VDD.n68 VSS 0.052f
C362 VDD.n69 VSS 0.0226f
C363 VDD.n70 VSS 0.00721f
C364 VDD.n71 VSS 0.0227f
C365 VDD.n72 VSS 0.052f
C366 VDD.n73 VSS 0.0226f
C367 VDD.n74 VSS 0.00721f
C368 VDD.n75 VSS 0.0227f
C369 VDD.n76 VSS 0.00637f
C370 VDD.n77 VSS 0.005f
C371 VDD.n78 VSS 0.00377f
C372 VDD.n79 VSS 5.39e-19
C373 VDD.n80 VSS 0.00305f
C374 VDD.n81 VSS 0.00305f
C375 VDD.n82 VSS 0.0146f
C376 VDD.n85 VSS 0.0118f
C377 VDD.n88 VSS 0.0266f
C378 VDD.n92 VSS 0.0118f
C379 VDD.n94 VSS 0.0118f
C380 VDD.n97 VSS 0.0266f
C381 VDD.n101 VSS 0.0118f
C382 VDD.n103 VSS 0.0118f
C383 VDD.n106 VSS 0.0266f
C384 VDD.n110 VSS 0.0118f
C385 VDD.n112 VSS 0.0118f
C386 VDD.n115 VSS 0.0266f
C387 VDD.n118 VSS 0.524f
C388 VDD.n119 VSS 0.023f
C389 VDD.n124 VSS 0.0266f
C390 VDD.n126 VSS 0.0118f
C391 VDD.n128 VSS 0.0118f
C392 VDD.n129 VSS 0.0197f
C393 VDD.n130 VSS 0.0197f
C394 VDD.n135 VSS 0.0266f
C395 VDD.n137 VSS 0.0118f
C396 VDD.n139 VSS 0.0118f
C397 VDD.n140 VSS 0.0197f
C398 VDD.n141 VSS 0.0197f
C399 VDD.n146 VSS 0.0266f
C400 VDD.n148 VSS 0.0118f
C401 VDD.n150 VSS 0.0118f
C402 VDD.n151 VSS 0.0197f
C403 VDD.n152 VSS 0.0197f
C404 VDD.n157 VSS 0.0266f
C405 VDD.n159 VSS 0.00315f
C406 VDD.n160 VSS 0.0146f
C407 VDD.n161 VSS 0.00305f
C408 VDD.n162 VSS 0.00305f
C409 VDD.n163 VSS 0.0104f
C410 VDD.n164 VSS 5.39e-19
C411 VDD.n165 VSS 0.00377f
C412 VDD.n166 VSS 0.00665f
C413 VDD.n167 VSS 0.00395f
C414 VDD.n168 VSS 5.39e-19
C415 VDD.n169 VSS 0.00537f
C416 VDD.n170 VSS 3.7e-19
C417 VDD.n171 VSS 0.0106f
C418 VDD.n172 VSS -0.0856f
C419 VDD.n173 VSS 0.0106f
C420 VDD.n174 VSS 0.00907f
C421 VDD.n175 VSS 0.00395f
C422 VDD.n176 VSS 0.00305f
C423 VDD.n177 VSS 0.00305f
C424 VDD.n178 VSS 0.00315f
C425 VDD.n179 VSS 0.00305f
C426 VDD.n180 VSS 0.0104f
C427 VDD.n181 VSS 0.00377f
C428 VDD.n182 VSS 0.005f
C429 VDD.n183 VSS -0.214f
C430 VDD.n184 VSS -0.106f
C431 VDD.n185 VSS 3.7e-19
C432 VDD.n186 VSS 0.00555f
C433 VDD.n187 VSS 0.00907f
C434 VDD.n188 VSS 0.00395f
C435 VDD.n189 VSS 0.0111f
C436 VDD.n190 VSS 0.0111f
C437 VDD.n191 VSS 0.00377f
C438 VDD.n192 VSS 0.00755f
C439 VDD.n193 VSS 0.00916f
C440 VDD.n194 VSS 0.00467f
C441 VDD.n195 VSS 0.00665f
C442 VDD.n196 VSS 0.00537f
C443 VDD.n197 VSS 0.00426f
C444 VDD.n198 VSS 0.0104f
C445 VDD.n199 VSS 0.00637f
C446 VDD.n200 VSS 0.00658f
C447 VDD.n201 VSS 3.7e-19
C448 VDD.n202 VSS 0.00555f
C449 VDD.n203 VSS 5.39e-19
C450 VDD.n204 VSS 0.00395f
C451 VDD.n205 VSS 3.59e-19
C452 VDD.n206 VSS 0.0118f
C453 VDD.n207 VSS 0.0146f
C454 VDD.n208 VSS 0.0111f
C455 VDD.n209 VSS 0.0111f
C456 VDD.n210 VSS 0.00377f
C457 VDD.n211 VSS 0.00755f
C458 VDD.n212 VSS 0.00916f
C459 VDD.n213 VSS 0.00377f
C460 VDD.n214 VSS 0.00467f
C461 VDD.n215 VSS 0.00665f
C462 VDD.n216 VSS -0.241f
C463 VDD.n217 VSS 0.00426f
C464 VDD.n218 VSS 0.0104f
C465 VDD.n219 VSS 0.00637f
C466 VDD.n220 VSS 0.00658f
C467 VDD.n221 VSS 3.7e-19
C468 VDD.n222 VSS 0.00555f
C469 VDD.n223 VSS 0.00907f
C470 VDD.n224 VSS 0.00426f
C471 VDD.n225 VSS 0.0104f
C472 VDD.n226 VSS 0.0104f
C473 VDD.n227 VSS 0.00555f
C474 VDD.n228 VSS 0.005f
C475 VDD.n229 VSS 0.00916f
C476 VDD.n230 VSS 0.00377f
C477 VDD.n231 VSS 0.00755f
C478 VDD.n232 VSS 5.39e-19
C479 VDD.n233 VSS 0.00305f
C480 VDD.n234 VSS 0.0111f
C481 VDD.n235 VSS 0.0111f
C482 VDD.n236 VSS 0.00315f
C483 VDD.n237 VSS 0.00305f
C484 VDD.n238 VSS 3.59e-19
C485 VDD.n239 VSS 0.00305f
C486 VDD.n240 VSS 0.00395f
C487 VDD.n241 VSS 0.00305f
C488 VDD.n242 VSS 0.00377f
C489 VDD.n243 VSS 0.0111f
C490 VDD.n244 VSS 0.0146f
C491 VDD.n245 VSS 0.0111f
C492 VDD.n246 VSS 0.00305f
C493 VDD.n247 VSS 0.0111f
C494 VDD.n248 VSS 0.0104f
C495 VDD.n249 VSS 0.00395f
C496 VDD.n250 VSS 0.00467f
C497 VDD.n251 VSS 0.00426f
C498 VDD.n252 VSS 3.7e-19
C499 VDD.n253 VSS 0.00637f
C500 VDD.n254 VSS 0.00658f
C501 VDD.n255 VSS 3.7e-19
C502 VDD.n256 VSS 0.00555f
C503 VDD.n257 VSS 0.00907f
C504 VDD.n258 VSS 0.0106f
C505 VDD.n259 VSS 0.0104f
C506 VDD.n260 VSS 0.00637f
C507 VDD.n261 VSS 0.00395f
C508 VDD.n262 VSS 0.00555f
C509 VDD.n263 VSS 0.00305f
C510 VDD.n264 VSS 0.0146f
C511 VDD.n265 VSS 0.00315f
C512 VDD.n266 VSS 0.00305f
C513 VDD.n267 VSS 0.0334f
C514 VDD.n268 VSS 0.0296f
C515 VDD.n269 VSS 5.39e-19
C516 VDD.n270 VSS 0.00377f
C517 VDD.n271 VSS 0.00395f
C518 VDD.n272 VSS 0.00305f
C519 VDD.n273 VSS 0.00755f
C520 VDD.n274 VSS 0.00395f
C521 VDD.n275 VSS 0.00916f
C522 VDD.n276 VSS 0.00377f
C523 VDD.n277 VSS 0.00889f
C524 VDD.n278 VSS 0.005f
C525 VDD.n279 VSS 0.00658f
C526 VDD.n280 VSS 0.00537f
C527 VDD.n281 VSS 0.00658f
C528 VDD.n282 VSS 0.0376f
C529 VDD.n283 VSS 0.0326f
C530 VDD.n284 VSS 0.0324f
C531 VDD.n285 VSS 0.0374f
C532 VDD.n286 VSS 0.00637f
C533 VDD.n287 VSS 3.7e-19
C534 VDD.n288 VSS -0.0856f
C535 VDD.n289 VSS 0.00377f
C536 VDD.n290 VSS 0.0104f
C537 VDD.n291 VSS 0.00467f
C538 VDD.n292 VSS 0.00665f
C539 VDD.n293 VSS -0.24f
C540 VDD.n294 VSS 0.00444f
C541 VDD.n295 VSS 0.0106f
C542 VDD.n296 VSS 0.0104f
C543 VDD.n297 VSS -0.222f
C544 VDD.n298 VSS 0.00555f
C545 VDD.n299 VSS 3.7e-19
C546 VDD.n300 VSS 0.00395f
C547 VDD.n301 VSS 0.00377f
C548 VDD.n302 VSS 0.00305f
C549 VDD.n303 VSS 0.0104f
C550 VDD.n304 VSS 0.00305f
C551 VDD.n305 VSS 0.00305f
C552 VDD.n306 VSS 0.00755f
C553 VDD.n307 VSS 0.00395f
C554 VDD.n308 VSS 0.00916f
C555 VDD.n309 VSS 0.00377f
C556 VDD.n310 VSS 0.00889f
C557 VDD.n311 VSS -0.0856f
C558 VDD.n312 VSS -0.0981f
C559 VDD.n313 VSS 0.00658f
C560 VDD.n314 VSS 0.005f
C561 VDD.n315 VSS 0.00467f
C562 VDD.n316 VSS 0.00665f
C563 VDD.n317 VSS 0.00555f
C564 VDD.n318 VSS 0.00444f
C565 VDD.n319 VSS 0.0106f
C566 VDD.n320 VSS 0.0104f
C567 VDD.n321 VSS 0.0104f
C568 VDD.n322 VSS -0.24f
C569 VDD.n323 VSS 3.7e-19
C570 VDD.n324 VSS 0.00395f
C571 VDD.n325 VSS 0.00377f
C572 VDD.n326 VSS 0.00305f
C573 VDD.n327 VSS 0.0104f
C574 VDD.n328 VSS 0.00305f
C575 VDD.n329 VSS 0.00305f
C576 VDD.n330 VSS 0.00755f
C577 VDD.n331 VSS 0.00395f
C578 VDD.n332 VSS 0.00916f
C579 VDD.n333 VSS 0.00377f
C580 VDD.n334 VSS 0.00889f
C581 VDD.n335 VSS 0.005f
C582 VDD.n336 VSS 0.00637f
C583 VDD.n337 VSS 0.00658f
C584 VDD.n338 VSS 0.005f
C585 VDD.n339 VSS 0.00467f
C586 VDD.n340 VSS 0.00665f
C587 VDD.n341 VSS 0.00555f
C588 VDD.n342 VSS 0.00444f
C589 VDD.n343 VSS 0.0106f
C590 VDD.n344 VSS -0.222f
C591 VDD.n345 VSS 0.00555f
C592 VDD.n346 VSS 0.00537f
C593 VDD.n347 VSS -0.106f
C594 VDD.n348 VSS 3.7e-19
C595 VDD.n349 VSS 0.00467f
C596 VDD.n350 VSS 0.00395f
C597 VDD.n351 VSS 0.00555f
C598 VDD.n352 VSS 0.0286f
C599 VDD.n353 VSS 0.0286f
C600 VDD.n354 VSS 0.00467f
C601 VDD.n355 VSS 0.0336f
C602 VDD.n356 VSS 0.0336f
C603 VDD.n357 VSS 0.00305f
C604 VDD.n358 VSS 3.59e-19
C605 VDD.n359 VSS 0.0118f
C606 VDD.n360 VSS 0.00315f
C607 VDD.n361 VSS 0.00305f
C608 VDD.n362 VSS 0.0355f
C609 VDD.n363 VSS 0.0355f
C610 VDD.n364 VSS 0.00315f
C611 VDD.n365 VSS 0.00305f
C612 VDD.n366 VSS 0.0146f
C613 VDD.n367 VSS 0.0111f
C614 VDD.n368 VSS 0.0104f
C615 VDD.n369 VSS 0.00467f
C616 VDD.n370 VSS 0.00426f
C617 VDD.n371 VSS 3.7e-19
C618 VDD.n372 VSS 0.00907f
C619 VDD.n373 VSS -0.214f
C620 VDD.n374 VSS 0.0104f
C621 VDD.n375 VSS 0.00637f
C622 VDD.n376 VSS 0.00395f
C623 VDD.n377 VSS 0.00555f
C624 VDD.n378 VSS 0.00305f
C625 VDD.n379 VSS 0.00315f
C626 VDD.n380 VSS 0.00305f
C627 VDD.n381 VSS 0.0146f
C628 VDD.n382 VSS 0.0111f
C629 VDD.n383 VSS 0.0104f
C630 VDD.n384 VSS 0.00467f
C631 VDD.n385 VSS 0.00426f
C632 VDD.n386 VSS 3.7e-19
C633 VDD.n387 VSS 0.00658f
C634 VDD.n388 VSS 0.00907f
C635 VDD.n389 VSS 0.0106f
C636 VDD.n390 VSS 0.0104f
C637 VDD.n391 VSS 0.00637f
C638 VDD.n392 VSS 0.00395f
C639 VDD.n393 VSS 0.00555f
C640 VDD.n394 VSS 0.00305f
C641 VDD.n395 VSS 0.00315f
C642 VDD.n396 VSS 0.00305f
C643 VDD.n397 VSS 0.0146f
C644 VDD.n398 VSS 0.0111f
C645 VDD.n399 VSS 0.0104f
C646 VDD.n400 VSS 0.00467f
C647 VDD.n401 VSS 0.00426f
C648 VDD.n402 VSS 3.7e-19
C649 VDD.n403 VSS 0.00658f
C650 VDD.n404 VSS 0.00907f
C651 VDD.n405 VSS 0.0106f
C652 VDD.n406 VSS 0.0104f
C653 VDD.n407 VSS 0.00637f
C654 VDD.n408 VSS 0.00395f
C655 VDD.n409 VSS 0.00555f
C656 VDD.n410 VSS 0.00305f
C657 VDD.n411 VSS 0.00315f
C658 VDD.n412 VSS 0.00305f
C659 VDD.n413 VSS 0.0146f
C660 VDD.n414 VSS 0.0111f
C661 VDD.n415 VSS 0.0104f
C662 VDD.n416 VSS 0.00467f
C663 VDD.n417 VSS 0.00426f
C664 VDD.n418 VSS 3.7e-19
C665 VDD.n419 VSS -0.106f
C666 VDD.n420 VSS 0.00907f
C667 VDD.n421 VSS -0.214f
C668 VDD.n422 VSS 0.0104f
C669 VDD.n423 VSS 0.00637f
C670 VDD.n424 VSS 0.00395f
C671 VDD.n425 VSS 0.00555f
C672 VDD.n426 VSS 0.00305f
C673 VDD.n427 VSS 0.00305f
C674 VDD.n428 VSS 0.0111f
C675 VDD.n429 VSS 0.0104f
C676 VDD.n430 VSS 0.00467f
C677 VDD.n431 VSS 0.00426f
C678 VDD.n432 VSS 3.7e-19
C679 VDD.n433 VSS 0.00658f
C680 VDD.n434 VSS 0.00907f
C681 VDD.n435 VSS 0.0106f
C682 VDD.n436 VSS 0.0104f
C683 VDD.n437 VSS 0.00637f
C684 VDD.n438 VSS 0.00395f
C685 VDD.n439 VSS 0.00555f
C686 VDD.n440 VSS 0.00305f
C687 VDD.n441 VSS 0.0146f
C688 VDD.n442 VSS 0.00315f
C689 VDD.n443 VSS 0.00305f
C690 VDD.n444 VSS 0.0334f
C691 VDD.n445 VSS 0.0296f
C692 VDD.n446 VSS 5.39e-19
C693 VDD.n447 VSS 0.00377f
C694 VDD.n448 VSS 0.00395f
C695 VDD.n449 VSS 0.00305f
C696 VDD.n450 VSS 0.00755f
C697 VDD.n451 VSS 0.00395f
C698 VDD.n452 VSS 0.00916f
C699 VDD.n453 VSS 0.00377f
C700 VDD.n454 VSS 0.00889f
C701 VDD.n455 VSS 0.005f
C702 VDD.n456 VSS 0.00658f
C703 VDD.n457 VSS 0.00537f
C704 VDD.n458 VSS 0.00658f
C705 VDD.n459 VSS 0.0376f
C706 VDD.n460 VSS 0.0326f
C707 VDD.n461 VSS 0.0324f
C708 VDD.n462 VSS 0.0374f
C709 VDD.n463 VSS 0.00637f
C710 VDD.n464 VSS 3.7e-19
C711 VDD.n465 VSS -0.0856f
C712 VDD.n466 VSS 0.00377f
C713 VDD.n467 VSS 0.0104f
C714 VDD.n468 VSS 0.00467f
C715 VDD.n469 VSS 0.00665f
C716 VDD.n470 VSS -0.24f
C717 VDD.n471 VSS 0.00444f
C718 VDD.n472 VSS 0.0106f
C719 VDD.n473 VSS 0.0104f
C720 VDD.n474 VSS -0.222f
C721 VDD.n475 VSS 0.00555f
C722 VDD.n476 VSS 3.7e-19
C723 VDD.n477 VSS 0.00395f
C724 VDD.n478 VSS 0.00377f
C725 VDD.n479 VSS 0.00305f
C726 VDD.n480 VSS 0.0104f
C727 VDD.n481 VSS 0.00305f
C728 VDD.n482 VSS 0.00305f
C729 VDD.n483 VSS 0.00755f
C730 VDD.n484 VSS 0.00395f
C731 VDD.n485 VSS 0.00916f
C732 VDD.n486 VSS 0.00377f
C733 VDD.n487 VSS 0.00889f
C734 VDD.n488 VSS -0.0856f
C735 VDD.n489 VSS -0.0981f
C736 VDD.n490 VSS 0.00658f
C737 VDD.n491 VSS 0.005f
C738 VDD.n492 VSS 0.00467f
C739 VDD.n493 VSS 0.00665f
C740 VDD.n494 VSS 0.00555f
C741 VDD.n495 VSS 0.00444f
C742 VDD.n496 VSS 0.0106f
C743 VDD.n497 VSS 0.0104f
C744 VDD.n498 VSS 0.0104f
C745 VDD.n499 VSS -0.24f
C746 VDD.n500 VSS 3.7e-19
C747 VDD.n501 VSS 0.00395f
C748 VDD.n502 VSS 0.00377f
C749 VDD.n503 VSS 0.00305f
C750 VDD.n504 VSS 0.0104f
C751 VDD.n505 VSS 0.00305f
C752 VDD.n506 VSS 0.00305f
C753 VDD.n507 VSS 0.00755f
C754 VDD.n508 VSS 0.00395f
C755 VDD.n509 VSS 0.00916f
C756 VDD.n510 VSS 0.00377f
C757 VDD.n511 VSS 0.00889f
C758 VDD.n512 VSS 0.005f
C759 VDD.n513 VSS 0.00637f
C760 VDD.n514 VSS 0.00658f
C761 VDD.n515 VSS 0.005f
C762 VDD.n516 VSS 0.00467f
C763 VDD.n517 VSS 0.00665f
C764 VDD.n518 VSS 0.00555f
C765 VDD.n519 VSS 0.00444f
C766 VDD.n520 VSS 0.0106f
C767 VDD.n521 VSS -0.222f
C768 VDD.n522 VSS 0.00555f
C769 VDD.n523 VSS 0.00537f
C770 VDD.n524 VSS -0.106f
C771 VDD.n525 VSS 3.7e-19
C772 VDD.n526 VSS 0.00467f
C773 VDD.n527 VSS 0.00395f
C774 VDD.n528 VSS 0.00555f
C775 VDD.n529 VSS 0.0286f
C776 VDD.n530 VSS 0.0286f
C777 VDD.n531 VSS 0.00467f
C778 VDD.n532 VSS 0.0336f
C779 VDD.n533 VSS 0.0336f
C780 VDD.n534 VSS 0.00305f
C781 VDD.n535 VSS 3.59e-19
C782 VDD.n536 VSS 0.0118f
C783 VDD.n537 VSS 0.00315f
C784 VDD.n538 VSS 0.00305f
C785 VDD.n539 VSS 0.0355f
C786 VDD.n540 VSS 0.0355f
C787 VDD.n541 VSS 0.00315f
C788 VDD.n542 VSS 0.00305f
C789 VDD.n543 VSS 0.0146f
C790 VDD.n544 VSS 0.0111f
C791 VDD.n545 VSS 0.0104f
C792 VDD.n546 VSS 0.00467f
C793 VDD.n547 VSS 0.00426f
C794 VDD.n548 VSS 3.7e-19
C795 VDD.n549 VSS 0.00907f
C796 VDD.n550 VSS -0.214f
C797 VDD.n551 VSS 0.0104f
C798 VDD.n552 VSS 0.00637f
C799 VDD.n553 VSS 0.00395f
C800 VDD.n554 VSS 0.00555f
C801 VDD.n555 VSS 0.00305f
C802 VDD.n556 VSS 0.00315f
C803 VDD.n557 VSS 0.00305f
C804 VDD.n558 VSS 0.0146f
C805 VDD.n559 VSS 0.0111f
C806 VDD.n560 VSS 0.0104f
C807 VDD.n561 VSS 0.00467f
C808 VDD.n562 VSS 0.00426f
C809 VDD.n563 VSS 3.7e-19
C810 VDD.n564 VSS 0.00658f
C811 VDD.n565 VSS 0.00907f
C812 VDD.n566 VSS 0.0106f
C813 VDD.n567 VSS 0.0104f
C814 VDD.n568 VSS 0.00637f
C815 VDD.n569 VSS 0.00395f
C816 VDD.n570 VSS 0.00555f
C817 VDD.n571 VSS 0.00305f
C818 VDD.n572 VSS 0.00315f
C819 VDD.n573 VSS 0.00305f
C820 VDD.n574 VSS 0.0146f
C821 VDD.n575 VSS 0.0111f
C822 VDD.n576 VSS 0.0104f
C823 VDD.n577 VSS 0.00467f
C824 VDD.n578 VSS 0.00426f
C825 VDD.n579 VSS 3.7e-19
C826 VDD.n580 VSS 0.00658f
C827 VDD.n581 VSS 0.00907f
C828 VDD.n582 VSS 0.0106f
C829 VDD.n583 VSS 0.0104f
C830 VDD.n584 VSS 0.00637f
C831 VDD.n585 VSS 0.00395f
C832 VDD.n586 VSS 0.00555f
C833 VDD.n587 VSS 0.00305f
C834 VDD.n588 VSS 0.00315f
C835 VDD.n589 VSS 0.00305f
C836 VDD.n590 VSS 0.0146f
C837 VDD.n591 VSS 0.0111f
C838 VDD.n592 VSS 0.0104f
C839 VDD.n593 VSS 0.00467f
C840 VDD.n594 VSS 0.00426f
C841 VDD.n595 VSS 3.7e-19
C842 VDD.n596 VSS -0.106f
C843 VDD.n597 VSS 0.00907f
C844 VDD.n598 VSS -0.214f
C845 VDD.n599 VSS 0.0104f
C846 VDD.n600 VSS 0.00637f
C847 VDD.n601 VSS 0.00395f
C848 VDD.n602 VSS 0.00555f
C849 VDD.n603 VSS 0.00305f
C850 VDD.n604 VSS 0.00305f
C851 VDD.n605 VSS 0.0111f
C852 VDD.n606 VSS 0.0104f
C853 VDD.n607 VSS 0.00467f
C854 VDD.n608 VSS 0.00426f
C855 VDD.n609 VSS 3.7e-19
C856 VDD.n610 VSS 0.00658f
C857 VDD.n611 VSS 0.00907f
C858 VDD.n612 VSS 0.0106f
C859 VDD.n613 VSS 0.0104f
C860 VDD.n614 VSS 0.00637f
C861 VDD.n615 VSS 0.00395f
C862 VDD.n616 VSS 0.00555f
C863 VDD.n617 VSS 0.00305f
C864 VDD.n618 VSS 0.0146f
C865 VDD.n619 VSS 0.00315f
C866 VDD.n620 VSS 0.00305f
C867 VDD.n621 VSS 0.0334f
C868 VDD.n622 VSS 0.0296f
C869 VDD.n623 VSS 5.39e-19
C870 VDD.n624 VSS 0.00377f
C871 VDD.n625 VSS 0.00395f
C872 VDD.n626 VSS 0.00305f
C873 VDD.n627 VSS 0.00755f
C874 VDD.n628 VSS 0.00395f
C875 VDD.n629 VSS 0.00916f
C876 VDD.n630 VSS 0.00377f
C877 VDD.n631 VSS 0.00889f
C878 VDD.n632 VSS 0.005f
C879 VDD.n633 VSS 0.00658f
C880 VDD.n634 VSS 0.00537f
C881 VDD.n635 VSS 0.00658f
C882 VDD.n636 VSS 0.0376f
C883 VDD.n637 VSS 0.0326f
C884 VDD.n638 VSS 0.0324f
C885 VDD.n639 VSS 0.0374f
C886 VDD.n640 VSS 0.00637f
C887 VDD.n641 VSS 3.7e-19
C888 VDD.n642 VSS -0.0856f
C889 VDD.n643 VSS 0.00377f
C890 VDD.n644 VSS 0.0104f
C891 VDD.n645 VSS 0.00467f
C892 VDD.n646 VSS 0.00665f
C893 VDD.n647 VSS -0.24f
C894 VDD.n648 VSS 0.00444f
C895 VDD.n649 VSS 0.0106f
C896 VDD.n650 VSS 0.0104f
C897 VDD.n651 VSS -0.222f
C898 VDD.n652 VSS 0.00555f
C899 VDD.n653 VSS 3.7e-19
C900 VDD.n654 VSS 0.00395f
C901 VDD.n655 VSS 0.00377f
C902 VDD.n656 VSS 0.00305f
C903 VDD.n657 VSS 0.0104f
C904 VDD.n658 VSS 0.00305f
C905 VDD.n659 VSS 0.00305f
C906 VDD.n660 VSS 0.00755f
C907 VDD.n661 VSS 0.00395f
C908 VDD.n662 VSS 0.00916f
C909 VDD.n663 VSS 0.00377f
C910 VDD.n664 VSS 0.00889f
C911 VDD.n665 VSS -0.0856f
C912 VDD.n666 VSS -0.0981f
C913 VDD.n667 VSS 0.00658f
C914 VDD.n668 VSS 0.005f
C915 VDD.n669 VSS 0.00467f
C916 VDD.n670 VSS 0.00665f
C917 VDD.n671 VSS 0.00555f
C918 VDD.n672 VSS 0.00444f
C919 VDD.n673 VSS 0.0106f
C920 VDD.n674 VSS 0.0104f
C921 VDD.n675 VSS 0.0104f
C922 VDD.n676 VSS -0.24f
C923 VDD.n677 VSS 3.7e-19
C924 VDD.n678 VSS 0.00395f
C925 VDD.n679 VSS 0.00377f
C926 VDD.n680 VSS 0.00305f
C927 VDD.n681 VSS 0.0104f
C928 VDD.n682 VSS 0.00305f
C929 VDD.n683 VSS 0.00305f
C930 VDD.n684 VSS 0.00755f
C931 VDD.n685 VSS 0.00395f
C932 VDD.n686 VSS 0.00916f
C933 VDD.n687 VSS 0.00377f
C934 VDD.n688 VSS 0.00889f
C935 VDD.n689 VSS 0.005f
C936 VDD.n690 VSS 0.00637f
C937 VDD.n691 VSS 0.00658f
C938 VDD.n692 VSS 0.005f
C939 VDD.n693 VSS 0.00467f
C940 VDD.n694 VSS 0.00665f
C941 VDD.n695 VSS 0.00555f
C942 VDD.n696 VSS 0.00444f
C943 VDD.n697 VSS 0.0106f
C944 VDD.n698 VSS -0.222f
C945 VDD.n699 VSS 0.00555f
C946 VDD.n700 VSS 0.00537f
C947 VDD.n701 VSS -0.106f
C948 VDD.n702 VSS 3.7e-19
C949 VDD.n703 VSS 0.00467f
C950 VDD.n704 VSS 0.00395f
C951 VDD.n705 VSS 0.00555f
C952 VDD.n706 VSS 0.0286f
C953 VDD.n707 VSS 0.0286f
C954 VDD.n708 VSS 0.00467f
C955 VDD.n709 VSS 0.0336f
C956 VDD.n710 VSS 0.0336f
C957 VDD.n711 VSS 0.00305f
C958 VDD.n712 VSS 3.59e-19
C959 VDD.n713 VSS 0.0118f
C960 VDD.n714 VSS 0.00315f
C961 VDD.n715 VSS 0.00305f
C962 VDD.n716 VSS 0.0355f
C963 VDD.n717 VSS 0.0355f
C964 VDD.n718 VSS 0.00315f
C965 VDD.n719 VSS 0.00305f
C966 VDD.n720 VSS 0.0146f
C967 VDD.n721 VSS 0.0111f
C968 VDD.n722 VSS 0.0104f
C969 VDD.n723 VSS 0.00467f
C970 VDD.n724 VSS 0.00426f
C971 VDD.n725 VSS 3.7e-19
C972 VDD.n726 VSS 0.00907f
C973 VDD.n727 VSS -0.214f
C974 VDD.n728 VSS 0.0104f
C975 VDD.n729 VSS 0.00637f
C976 VDD.n730 VSS 0.00395f
C977 VDD.n731 VSS 0.00555f
C978 VDD.n732 VSS 0.00305f
C979 VDD.n733 VSS 0.00315f
C980 VDD.n734 VSS 0.00305f
C981 VDD.n735 VSS 0.0146f
C982 VDD.n736 VSS 0.0111f
C983 VDD.n737 VSS 0.0104f
C984 VDD.n738 VSS 0.00467f
C985 VDD.n739 VSS 0.00426f
C986 VDD.n740 VSS 3.7e-19
C987 VDD.n741 VSS 0.00658f
C988 VDD.n742 VSS 0.00907f
C989 VDD.n743 VSS 0.0106f
C990 VDD.n744 VSS 0.0104f
C991 VDD.n745 VSS 0.00637f
C992 VDD.n746 VSS 0.00395f
C993 VDD.n747 VSS 0.00555f
C994 VDD.n748 VSS 0.00305f
C995 VDD.n749 VSS 0.00315f
C996 VDD.n750 VSS 0.00305f
C997 VDD.n751 VSS 0.0146f
C998 VDD.n752 VSS 0.0111f
C999 VDD.n753 VSS 0.0104f
C1000 VDD.n754 VSS 0.00467f
C1001 VDD.n755 VSS 0.00426f
C1002 VDD.n756 VSS 3.7e-19
C1003 VDD.n757 VSS 0.00658f
C1004 VDD.n758 VSS 0.00907f
C1005 VDD.n759 VSS 0.0106f
C1006 VDD.n760 VSS 0.0104f
C1007 VDD.n761 VSS 0.00637f
C1008 VDD.n762 VSS 0.00395f
C1009 VDD.n763 VSS 0.00555f
C1010 VDD.n764 VSS 0.00305f
C1011 VDD.n765 VSS 0.00315f
C1012 VDD.n766 VSS 0.00305f
C1013 VDD.n767 VSS 0.0146f
C1014 VDD.n768 VSS 0.0111f
C1015 VDD.n769 VSS 0.0104f
C1016 VDD.n770 VSS 0.00467f
C1017 VDD.n771 VSS 0.00426f
C1018 VDD.n772 VSS 3.7e-19
C1019 VDD.n773 VSS -0.106f
C1020 VDD.n774 VSS 0.00907f
C1021 VDD.n775 VSS -0.214f
C1022 VDD.n776 VSS 0.0104f
C1023 VDD.n777 VSS 0.00637f
C1024 VDD.n778 VSS 0.00395f
C1025 VDD.n779 VSS 0.00555f
C1026 VDD.n780 VSS 0.00305f
C1027 VDD.n781 VSS 0.00305f
C1028 VDD.n782 VSS 0.0111f
C1029 VDD.n783 VSS 0.0104f
C1030 VDD.n784 VSS 0.00467f
C1031 VDD.n785 VSS 0.00426f
C1032 VDD.n786 VSS 3.7e-19
C1033 VDD.n787 VSS 0.00658f
C1034 VDD.n788 VSS 0.00907f
C1035 VDD.n789 VSS 0.0106f
C1036 VDD.n790 VSS 0.0104f
C1037 VDD.n791 VSS 0.00637f
C1038 VDD.n792 VSS 0.00395f
C1039 VDD.n793 VSS 0.00555f
C1040 VDD.n794 VSS 0.00305f
C1041 VDD.n795 VSS 0.0146f
C1042 VDD.n796 VSS 0.00315f
C1043 VDD.n797 VSS 0.00305f
C1044 VDD.n798 VSS 0.0334f
C1045 VDD.n799 VSS 0.0296f
C1046 VDD.n800 VSS 5.39e-19
C1047 VDD.n801 VSS 0.00377f
C1048 VDD.n802 VSS 0.00395f
C1049 VDD.n803 VSS 0.00305f
C1050 VDD.n804 VSS 0.00755f
C1051 VDD.n805 VSS 0.00395f
C1052 VDD.n806 VSS 0.00916f
C1053 VDD.n807 VSS 0.00377f
C1054 VDD.n808 VSS 0.00889f
C1055 VDD.n809 VSS 0.005f
C1056 VDD.n810 VSS 0.00658f
C1057 VDD.n811 VSS 0.00537f
C1058 VDD.n812 VSS 0.00658f
C1059 VDD.n813 VSS 0.0376f
C1060 VDD.n814 VSS 0.0326f
C1061 VDD.n815 VSS 0.0324f
C1062 VDD.n816 VSS 0.0374f
C1063 VDD.n817 VSS 0.00637f
C1064 VDD.n818 VSS 3.7e-19
C1065 VDD.n819 VSS -0.0856f
C1066 VDD.n820 VSS 0.00377f
C1067 VDD.n821 VSS 0.0104f
C1068 VDD.n822 VSS 0.00467f
C1069 VDD.n823 VSS 0.00665f
C1070 VDD.n824 VSS -0.24f
C1071 VDD.n825 VSS 0.00444f
C1072 VDD.n826 VSS 0.0106f
C1073 VDD.n827 VSS 0.0104f
C1074 VDD.n828 VSS -0.222f
C1075 VDD.n829 VSS 0.00555f
C1076 VDD.n830 VSS 3.7e-19
C1077 VDD.n831 VSS 0.00395f
C1078 VDD.n832 VSS 0.00377f
C1079 VDD.n833 VSS 0.00305f
C1080 VDD.n834 VSS 0.0104f
C1081 VDD.n835 VSS 0.00305f
C1082 VDD.n836 VSS 0.00305f
C1083 VDD.n837 VSS 0.00755f
C1084 VDD.n838 VSS 0.00395f
C1085 VDD.n839 VSS 0.00916f
C1086 VDD.n840 VSS 0.00377f
C1087 VDD.n841 VSS 0.00889f
C1088 VDD.n842 VSS -0.0856f
C1089 VDD.n843 VSS -0.0981f
C1090 VDD.n844 VSS 0.00658f
C1091 VDD.n845 VSS 0.005f
C1092 VDD.n846 VSS 0.00467f
C1093 VDD.n847 VSS 0.00665f
C1094 VDD.n848 VSS 0.00555f
C1095 VDD.n849 VSS 0.00444f
C1096 VDD.n850 VSS 0.0106f
C1097 VDD.n851 VSS 0.0104f
C1098 VDD.n852 VSS 0.0104f
C1099 VDD.n853 VSS -0.24f
C1100 VDD.n854 VSS 3.7e-19
C1101 VDD.n855 VSS 0.00395f
C1102 VDD.n856 VSS 0.00377f
C1103 VDD.n857 VSS 0.00305f
C1104 VDD.n858 VSS 0.0104f
C1105 VDD.n859 VSS 0.00305f
C1106 VDD.n860 VSS 0.00305f
C1107 VDD.n861 VSS 0.00755f
C1108 VDD.n862 VSS 0.0586f
C1109 VDD.n863 VSS 0.0479f
C1110 VDD.n864 VSS 0.00916f
C1111 VDD.n865 VSS 0.00377f
C1112 VDD.n866 VSS 0.00889f
C1113 VDD.n867 VSS 0.005f
C1114 VDD.n868 VSS 0.00637f
C1115 VDD.n869 VSS 0.00658f
C1116 VDD.n870 VSS 0.005f
C1117 VDD.n871 VSS 0.00467f
C1118 VDD.n872 VSS 0.00665f
C1119 VDD.n873 VSS 0.00555f
C1120 VDD.n874 VSS 0.00444f
C1121 VDD.n875 VSS 0.0106f
C1122 VDD.n876 VSS -0.222f
C1123 VDD.n877 VSS 0.00661f
C1124 VDD.n878 VSS 3.7e-19
C1125 VDD.n879 VSS 0.0656f
C1126 VDD.n880 VSS 0.00467f
C1127 VDD.n881 VSS -0.24f
C1128 VDD.n882 VSS 0.0108f
C1129 VDD.n883 VSS 3.7e-19
C1130 VDD.n884 VSS 0.00395f
C1131 VDD.n885 VSS 0.00377f
C1132 VDD.n886 VSS 0.00305f
C1133 VDD.n887 VSS 0.0104f
C1134 VDD.n888 VSS 0.00305f
C1135 VDD.n889 VSS 0.00305f
C1136 VDD.n891 VSS 0.0357f
C1137 VDD.n892 VSS 0.0268f
C1138 VDD.n893 VSS 0.00315f
C1139 VDD.n894 VSS 0.00305f
C1140 VDD.n895 VSS 0.0108f
C1141 VDD.n896 VSS 0.00665f
C1142 VDD.n897 VSS 0.00916f
C1143 VDD.n898 VSS 0.00755f
C1144 VDD.n899 VSS 0.00377f
C1145 VDD.n900 VSS 0.0111f
C1146 VDD.n901 VSS 0.0111f
C1147 VDD.n902 VSS 0.0146f
C1148 VDD.n903 VSS 0.0118f
C1149 VDD.n904 VSS 0.00305f
C1150 VDD.n905 VSS 0.00755f
C1151 VDD.n906 VSS 0.00395f
C1152 VDD.n907 VSS 0.00916f
C1153 VDD.n908 VSS 0.00377f
C1154 VDD.n909 VSS 0.00889f
C1155 VDD.n910 VSS 0.005f
C1156 VDD.n911 VSS 0.00661f
C1157 VDD.n912 VSS 0.00683f
C1158 VDD.n913 VSS 0.005f
C1159 VDD.n914 VSS 0.00467f
C1160 VDD.n915 VSS 0.00665f
C1161 VDD.n916 VSS 0.00555f
C1162 VDD.n917 VSS 0.00444f
C1163 VDD.n918 VSS 0.011f
C1164 VDD.n919 VSS -0.221f
C1165 VDD.n920 VSS 0.0108f
C1166 VDD.n921 VSS 0.00555f
C1167 VDD.n922 VSS 3.7e-19
C1168 VDD.n923 VSS 0.00395f
C1169 VDD.n924 VSS 0.00377f
C1170 VDD.n925 VSS 0.00305f
C1171 VDD.n926 VSS 0.0104f
C1172 VDD.n927 VSS 0.00305f
C1173 VDD.n928 VSS 0.00305f
C1174 VDD.n930 VSS 0.00315f
C1175 VDD.n931 VSS 3.59e-19
C1176 VDD.n932 VSS 0.00305f
C1177 VDD.n933 VSS 0.0104f
C1178 VDD.n934 VSS 0.00467f
C1179 VDD.n935 VSS 0.00665f
C1180 VDD.n936 VSS 0.00916f
C1181 VDD.n937 VSS 0.00755f
C1182 VDD.n938 VSS 0.00377f
C1183 VDD.n939 VSS 0.0111f
C1184 VDD.n940 VSS 0.0111f
C1185 VDD.n941 VSS 0.0146f
C1186 VDD.n942 VSS 0.0118f
C1187 VDD.n943 VSS 0.00305f
C1188 VDD.n944 VSS 0.00755f
C1189 VDD.n945 VSS 0.00395f
C1190 VDD.n946 VSS 0.00916f
C1191 VDD.n947 VSS 0.00377f
C1192 VDD.n948 VSS 0.00889f
C1193 VDD.n949 VSS 0.005f
C1194 VDD.n950 VSS 0.00661f
C1195 VDD.n951 VSS 0.00683f
C1196 VDD.n952 VSS -0.0856f
C1197 VDD.n953 VSS 0.00467f
C1198 VDD.n954 VSS 0.00665f
C1199 VDD.n955 VSS -0.24f
C1200 VDD.n956 VSS 0.00444f
C1201 VDD.n957 VSS 0.011f
C1202 VDD.n958 VSS 0.0108f
C1203 VDD.n959 VSS -0.221f
C1204 VDD.n960 VSS 0.00555f
C1205 VDD.n961 VSS 3.7e-19
C1206 VDD.n962 VSS 0.00395f
C1207 VDD.n963 VSS 0.00377f
C1208 VDD.n964 VSS 0.00305f
C1209 VDD.n965 VSS 0.018f
C1210 VDD.n966 VSS 0.00305f
C1211 VDD.n967 VSS 0.00344f
C1212 VDD.t4 VSS 0.00664f
C1213 VDD.n968 VSS 0.0138f
C1214 VDD.n969 VSS 0.00843f
C1215 VDD.n970 VSS 0.00702f
C1216 VDD.n971 VSS 0.0302f
C1217 VDD.n972 VSS 0.00467f
C1218 VDD.n973 VSS 0.00887f
C1219 VDD.n974 VSS 0.00555f
C1220 VDD.n975 VSS -0.0978f
C1221 VDD.n976 VSS 0.005f
C1222 VDD.n977 VSS 0.00683f
C1223 VDD.n978 VSS 0.00727f
C1224 VDD.n979 VSS 0.00872f
C1225 VDD.n980 VSS 0.00928f
C1226 VDD.n981 VSS 0.0148f
C1227 VDD.n982 VSS 0.014f
C1228 VDD.n983 VSS 0.0126f
C1229 VDD.n984 VSS 0.00121f
C1230 VDD.n985 VSS 0.0197f
C1231 VDD.n986 VSS 0.041f
C1232 VDD.n987 VSS 0.0659f
C1233 VDD.n988 VSS 0.0351f
C1234 VDD.n989 VSS 0.0351f
C1235 VDD.t3 VSS 0.287f
C1236 VDD.n990 VSS 0.00945f
C1237 VDD.n991 VSS 0.0093f
C1238 VDD.n992 VSS 0.0925f
C1239 VDD.n993 VSS 0.536f
C1240 VDD.t13 VSS 1.89f
C1241 VDD.n994 VSS 0.00945f
C1242 VDD.n995 VSS 0.0093f
C1243 VDD.n996 VSS 0.0925f
C1244 VDD.n997 VSS 0.00945f
C1245 VDD.n998 VSS 0.0093f
C1246 VDD.n999 VSS 0.0925f
C1247 VDD.n1000 VSS 1.21f
C1248 VDD.n1001 VSS 1.06f
C1249 VDD.t17 VSS 1.18f
C1250 VDD.n1002 VSS 1.81f
C1251 VDD.n1003 VSS 0.0316f
C1252 VDD.n1004 VSS 0.0316f
C1253 VDD.n1005 VSS 0.0326f
C1254 VDD.n1006 VSS 0.0326f
C1255 VDD.n1007 VSS 0.524f
C1256 VDD.t7 VSS 1.25f
C1257 VDD.n1008 VSS 2.04f
C1258 VDD.n1009 VSS 1.4f
C1259 VDD.n1010 VSS 0.287f
C1260 VDD.n1011 VSS 0.0378f
C1261 VDD.n1012 VSS 0.0415f
C1262 VDD.n1013 VSS 0.0546f
C1263 VDD.n1014 VSS 0.0116f
C1264 VDD.n1015 VSS 0.0197f
C1265 VDD.n1016 VSS 0.00315f
C1266 VDD.n1018 VSS 0.00315f
C1267 VDD.n1019 VSS 3.59e-19
C1268 VDD.n1020 VSS 0.00305f
C1269 VDD.n1021 VSS 0.0104f
C1270 VDD.n1022 VSS 0.00467f
C1271 VDD.n1023 VSS 0.00665f
C1272 VDD.n1024 VSS 0.00916f
C1273 VDD.n1025 VSS 0.00755f
C1274 VDD.n1026 VSS 0.00377f
C1275 VDD.n1027 VSS 0.0111f
C1276 VDD.n1028 VSS 0.0111f
C1277 VDD.n1029 VSS 0.0146f
C1278 VDD.n1031 VSS 0.0118f
C1279 VDD.n1032 VSS 3.59e-19
C1280 VDD.n1033 VSS 0.00395f
C1281 VDD.n1034 VSS 5.39e-19
C1282 VDD.n1035 VSS 0.00537f
C1283 VDD.n1036 VSS 0.00889f
C1284 VDD.n1037 VSS 0.00444f
C1285 VDD.n1038 VSS 0.011f
C1286 VDD.n1039 VSS 0.00683f
C1287 VDD.n1040 VSS 0.00661f
C1288 VDD.n1041 VSS 3.7e-19
C1289 VDD.n1042 VSS 0.00537f
C1290 VDD.n1043 VSS 5.39e-19
C1291 VDD.n1044 VSS 0.00395f
C1292 VDD.n1045 VSS 0.00305f
C1293 VDD.n1046 VSS 0.00377f
C1294 VDD.n1047 VSS 0.0111f
C1295 VDD.n1048 VSS 0.0111f
C1296 VDD.n1049 VSS 0.0146f
C1297 VDD.n1050 VSS 0.00315f
C1298 VDD.n1052 VSS 0.0118f
C1299 VDD.n1053 VSS 3.59e-19
C1300 VDD.n1054 VSS 0.00395f
C1301 VDD.n1055 VSS 5.39e-19
C1302 VDD.n1056 VSS 0.00537f
C1303 VDD.n1057 VSS 0.00889f
C1304 VDD.n1058 VSS 0.00444f
C1305 VDD.n1059 VSS 0.011f
C1306 VDD.n1060 VSS 0.00683f
C1307 VDD.n1061 VSS -0.0978f
C1308 VDD.n1062 VSS 3.7e-19
C1309 VDD.n1063 VSS 0.00537f
C1310 VDD.n1064 VSS 5.39e-19
C1311 VDD.n1065 VSS 0.00395f
C1312 VDD.n1066 VSS 0.00305f
C1313 VDD.n1067 VSS 0.00377f
C1314 VDD.n1068 VSS 0.0111f
C1315 VDD.n1069 VSS 0.0111f
C1316 VDD.n1070 VSS 0.0146f
C1317 VDD.n1071 VSS 0.00315f
C1318 VDD.n1073 VSS 0.0118f
C1319 VDD.n1074 VSS 3.59e-19
C1320 VDD.n1075 VSS 0.00395f
C1321 VDD.n1076 VSS 5.39e-19
C1322 VDD.n1077 VSS 0.00537f
C1323 VDD.n1078 VSS 0.00889f
C1324 VDD.n1079 VSS 0.00444f
C1325 VDD.n1080 VSS 0.011f
C1326 VDD.n1081 VSS 0.00683f
C1327 VDD.n1082 VSS -0.0856f
C1328 VDD.n1083 VSS 0.00377f
C1329 VDD.n1084 VSS 0.0493f
C1330 VDD.n1085 VSS 0.0499f
C1331 VDD.n1086 VSS 0.0443f
C1332 VDD.n1087 VSS 0.0443f
C1333 VDD.n1088 VSS 0.0453f
C1334 VDD.n1089 VSS 0.0281f
C1335 VDD.n1090 VSS 0.00658f
C1336 VDD.n1091 VSS -0.0981f
C1337 VDD.n1092 VSS 3.7e-19
C1338 VDD.n1093 VSS 0.00537f
C1339 VDD.n1094 VSS 5.39e-19
C1340 VDD.n1095 VSS 0.00395f
C1341 VDD.n1096 VSS 0.00305f
C1342 VDD.n1097 VSS 0.00377f
C1343 VDD.n1098 VSS 0.0111f
C1344 VDD.n1099 VSS 0.0111f
C1345 VDD.n1100 VSS 0.0146f
C1346 VDD.n1101 VSS 0.00315f
C1347 VDD.n1102 VSS 0.00305f
C1348 VDD.n1103 VSS 3.59e-19
C1349 VDD.n1104 VSS 0.0118f
C1350 VDD.n1105 VSS 0.00315f
C1351 VDD.n1106 VSS 0.00305f
C1352 VDD.n1107 VSS 0.0104f
C1353 VDD.n1108 VSS 0.00467f
C1354 VDD.n1109 VSS 0.00665f
C1355 VDD.n1110 VSS 0.00916f
C1356 VDD.n1111 VSS 0.00755f
C1357 VDD.n1112 VSS 0.00377f
C1358 VDD.n1113 VSS 0.0111f
C1359 VDD.n1114 VSS 0.0111f
C1360 VDD.n1115 VSS 0.0146f
C1361 VDD.n1116 VSS 0.0118f
C1362 VDD.n1117 VSS 3.59e-19
C1363 VDD.n1118 VSS 0.00395f
C1364 VDD.n1119 VSS 5.39e-19
C1365 VDD.n1120 VSS 0.00537f
C1366 VDD.n1121 VSS 0.00889f
C1367 VDD.n1122 VSS 0.00444f
C1368 VDD.n1123 VSS 0.0106f
C1369 VDD.n1124 VSS 0.00658f
C1370 VDD.n1125 VSS 0.00637f
C1371 VDD.n1126 VSS 3.7e-19
C1372 VDD.n1127 VSS 0.00537f
C1373 VDD.n1128 VSS 5.39e-19
C1374 VDD.n1129 VSS 0.00395f
C1375 VDD.n1130 VSS 0.00305f
C1376 VDD.n1131 VSS 0.00377f
C1377 VDD.n1132 VSS 0.0111f
C1378 VDD.n1133 VSS 0.0111f
C1379 VDD.n1134 VSS 0.0146f
C1380 VDD.n1135 VSS 0.00315f
C1381 VDD.n1136 VSS 0.00305f
C1382 VDD.n1137 VSS 3.59e-19
C1383 VDD.n1138 VSS 0.0118f
C1384 VDD.n1139 VSS 0.00315f
C1385 VDD.n1140 VSS 0.00305f
C1386 VDD.n1141 VSS 0.0104f
C1387 VDD.n1142 VSS 0.00467f
C1388 VDD.n1143 VSS 0.00665f
C1389 VDD.n1144 VSS 0.00916f
C1390 VDD.n1145 VSS 0.00755f
C1391 VDD.n1146 VSS 0.00377f
C1392 VDD.n1147 VSS 0.0111f
C1393 VDD.n1148 VSS 0.0111f
C1394 VDD.n1149 VSS 0.0146f
C1395 VDD.n1150 VSS 0.0118f
C1396 VDD.n1151 VSS 3.59e-19
C1397 VDD.n1152 VSS 0.00395f
C1398 VDD.n1153 VSS 5.39e-19
C1399 VDD.n1154 VSS 0.00537f
C1400 VDD.n1155 VSS 0.00889f
C1401 VDD.n1156 VSS 0.00444f
C1402 VDD.n1157 VSS 0.0106f
C1403 VDD.n1158 VSS 0.00658f
C1404 VDD.n1159 VSS 0.00637f
C1405 VDD.n1160 VSS 3.7e-19
C1406 VDD.n1161 VSS 0.00537f
C1407 VDD.n1162 VSS 5.39e-19
C1408 VDD.n1163 VSS 0.00395f
C1409 VDD.n1164 VSS 0.00305f
C1410 VDD.n1165 VSS 0.00377f
C1411 VDD.n1166 VSS 0.0111f
C1412 VDD.n1167 VSS 0.0111f
C1413 VDD.n1168 VSS 0.0146f
C1414 VDD.n1169 VSS 0.00315f
C1415 VDD.n1170 VSS 0.00305f
C1416 VDD.n1171 VSS 6e-19
C1417 VDD.n1172 VSS 0.00305f
C1418 VDD.n1173 VSS 0.00305f
C1419 VDD.n1174 VSS 0.00395f
C1420 VDD.n1175 VSS 0.0325f
C1421 VDD.n1176 VSS 0.0325f
C1422 VDD.n1177 VSS 0.0296f
C1423 VDD.n1178 VSS 0.00377f
C1424 VDD.n1179 VSS 0.0334f
C1425 VDD.n1180 VSS 0.00305f
C1426 VDD.n1181 VSS 6e-19
C1427 VDD.n1182 VSS 0.00395f
C1428 VDD.n1183 VSS 5.39e-19
C1429 VDD.n1184 VSS 0.00377f
C1430 VDD.n1185 VSS -0.0856f
C1431 VDD.n1186 VSS -0.241f
C1432 VDD.n1187 VSS 0.00665f
C1433 VDD.n1188 VSS 0.00916f
C1434 VDD.n1189 VSS 0.00755f
C1435 VDD.n1190 VSS 0.00377f
C1436 VDD.n1191 VSS 0.0111f
C1437 VDD.n1192 VSS 0.00305f
C1438 VDD.n1193 VSS 0.00315f
C1439 VDD.n1194 VSS 0.0118f
C1440 VDD.n1195 VSS 3.59e-19
C1441 VDD.n1196 VSS 0.00395f
C1442 VDD.n1197 VSS 5.39e-19
C1443 VDD.n1198 VSS 0.00377f
C1444 VDD.n1199 VSS 0.005f
C1445 VDD.n1200 VSS 0.00537f
C1446 VDD.n1201 VSS 0.00665f
C1447 VDD.n1202 VSS 0.00916f
C1448 VDD.n1203 VSS 0.00755f
C1449 VDD.n1204 VSS 0.00377f
C1450 VDD.n1205 VSS 0.0111f
C1451 VDD.n1206 VSS 0.00305f
C1452 VDD.n1207 VSS 3.59e-19
C1453 VDD.n1208 VSS 0.00395f
C1454 VDD.n1209 VSS 5.39e-19
C1455 VDD.n1210 VSS 0.00377f
C1456 VDD.n1211 VSS 0.005f
C1457 VDD.n1212 VSS 0.00537f
C1458 VDD.n1213 VSS 0.00665f
C1459 VDD.n1214 VSS 0.00916f
C1460 VDD.n1215 VSS 0.00755f
C1461 VDD.n1216 VSS 0.00377f
C1462 VDD.n1217 VSS 0.0111f
C1463 VDD.n1218 VSS 0.00305f
C1464 VDD.n1219 VSS 3.59e-19
C1465 VDD.n1220 VSS 0.00395f
C1466 VDD.n1221 VSS 5.39e-19
C1467 VDD.n1222 VSS 0.00377f
C1468 VDD.n1223 VSS -0.0856f
C1469 VDD.n1224 VSS -0.241f
C1470 VDD.n1225 VSS 0.00665f
C1471 VDD.n1226 VSS 0.00916f
C1472 VDD.n1227 VSS 0.00755f
C1473 VDD.n1228 VSS 0.00377f
C1474 VDD.n1229 VSS 0.0111f
C1475 VDD.n1230 VSS 0.00305f
C1476 VDD.n1231 VSS 3.59e-19
C1477 VDD.n1232 VSS 0.00395f
C1478 VDD.n1233 VSS 5.39e-19
C1479 VDD.n1234 VSS 0.00377f
C1480 VDD.n1235 VSS 0.005f
C1481 VDD.n1236 VSS 0.00537f
C1482 VDD.n1237 VSS 0.00665f
C1483 VDD.n1238 VSS 0.00916f
C1484 VDD.n1239 VSS 0.00755f
C1485 VDD.n1240 VSS 0.00377f
C1486 VDD.n1241 VSS 0.0111f
C1487 VDD.n1242 VSS 0.00305f
C1488 VDD.n1243 VSS 3.59e-19
C1489 VDD.n1244 VSS 0.00395f
C1490 VDD.n1245 VSS 5.39e-19
C1491 VDD.n1246 VSS 0.00377f
C1492 VDD.n1247 VSS 0.005f
C1493 VDD.n1248 VSS 0.00637f
C1494 VDD.n1249 VSS 0.00658f
C1495 VDD.n1250 VSS 0.0274f
C1496 VDD.n1251 VSS 0.0276f
C1497 VDD.n1252 VSS 0.028f
C1498 VDD.n1253 VSS 0.00658f
C1499 VDD.n1254 VSS -0.0981f
C1500 VDD.n1255 VSS 3.7e-19
C1501 VDD.n1256 VSS 0.00537f
C1502 VDD.n1257 VSS 5.39e-19
C1503 VDD.n1258 VSS 0.00395f
C1504 VDD.n1259 VSS 0.00305f
C1505 VDD.n1260 VSS 0.00377f
C1506 VDD.n1261 VSS 0.0111f
C1507 VDD.n1262 VSS 0.0111f
C1508 VDD.n1263 VSS 0.0146f
C1509 VDD.n1264 VSS 0.00315f
C1510 VDD.n1265 VSS 0.00305f
C1511 VDD.n1266 VSS 3.59e-19
C1512 VDD.n1267 VSS 0.0118f
C1513 VDD.n1268 VSS 0.00315f
C1514 VDD.n1269 VSS 0.00305f
C1515 VDD.n1270 VSS 0.0104f
C1516 VDD.n1271 VSS 0.00467f
C1517 VDD.n1272 VSS 0.00665f
C1518 VDD.n1273 VSS 0.00916f
C1519 VDD.n1274 VSS 0.00755f
C1520 VDD.n1275 VSS 0.00377f
C1521 VDD.n1276 VSS 0.0111f
C1522 VDD.n1277 VSS 0.0111f
C1523 VDD.n1278 VSS 0.0146f
C1524 VDD.n1279 VSS 0.0118f
C1525 VDD.n1280 VSS 3.59e-19
C1526 VDD.n1281 VSS 0.00395f
C1527 VDD.n1282 VSS 5.39e-19
C1528 VDD.n1283 VSS 0.00537f
C1529 VDD.n1284 VSS 0.00889f
C1530 VDD.n1285 VSS 0.00444f
C1531 VDD.n1286 VSS 0.0106f
C1532 VDD.n1287 VSS 0.00658f
C1533 VDD.n1288 VSS 0.00637f
C1534 VDD.n1289 VSS 3.7e-19
C1535 VDD.n1290 VSS 0.00537f
C1536 VDD.n1291 VSS 5.39e-19
C1537 VDD.n1292 VSS 0.00395f
C1538 VDD.n1293 VSS 0.00305f
C1539 VDD.n1294 VSS 0.00377f
C1540 VDD.n1295 VSS 0.0111f
C1541 VDD.n1296 VSS 0.0111f
C1542 VDD.n1297 VSS 0.0146f
C1543 VDD.n1298 VSS 0.00315f
C1544 VDD.n1299 VSS 0.00305f
C1545 VDD.n1300 VSS 3.59e-19
C1546 VDD.n1301 VSS 0.0118f
C1547 VDD.n1302 VSS 0.00315f
C1548 VDD.n1303 VSS 0.00305f
C1549 VDD.n1304 VSS 0.0104f
C1550 VDD.n1305 VSS 0.00467f
C1551 VDD.n1306 VSS 0.00665f
C1552 VDD.n1307 VSS 0.00916f
C1553 VDD.n1308 VSS 0.00755f
C1554 VDD.n1309 VSS 0.00377f
C1555 VDD.n1310 VSS 0.0111f
C1556 VDD.n1311 VSS 0.0111f
C1557 VDD.n1312 VSS 0.0146f
C1558 VDD.n1313 VSS 0.0118f
C1559 VDD.n1314 VSS 3.59e-19
C1560 VDD.n1315 VSS 0.00395f
C1561 VDD.n1316 VSS 5.39e-19
C1562 VDD.n1317 VSS 0.00537f
C1563 VDD.n1318 VSS 0.00889f
C1564 VDD.n1319 VSS 0.00444f
C1565 VDD.n1320 VSS 0.0106f
C1566 VDD.n1321 VSS 0.00658f
C1567 VDD.n1322 VSS 0.00637f
C1568 VDD.n1323 VSS 3.7e-19
C1569 VDD.n1324 VSS 0.00537f
C1570 VDD.n1325 VSS 5.39e-19
C1571 VDD.n1326 VSS 0.00395f
C1572 VDD.n1327 VSS 0.00305f
C1573 VDD.n1328 VSS 0.00377f
C1574 VDD.n1329 VSS 0.0111f
C1575 VDD.n1330 VSS 0.0111f
C1576 VDD.n1331 VSS 0.0146f
C1577 VDD.n1332 VSS 0.00315f
C1578 VDD.n1333 VSS 0.00305f
C1579 VDD.n1334 VSS 6e-19
C1580 VDD.n1335 VSS 0.00305f
C1581 VDD.n1336 VSS 0.00305f
C1582 VDD.n1337 VSS 0.00395f
C1583 VDD.n1338 VSS 0.0325f
C1584 VDD.n1339 VSS 0.0325f
C1585 VDD.n1340 VSS 0.0296f
C1586 VDD.n1341 VSS 0.00377f
C1587 VDD.n1342 VSS 0.0334f
C1588 VDD.n1343 VSS 0.00305f
C1589 VDD.n1344 VSS 6e-19
C1590 VDD.n1345 VSS 0.00395f
C1591 VDD.n1346 VSS 5.39e-19
C1592 VDD.n1347 VSS 0.00377f
C1593 VDD.n1348 VSS -0.0856f
C1594 VDD.n1349 VSS -0.241f
C1595 VDD.n1350 VSS 0.00665f
C1596 VDD.n1351 VSS 0.00916f
C1597 VDD.n1352 VSS 0.00755f
C1598 VDD.n1353 VSS 0.00377f
C1599 VDD.n1354 VSS 0.0111f
C1600 VDD.n1355 VSS 0.00305f
C1601 VDD.n1356 VSS 0.00315f
C1602 VDD.n1357 VSS 0.0118f
C1603 VDD.n1358 VSS 3.59e-19
C1604 VDD.n1359 VSS 0.00395f
C1605 VDD.n1360 VSS 5.39e-19
C1606 VDD.n1361 VSS 0.00377f
C1607 VDD.n1362 VSS 0.005f
C1608 VDD.n1363 VSS 0.00537f
C1609 VDD.n1364 VSS 0.00665f
C1610 VDD.n1365 VSS 0.00916f
C1611 VDD.n1366 VSS 0.00755f
C1612 VDD.n1367 VSS 0.00377f
C1613 VDD.n1368 VSS 0.0111f
C1614 VDD.n1369 VSS 0.00305f
C1615 VDD.n1370 VSS 3.59e-19
C1616 VDD.n1371 VSS 0.00395f
C1617 VDD.n1372 VSS 5.39e-19
C1618 VDD.n1373 VSS 0.00377f
C1619 VDD.n1374 VSS 0.005f
C1620 VDD.n1375 VSS 0.00537f
C1621 VDD.n1376 VSS 0.00665f
C1622 VDD.n1377 VSS 0.00916f
C1623 VDD.n1378 VSS 0.00755f
C1624 VDD.n1379 VSS 0.00377f
C1625 VDD.n1380 VSS 0.0111f
C1626 VDD.n1381 VSS 0.00305f
C1627 VDD.n1382 VSS 3.59e-19
C1628 VDD.n1383 VSS 0.00395f
C1629 VDD.n1384 VSS 5.39e-19
C1630 VDD.n1385 VSS 0.00377f
C1631 VDD.n1386 VSS -0.0856f
C1632 VDD.n1387 VSS -0.241f
C1633 VDD.n1388 VSS 0.00665f
C1634 VDD.n1389 VSS 0.00916f
C1635 VDD.n1390 VSS 0.00755f
C1636 VDD.n1391 VSS 0.00377f
C1637 VDD.n1392 VSS 0.0111f
C1638 VDD.n1393 VSS 0.00305f
C1639 VDD.n1394 VSS 3.59e-19
C1640 VDD.n1395 VSS 0.00395f
C1641 VDD.n1396 VSS 5.39e-19
C1642 VDD.n1397 VSS 0.00377f
C1643 VDD.n1398 VSS 0.005f
C1644 VDD.n1399 VSS 0.00537f
C1645 VDD.n1400 VSS 0.00665f
C1646 VDD.n1401 VSS 0.00916f
C1647 VDD.n1402 VSS 0.00755f
C1648 VDD.n1403 VSS 0.00377f
C1649 VDD.n1404 VSS 0.0111f
C1650 VDD.n1405 VSS 0.00305f
C1651 VDD.n1406 VSS 3.59e-19
C1652 VDD.n1407 VSS 0.00395f
C1653 VDD.n1408 VSS 5.39e-19
C1654 VDD.n1409 VSS 0.00377f
C1655 VDD.n1410 VSS 0.005f
C1656 VDD.n1411 VSS 0.00637f
C1657 VDD.n1412 VSS 0.00658f
C1658 VDD.n1413 VSS 0.0274f
C1659 VDD.n1414 VSS 0.0276f
C1660 VDD.n1415 VSS 0.028f
C1661 VDD.n1416 VSS 0.00658f
C1662 VDD.n1417 VSS -0.0981f
C1663 VDD.n1418 VSS 3.7e-19
C1664 VDD.n1419 VSS 0.00537f
C1665 VDD.n1420 VSS 5.39e-19
C1666 VDD.n1421 VSS 0.00395f
C1667 VDD.n1422 VSS 0.00305f
C1668 VDD.n1423 VSS 0.00377f
C1669 VDD.n1424 VSS 0.0111f
C1670 VDD.n1425 VSS 0.0111f
C1671 VDD.n1426 VSS 0.0146f
C1672 VDD.n1427 VSS 0.00315f
C1673 VDD.n1428 VSS 0.00305f
C1674 VDD.n1429 VSS 3.59e-19
C1675 VDD.n1430 VSS 0.0118f
C1676 VDD.n1431 VSS 0.00315f
C1677 VDD.n1432 VSS 0.00305f
C1678 VDD.n1433 VSS 0.0104f
C1679 VDD.n1434 VSS 0.00467f
C1680 VDD.n1435 VSS 0.00665f
C1681 VDD.n1436 VSS 0.00916f
C1682 VDD.n1437 VSS 0.00755f
C1683 VDD.n1438 VSS 0.00377f
C1684 VDD.n1439 VSS 0.0111f
C1685 VDD.n1440 VSS 0.0111f
C1686 VDD.n1441 VSS 0.0146f
C1687 VDD.n1442 VSS 0.0118f
C1688 VDD.n1443 VSS 3.59e-19
C1689 VDD.n1444 VSS 0.00395f
C1690 VDD.n1445 VSS 5.39e-19
C1691 VDD.n1446 VSS 0.00537f
C1692 VDD.n1447 VSS 0.00889f
C1693 VDD.n1448 VSS 0.00444f
C1694 VDD.n1449 VSS 0.0106f
C1695 VDD.n1450 VSS 0.00658f
C1696 VDD.n1451 VSS 0.00637f
C1697 VDD.n1452 VSS 3.7e-19
C1698 VDD.n1453 VSS 0.00537f
C1699 VDD.n1454 VSS 5.39e-19
C1700 VDD.n1455 VSS 0.00395f
C1701 VDD.n1456 VSS 0.00305f
C1702 VDD.n1457 VSS 0.00377f
C1703 VDD.n1458 VSS 0.0111f
C1704 VDD.n1459 VSS 0.0111f
C1705 VDD.n1460 VSS 0.0146f
C1706 VDD.n1461 VSS 0.00315f
C1707 VDD.n1462 VSS 0.00305f
C1708 VDD.n1463 VSS 3.59e-19
C1709 VDD.n1464 VSS 0.0118f
C1710 VDD.n1465 VSS 0.00315f
C1711 VDD.n1466 VSS 0.00305f
C1712 VDD.n1467 VSS 0.0104f
C1713 VDD.n1468 VSS 0.00467f
C1714 VDD.n1469 VSS 0.00665f
C1715 VDD.n1470 VSS 0.00916f
C1716 VDD.n1471 VSS 0.00755f
C1717 VDD.n1472 VSS 0.00377f
C1718 VDD.n1473 VSS 0.0111f
C1719 VDD.n1474 VSS 0.0111f
C1720 VDD.n1475 VSS 0.0146f
C1721 VDD.n1476 VSS 0.0118f
C1722 VDD.n1477 VSS 3.59e-19
C1723 VDD.n1478 VSS 0.00395f
C1724 VDD.n1479 VSS 5.39e-19
C1725 VDD.n1480 VSS 0.00537f
C1726 VDD.n1481 VSS 0.00889f
C1727 VDD.n1482 VSS 0.00444f
C1728 VDD.n1483 VSS 0.0106f
C1729 VDD.n1484 VSS 0.00658f
C1730 VDD.n1485 VSS 0.00637f
C1731 VDD.n1486 VSS 3.7e-19
C1732 VDD.n1487 VSS 0.00537f
C1733 VDD.n1488 VSS 5.39e-19
C1734 VDD.n1489 VSS 0.00395f
C1735 VDD.n1490 VSS 0.00305f
C1736 VDD.n1491 VSS 0.00377f
C1737 VDD.n1492 VSS 0.0111f
C1738 VDD.n1493 VSS 0.0111f
C1739 VDD.n1494 VSS 0.0146f
C1740 VDD.n1495 VSS 0.00315f
C1741 VDD.n1496 VSS 0.00305f
C1742 VDD.n1497 VSS 6e-19
C1743 VDD.n1498 VSS 0.00305f
C1744 VDD.n1499 VSS 0.00305f
C1745 VDD.n1500 VSS 0.00395f
C1746 VDD.n1501 VSS 0.0325f
C1747 VDD.n1502 VSS 0.0325f
C1748 VDD.n1503 VSS 0.0296f
C1749 VDD.n1504 VSS 0.00377f
C1750 VDD.n1505 VSS 0.0334f
C1751 VDD.n1506 VSS 0.00305f
C1752 VDD.n1507 VSS 6e-19
C1753 VDD.n1508 VSS 0.00395f
C1754 VDD.n1509 VSS 5.39e-19
C1755 VDD.n1510 VSS 0.00377f
C1756 VDD.n1511 VSS -0.0856f
C1757 VDD.n1512 VSS -0.241f
C1758 VDD.n1513 VSS 0.00665f
C1759 VDD.n1514 VSS 0.00916f
C1760 VDD.n1515 VSS 0.00755f
C1761 VDD.n1516 VSS 0.00377f
C1762 VDD.n1517 VSS 0.0111f
C1763 VDD.n1518 VSS 0.00305f
C1764 VDD.n1519 VSS 0.00315f
C1765 VDD.n1520 VSS 0.0118f
C1766 VDD.n1521 VSS 3.59e-19
C1767 VDD.n1522 VSS 0.00395f
C1768 VDD.n1523 VSS 5.39e-19
C1769 VDD.n1524 VSS 0.00377f
C1770 VDD.n1525 VSS 0.005f
C1771 VDD.n1526 VSS 0.00537f
C1772 VDD.n1527 VSS 0.00665f
C1773 VDD.n1528 VSS 0.00916f
C1774 VDD.n1529 VSS 0.00755f
C1775 VDD.n1530 VSS 0.00377f
C1776 VDD.n1531 VSS 0.0111f
C1777 VDD.n1532 VSS 0.00305f
C1778 VDD.n1533 VSS 3.59e-19
C1779 VDD.n1534 VSS 0.00395f
C1780 VDD.n1535 VSS 5.39e-19
C1781 VDD.n1536 VSS 0.00377f
C1782 VDD.n1537 VSS 0.005f
C1783 VDD.n1538 VSS 0.00537f
C1784 VDD.n1539 VSS 0.00665f
C1785 VDD.n1540 VSS 0.00916f
C1786 VDD.n1541 VSS 0.00755f
C1787 VDD.n1542 VSS 0.00377f
C1788 VDD.n1543 VSS 0.0111f
C1789 VDD.n1544 VSS 0.00305f
C1790 VDD.n1545 VSS 3.59e-19
C1791 VDD.n1546 VSS 0.00395f
C1792 VDD.n1547 VSS 5.39e-19
C1793 VDD.n1548 VSS 0.00377f
C1794 VDD.n1549 VSS -0.0856f
C1795 VDD.n1550 VSS -0.241f
C1796 VDD.n1551 VSS 0.00665f
C1797 VDD.n1552 VSS 0.00916f
C1798 VDD.n1553 VSS 0.00755f
C1799 VDD.n1554 VSS 0.00377f
C1800 VDD.n1555 VSS 0.0111f
C1801 VDD.n1556 VSS 0.00305f
C1802 VDD.n1557 VSS 3.59e-19
C1803 VDD.n1558 VSS 0.00395f
C1804 VDD.n1559 VSS 5.39e-19
C1805 VDD.n1560 VSS 0.00377f
C1806 VDD.n1561 VSS 0.005f
C1807 VDD.n1562 VSS 0.00537f
C1808 VDD.n1563 VSS 0.00665f
C1809 VDD.n1564 VSS 0.00916f
C1810 VDD.n1565 VSS 0.00755f
C1811 VDD.n1566 VSS 0.00377f
C1812 VDD.n1567 VSS 0.0111f
C1813 VDD.n1568 VSS 0.00305f
C1814 VDD.n1569 VSS 3.59e-19
C1815 VDD.n1570 VSS 0.00395f
C1816 VDD.n1571 VSS 5.39e-19
C1817 VDD.n1572 VSS 0.00377f
C1818 VDD.n1573 VSS 0.005f
C1819 VDD.n1574 VSS 0.00637f
C1820 VDD.n1575 VSS 0.00658f
C1821 VDD.n1576 VSS 0.0274f
C1822 VDD.n1577 VSS 0.0276f
C1823 VDD.n1578 VSS 0.028f
C1824 VDD.n1579 VSS 0.00658f
C1825 VDD.n1580 VSS -0.0981f
C1826 VDD.n1581 VSS 3.7e-19
C1827 VDD.n1582 VSS 0.00537f
C1828 VDD.n1583 VSS 5.39e-19
C1829 VDD.n1584 VSS 0.00395f
C1830 VDD.n1585 VSS 0.00305f
C1831 VDD.n1586 VSS 0.00377f
C1832 VDD.n1587 VSS 0.0111f
C1833 VDD.n1588 VSS 0.0111f
C1834 VDD.n1589 VSS 0.0146f
C1835 VDD.n1590 VSS 0.00315f
C1836 VDD.n1591 VSS 0.00305f
C1837 VDD.n1592 VSS 3.59e-19
C1838 VDD.n1593 VSS 0.0118f
C1839 VDD.n1594 VSS 0.00315f
C1840 VDD.n1595 VSS 0.00305f
C1841 VDD.n1596 VSS 0.0104f
C1842 VDD.n1597 VSS 0.00467f
C1843 VDD.n1598 VSS 0.00665f
C1844 VDD.n1599 VSS 0.00916f
C1845 VDD.n1600 VSS 0.00755f
C1846 VDD.n1601 VSS 0.00377f
C1847 VDD.n1602 VSS 0.0111f
C1848 VDD.n1603 VSS 0.0111f
C1849 VDD.n1604 VSS 0.0146f
C1850 VDD.n1605 VSS 0.0118f
C1851 VDD.n1606 VSS 3.59e-19
C1852 VDD.n1607 VSS 0.00395f
C1853 VDD.n1608 VSS 5.39e-19
C1854 VDD.n1609 VSS 0.00537f
C1855 VDD.n1610 VSS 0.00889f
C1856 VDD.n1611 VSS 0.00444f
C1857 VDD.n1612 VSS 0.0106f
C1858 VDD.n1613 VSS 0.00658f
C1859 VDD.n1614 VSS 0.00637f
C1860 VDD.n1615 VSS 3.7e-19
C1861 VDD.n1616 VSS 0.00537f
C1862 VDD.n1617 VSS 5.39e-19
C1863 VDD.n1618 VSS 0.00395f
C1864 VDD.n1619 VSS 0.00305f
C1865 VDD.n1620 VSS 0.00377f
C1866 VDD.n1621 VSS 0.0111f
C1867 VDD.n1622 VSS 0.0111f
C1868 VDD.n1623 VSS 0.0146f
C1869 VDD.n1624 VSS 0.00315f
C1870 VDD.n1625 VSS 0.00305f
C1871 VDD.n1626 VSS 3.59e-19
C1872 VDD.n1627 VSS 0.0118f
C1873 VDD.n1628 VSS 0.00315f
C1874 VDD.n1629 VSS 0.00305f
C1875 VDD.n1630 VSS 0.0104f
C1876 VDD.n1631 VSS 0.00467f
C1877 VDD.n1632 VSS 0.00665f
C1878 VDD.n1633 VSS 0.00916f
C1879 VDD.n1634 VSS 0.00755f
C1880 VDD.n1635 VSS 0.00377f
C1881 VDD.n1636 VSS 0.0111f
C1882 VDD.n1637 VSS 0.0111f
C1883 VDD.n1638 VSS 0.0146f
C1884 VDD.n1639 VSS 0.0118f
C1885 VDD.n1640 VSS 3.59e-19
C1886 VDD.n1641 VSS 0.00395f
C1887 VDD.n1642 VSS 5.39e-19
C1888 VDD.n1643 VSS 0.00537f
C1889 VDD.n1644 VSS 0.00889f
C1890 VDD.n1645 VSS 0.00444f
C1891 VDD.n1646 VSS 0.0106f
C1892 VDD.n1647 VSS 0.00658f
C1893 VDD.n1648 VSS 0.00637f
C1894 VDD.n1649 VSS 3.7e-19
C1895 VDD.n1650 VSS 0.00537f
C1896 VDD.n1651 VSS 5.39e-19
C1897 VDD.n1652 VSS 0.00395f
C1898 VDD.n1653 VSS 0.00305f
C1899 VDD.n1654 VSS 0.00377f
C1900 VDD.n1655 VSS 0.0111f
C1901 VDD.n1656 VSS 0.0111f
C1902 VDD.n1657 VSS 0.0146f
C1903 VDD.n1658 VSS 0.00315f
C1904 VDD.n1659 VSS 0.00305f
C1905 VDD.n1660 VSS 6e-19
C1906 VDD.n1661 VSS 0.00305f
C1907 VDD.n1662 VSS 0.00305f
C1908 VDD.n1663 VSS 0.00395f
C1909 VDD.n1664 VSS 0.0325f
C1910 VDD.n1665 VSS 0.0325f
C1911 VDD.n1666 VSS 0.0296f
C1912 VDD.n1667 VSS 0.00377f
C1913 VDD.n1668 VSS 0.0334f
C1914 VDD.n1669 VSS 0.00305f
C1915 VDD.n1670 VSS 6e-19
C1916 VDD.n1671 VSS 0.00395f
C1917 VDD.n1672 VSS 5.39e-19
C1918 VDD.n1673 VSS 0.00377f
C1919 VDD.n1674 VSS -0.0856f
C1920 VDD.n1675 VSS -0.241f
C1921 VDD.n1676 VSS 0.00665f
C1922 VDD.n1677 VSS 0.00916f
C1923 VDD.n1678 VSS 0.00755f
C1924 VDD.n1679 VSS 0.00377f
C1925 VDD.n1680 VSS 0.0111f
C1926 VDD.n1681 VSS 0.00305f
C1927 VDD.n1682 VSS 0.00315f
C1928 VDD.n1683 VSS 0.0118f
C1929 VDD.n1684 VSS 3.59e-19
C1930 VDD.n1685 VSS 0.00395f
C1931 VDD.n1686 VSS 0.0104f
C1932 VDD.n1687 VSS 0.00467f
C1933 VDD.n1688 VSS 0.00665f
C1934 VDD.n1689 VSS 0.00537f
C1935 VDD.n1690 VSS 0.00426f
C1936 VDD.n1691 VSS 0.00907f
C1937 VDD.n1692 VSS -0.214f
C1938 VDD.n1693 VSS -0.106f
C1939 VDD.n1694 VSS 0.00637f
C1940 VDD.n1695 VSS 0.005f
C1941 VDD.n1696 VSS 0.00377f
C1942 VDD.n1697 VSS 0.00467f
C1943 VDD.n1698 VSS 0.0104f
C1944 VDD.n1699 VSS 0.00755f
C1945 VDD.n1700 VSS 0.00916f
C1946 VDD.n1701 VSS 0.00395f
C1947 VDD.n1702 VSS 0.00305f
C1948 VDD.n1703 VSS 0.00395f
C1949 VDD.n1704 VSS 3.59e-19
C1950 VDD.n1705 VSS 0.0118f
C1951 VDD.n1706 VSS 2.89f
C1952 VDD.n1707 VSS 0.023f
C1953 VDD.n1708 VSS 0.0586f
C1954 VDD.n1709 VSS 0.0479f
C1955 VDD.n1710 VSS 0.0443f
C1956 VDD.n1711 VSS 0.0453f
C1957 VDD.n1712 VSS 0.00661f
C1958 VDD.n1713 VSS 0.175f
C1959 VDD.n1714 VSS 0.0123f
C1960 VDD.n1715 VSS 0.0987f
C1961 VDD.n1716 VSS 0.0987f
C1962 VDD.n1717 VSS 0.0123f
C1963 VDD.n1718 VSS 0.106f
C1964 VDD.n1719 VSS 0.106f
C1965 VDD.n1720 VSS 0.0123f
C1966 VDD.n1721 VSS 0.121f
C1967 VDD.n1722 VSS 0.121f
C1968 VDD.n1723 VSS 0.0123f
C1969 VDD.n1724 VSS 0.11f
C1970 VDD.n1725 VSS 0.052f
C1971 VDD.n1726 VSS 0.11f
C1972 VDD.n1727 VSS 0.0123f
C1973 VDD.n1728 VSS 0.00721f
C1974 VDD.n1729 VSS 0.0093f
C1975 VDD.n1730 VSS 0.0925f
C1976 VDD.n1731 VSS 0.823f
C1977 VDD.n1732 VSS 1.39f
C1978 VDD.t14 VSS 1.42f
C1979 VDD.n1733 VSS 1.27f
C1980 VDD.n1734 VSS 0.038f
C1981 VDD.n1735 VSS 0.038f
C1982 VDD.n1736 VSS 0.0393f
C1983 VDD.n1737 VSS 0.0589f
C1984 VDD.n1738 VSS 0.0366f
C1985 VDD.n1739 VSS 0.558f
C1986 VDD.n1740 VSS 0.61f
C1987 VDD.t11 VSS 0.142f
C1988 VDD.n1741 VSS 0.0719f
C1989 VDD.n1742 VSS 0.0357f
C1990 VDD.n1743 VSS 0.00867f
C1991 VDD.n1744 VSS 0.00444f
C1992 VDD.n1745 VSS 0.0163f
C1993 VDD.n1746 VSS 0.0221f
C1994 VDD.n1747 VSS 0.0311f
C1995 VDD.n1748 VSS 0.0196f
C1996 VDD.n1749 VSS 0.0225f
C1997 VDD.n1750 VSS 9.27e-19
C1998 VDD.n1751 VSS 0.0297f
C1999 VDD.n1752 VSS 0.0227f
C2000 VDD.n1753 VSS 0.0273f
C2001 VDD.n1754 VSS 0.00455f
C2002 VDD.n1755 VSS 0.0141f
C2003 VDD.n1756 VSS 0.00524f
C2004 VDD.n1757 VSS 0.00549f
C2005 VDD.n1758 VSS 0.00209f
C2006 VDD.n1759 VSS 0.00159f
C2007 VDD.n1760 VSS 0.0147f
C2008 VDD.n1761 VSS 0.00301f
C2009 VDD.n1762 VSS 0.00185f
C2010 VDD.n1763 VSS 0.017f
C2011 VDD.n1764 VSS 0.0859f
C2012 VDD.t5 VSS 0.117f
C2013 VDD.n1765 VSS 0.106f
C2014 VDD.n1766 VSS 0.023f
C2015 VDD.n1767 VSS 0.00867f
C2016 VDD.n1768 VSS 0.0588f
C2017 VDD.n1769 VSS 0.0163f
C2018 x5[7].floating.n0 VSS -7.97f
C2019 x5[7].floating.n1 VSS -28.8f
C2020 x5[7].floating.n2 VSS 3.82f
C2021 x5[7].floating.n3 VSS -7.06f
C2022 x5[7].floating.n4 VSS -28.3f
C2023 x5[7].floating.n5 VSS 52.6f
C2024 x5[7].floating.n6 VSS -28.3f
C2025 x5[7].floating.n7 VSS -7.06f
C2026 x5[7].floating.n8 VSS 3.82f
C2027 x5[7].floating.n9 VSS -28.8f
C2028 x5[7].floating.n10 VSS -8f
C2029 x5[7].floating.n11 VSS 2.2f
C2030 x5[7].floating.t5 VSS 0.857f
C2031 x5[7].floating.n12 VSS 6.64f
C2032 x5[7].floating.n13 VSS 1.21f
C2033 x5[7].floating.n14 VSS 1.16f
C2034 x5[7].floating.n15 VSS 2.18f
C2035 x5[7].floating.n16 VSS 1.06f
C2036 x5[7].floating.n17 VSS 0.365f
C2037 x5[7].floating.n18 VSS 1.06f
C2038 x5[7].floating.n19 VSS 2.8f
C2039 x5[7].floating.n20 VSS 51.3f
C2040 x5[7].floating.n21 VSS 2.78f
C2041 x5[7].floating.n22 VSS 1.06f
C2042 x5[7].floating.n23 VSS 0.363f
C2043 x5[7].floating.t2 VSS 0.857f
C2044 x5[7].floating.n24 VSS 6.47f
C2045 x5[7].floating.n25 VSS 1.15f
C2046 x5[7].floating.n26 VSS 1.36f
C2047 x5[7].floating.n27 VSS 2.2f
C2048 x5[7].floating.n28 VSS 1.06f
C2049 x5[7].floating.n29 VSS 2.22f
C2050 x5[7].floating.n30 VSS -7.97f
C2051 x5[7].floating.n31 VSS -28.8f
C2052 x5[7].floating.n32 VSS 3.82f
C2053 x5[7].floating.n33 VSS -7.06f
C2054 x5[7].floating.n34 VSS -28.3f
C2055 x5[7].floating.n35 VSS 52.6f
C2056 x5[7].floating.n36 VSS -28.3f
C2057 x5[7].floating.n37 VSS -7.06f
C2058 x5[7].floating.n38 VSS 3.82f
C2059 x5[7].floating.n39 VSS -28.8f
C2060 x5[7].floating.n40 VSS -8f
C2061 x5[7].floating.n41 VSS 2.2f
C2062 x5[7].floating.t1 VSS 0.857f
C2063 x5[7].floating.n42 VSS 6.64f
C2064 x5[7].floating.n43 VSS 1.21f
C2065 x5[7].floating.n44 VSS 1.16f
C2066 x5[7].floating.n45 VSS 2.18f
C2067 x5[7].floating.n46 VSS 1.06f
C2068 x5[7].floating.n47 VSS 0.365f
C2069 x5[7].floating.n48 VSS 1.06f
C2070 x5[7].floating.n49 VSS 2.8f
C2071 x5[7].floating.n50 VSS 51.3f
C2072 x5[7].floating.n51 VSS 2.78f
C2073 x5[7].floating.n52 VSS 1.06f
C2074 x5[7].floating.n53 VSS 0.363f
C2075 x5[7].floating.t3 VSS 0.857f
C2076 x5[7].floating.n54 VSS 6.47f
C2077 x5[7].floating.n55 VSS 1.15f
C2078 x5[7].floating.n56 VSS 1.36f
C2079 x5[7].floating.n57 VSS 2.2f
C2080 x5[7].floating.n58 VSS 1.06f
C2081 x5[7].floating.n59 VSS -15.2f
C2082 x5[7].floating.n60 VSS -15.1f
C2083 x5[7].floating.n61 VSS -41.5f
C2084 x5[7].floating.n62 VSS 0.765f
C2085 x5[7].floating.n63 VSS 2.46f
C2086 x5[7].floating.n64 VSS 51.4f
C2087 x5[7].floating.n65 VSS 2.46f
C2088 x5[7].floating.n66 VSS 0.765f
C2089 x5[7].floating.n67 VSS -33.4f
C2090 x5[7].floating.n68 VSS -4.55f
C2091 x5[7].floating.n69 VSS 3.82f
C2092 x5[7].floating.n70 VSS -28.8f
C2093 x5[7].floating.n71 VSS -7.06f
C2094 x5[7].floating.n72 VSS 2.68f
C2095 x5[7].floating.n73 VSS 51.9f
C2096 x5[7].floating.n74 VSS 3.23f
C2097 x5[7].floating.n75 VSS -7.82f
C2098 x5[7].floating.n76 VSS -28.8f
C2099 x5[7].floating.n77 VSS 3.82f
C2100 x5[7].floating.n78 VSS -5f
C2101 x5[7].floating.n79 VSS -32.9f
C2102 x5[7].floating.n80 VSS 0.765f
C2103 x5[7].floating.n81 VSS 2.46f
C2104 x5[7].floating.n82 VSS 2.68f
C2105 x5[7].floating.n83 VSS -7.06f
C2106 x5[7].floating.n84 VSS -28.8f
C2107 x5[7].floating.n85 VSS 3.82f
C2108 x5[7].floating.n86 VSS -4.55f
C2109 x5[7].floating.n87 VSS -33.4f
C2110 x5[7].floating.n88 VSS 0.765f
C2111 x5[7].floating.n89 VSS 2.46f
C2112 x5[7].floating.n90 VSS 51.4f
C2113 x5[7].floating.n91 VSS 51.3f
C2114 x5[7].floating.n92 VSS 2.8f
C2115 x5[7].floating.n93 VSS 1.06f
C2116 x5[7].floating.n94 VSS 0.365f
C2117 x5[7].floating.t7 VSS 0.857f
C2118 x5[7].floating.n95 VSS 6.64f
C2119 x5[7].floating.n96 VSS 1.21f
C2120 x5[7].floating.n97 VSS 1.16f
C2121 x5[7].floating.n98 VSS 2.18f
C2122 x5[7].floating.n99 VSS 1.06f
C2123 x5[7].floating.n100 VSS 2.2f
C2124 x5[7].floating.n101 VSS -8f
C2125 x5[7].floating.n102 VSS -28.8f
C2126 x5[7].floating.n103 VSS 3.82f
C2127 x5[7].floating.n104 VSS -7.06f
C2128 x5[7].floating.n105 VSS -28.3f
C2129 x5[7].floating.n106 VSS 2.78f
C2130 x5[7].floating.n107 VSS 1.06f
C2131 x5[7].floating.n108 VSS 0.363f
C2132 x5[7].floating.t6 VSS 0.857f
C2133 x5[7].floating.n109 VSS 6.47f
C2134 x5[7].floating.n110 VSS 1.15f
C2135 x5[7].floating.n111 VSS 1.36f
C2136 x5[7].floating.n112 VSS 2.2f
C2137 x5[7].floating.n113 VSS 1.06f
C2138 x5[7].floating.n114 VSS 2.22f
C2139 x5[7].floating.n115 VSS -7.97f
C2140 x5[7].floating.n116 VSS -28.8f
C2141 x5[7].floating.n117 VSS 3.82f
C2142 x5[7].floating.n118 VSS -7.06f
C2143 x5[7].floating.n119 VSS -28.3f
C2144 x5[7].floating.n120 VSS 52.6f
C2145 x5[7].floating.n121 VSS 51.9f
C2146 x5[7].floating.n122 VSS 3.23f
C2147 x5[7].floating.n123 VSS -7.82f
C2148 x5[7].floating.n124 VSS -28.8f
C2149 x5[7].floating.n125 VSS 3.82f
C2150 x5[7].floating.n126 VSS -5f
C2151 x5[7].floating.n127 VSS -32.9f
C2152 x5[7].floating.n128 VSS 0.765f
C2153 x5[7].floating.n129 VSS 2.46f
C2154 x5[7].floating.n130 VSS 51.4f
C2155 x5[7].floating.n131 VSS 2.46f
C2156 x5[7].floating.n132 VSS 0.765f
C2157 x5[7].floating.n133 VSS -33.4f
C2158 x5[7].floating.n134 VSS -4.55f
C2159 x5[7].floating.n135 VSS 3.82f
C2160 x5[7].floating.n136 VSS -28.8f
C2161 x5[7].floating.n137 VSS -7.06f
C2162 x5[7].floating.n138 VSS 2.68f
C2163 x5[7].floating.n139 VSS 51.9f
C2164 x5[7].floating.n140 VSS 3.23f
C2165 x5[7].floating.n141 VSS 2.22f
C2166 x5[7].floating.t4 VSS 0.857f
C2167 x5[7].floating.n142 VSS 6.47f
C2168 x5[7].floating.n143 VSS 1.15f
C2169 x5[7].floating.n144 VSS 1.36f
C2170 x5[7].floating.n145 VSS 2.2f
C2171 x5[7].floating.n146 VSS 1.06f
C2172 x5[7].floating.n147 VSS 0.363f
C2173 x5[7].floating.n148 VSS 1.06f
C2174 x5[7].floating.n149 VSS 2.78f
C2175 x5[7].floating.n150 VSS 51.3f
C2176 x5[7].floating.n151 VSS 2.8f
C2177 x5[7].floating.n152 VSS 1.06f
C2178 x5[7].floating.n153 VSS 0.365f
C2179 x5[7].floating.t0 VSS 0.857f
C2180 x5[7].floating.n154 VSS 7.14f
C2181 x5[7].floating.n155 VSS 1.21f
C2182 x5[7].floating.n156 VSS 1.16f
C2183 x5[7].floating.n157 VSS 1.67f
C2184 x5[7].floating.n158 VSS 1.06f
C2185 x5[7].floating.n159 VSS -17.3f
C2186 x5[7].floating.n160 VSS -17.2f
C2187 x5[7].floating.n161 VSS -43.5f
C2188 x5[7].floating.n162 VSS 0.765f
C2189 x5[7].floating.n163 VSS 2.46f
C2190 x5[7].floating.n164 VSS 51.4f
C2191 x5[7].floating.n165 VSS 2.46f
C2192 x5[7].floating.n166 VSS 0.765f
C2193 x5[7].floating.n167 VSS -32.9f
C2194 x5[7].floating.n168 VSS -5f
C2195 x5[7].floating.n169 VSS 3.82f
C2196 x5[7].floating.n170 VSS -28.8f
C2197 x5[7].floating.n171 VSS -7.82f
C2198 x10.Y.t1 VSS 0.0462f
C2199 x10.Y.t6 VSS 0.0167f
C2200 x10.Y.t8 VSS 0.0167f
C2201 x10.Y.t7 VSS 0.0167f
C2202 x10.Y.t2 VSS 0.0167f
C2203 x10.Y.t3 VSS 0.0167f
C2204 x10.Y.t4 VSS 0.0167f
C2205 x10.Y.t5 VSS 0.0167f
C2206 x10.Y.t9 VSS 0.0167f
C2207 x10.Y.n0 VSS 0.222f
C2208 x10.Y.n1 VSS 0.0366f
C2209 x10.Y.t0 VSS 0.0174f
C2210 x10.Y.n2 VSS 0.0188f
C2211 x10.Y.n3 VSS 0.0186f
C2212 x10.Y.n4 VSS 0.0151f
C2213 x10.Y.n5 VSS 0.0211f
.ends

