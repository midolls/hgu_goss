magic
tech sky130A
magscale 1 2
timestamp 1699109709
<< error_p >>
rect 917 1685 975 1691
rect 917 1651 929 1685
rect 917 1645 975 1651
<< nmos >>
rect 931 1723 961 1807
<< ndiff >>
rect 873 1795 931 1807
rect 873 1735 885 1795
rect 919 1735 931 1795
rect 873 1723 931 1735
rect 961 1723 1019 1807
<< ndiffc >>
rect 885 1735 919 1795
<< psubdiff >>
rect 540 598 872 614
rect 540 564 566 598
rect 600 564 646 598
rect 680 564 726 598
rect 760 564 806 598
rect 840 564 872 598
rect 540 546 872 564
<< psubdiffcont >>
rect 566 564 600 598
rect 646 564 680 598
rect 726 564 760 598
rect 806 564 840 598
<< poly >>
rect 931 1807 961 1833
rect 931 1701 961 1723
rect 913 1685 979 1701
rect 913 1651 929 1685
rect 963 1651 979 1685
rect 913 1635 979 1651
<< polycont >>
rect 929 1651 963 1685
<< locali >>
rect 885 1795 919 1811
rect 885 1719 919 1735
rect 913 1651 929 1685
rect 963 1651 979 1685
rect 540 598 872 614
rect 540 564 566 598
rect 600 564 646 598
rect 680 564 726 598
rect 760 564 806 598
rect 840 564 872 598
rect 540 546 872 564
<< viali >>
rect 885 1735 919 1795
rect 929 1651 963 1685
rect 566 564 600 598
rect 646 564 680 598
rect 726 564 760 598
rect 806 564 840 598
<< metal1 >>
rect 879 1797 925 1807
rect 857 1733 866 1797
rect 930 1733 939 1797
rect 857 1732 939 1733
rect 879 1723 925 1732
rect 917 1685 975 1691
rect 917 1651 929 1685
rect 963 1651 975 1685
rect 917 1645 975 1651
rect 540 608 872 614
rect 540 556 558 608
rect 610 556 638 608
rect 690 556 718 608
rect 770 556 798 608
rect 850 556 872 608
rect 540 546 872 556
<< via1 >>
rect 866 1795 930 1797
rect 866 1735 885 1795
rect 885 1735 919 1795
rect 919 1735 930 1795
rect 866 1733 930 1735
rect 558 598 610 608
rect 558 564 566 598
rect 566 564 600 598
rect 600 564 610 598
rect 558 556 610 564
rect 638 598 690 608
rect 638 564 646 598
rect 646 564 680 598
rect 680 564 690 598
rect 638 556 690 564
rect 718 598 770 608
rect 718 564 726 598
rect 726 564 760 598
rect 760 564 770 598
rect 718 556 770 564
rect 798 598 850 608
rect 798 564 806 598
rect 806 564 840 598
rect 840 564 850 598
rect 798 556 850 564
<< metal2 >>
rect 857 1733 866 1797
rect 930 1733 939 1797
rect 857 1732 939 1733
rect 540 610 872 614
rect 540 554 556 610
rect 612 554 636 610
rect 692 554 716 610
rect 772 554 796 610
rect 852 554 872 610
rect 540 546 872 554
<< via2 >>
rect 866 1733 930 1797
rect 556 608 612 610
rect 556 556 558 608
rect 558 556 610 608
rect 610 556 612 608
rect 556 554 612 556
rect 636 608 692 610
rect 636 556 638 608
rect 638 556 690 608
rect 690 556 692 608
rect 636 554 692 556
rect 716 608 772 610
rect 716 556 718 608
rect 718 556 770 608
rect 770 556 772 608
rect 716 554 772 556
rect 796 608 852 610
rect 796 556 798 608
rect 798 556 850 608
rect 850 556 852 608
rect 796 554 852 556
<< metal3 >>
rect 857 1797 939 1803
rect 857 1776 866 1797
rect 368 1774 866 1776
rect 930 1776 939 1797
rect 930 1774 1040 1776
rect 368 1710 472 1774
rect 536 1710 552 1774
rect 616 1710 632 1774
rect 696 1710 712 1774
rect 776 1710 792 1774
rect 856 1733 866 1774
rect 856 1710 872 1733
rect 936 1710 1040 1774
rect 368 1708 1040 1710
rect 368 1554 434 1708
rect 368 1490 369 1554
rect 433 1490 434 1554
rect 368 1474 434 1490
rect 368 1410 369 1474
rect 433 1410 434 1474
rect 368 1394 434 1410
rect 368 1330 369 1394
rect 433 1330 434 1394
rect 368 1314 434 1330
rect 368 1250 369 1314
rect 433 1250 434 1314
rect 368 1234 434 1250
rect 368 1170 369 1234
rect 433 1170 434 1234
rect 368 1154 434 1170
rect 368 1090 369 1154
rect 433 1090 434 1154
rect 368 1074 434 1090
rect 368 1010 369 1074
rect 433 1010 434 1074
rect 368 994 434 1010
rect 368 930 369 994
rect 433 930 434 994
rect 368 914 434 930
rect 368 850 369 914
rect 433 850 434 914
rect 368 834 434 850
rect 368 770 369 834
rect 433 770 434 834
rect 368 680 434 770
rect 494 676 554 1708
rect 614 616 674 1646
rect 734 676 794 1708
rect 854 616 914 1646
rect 974 1554 1040 1708
rect 974 1490 975 1554
rect 1039 1490 1040 1554
rect 974 1474 1040 1490
rect 974 1410 975 1474
rect 1039 1410 1040 1474
rect 974 1394 1040 1410
rect 974 1330 975 1394
rect 1039 1330 1040 1394
rect 974 1314 1040 1330
rect 974 1250 975 1314
rect 1039 1250 1040 1314
rect 974 1234 1040 1250
rect 974 1170 975 1234
rect 1039 1170 1040 1234
rect 974 1154 1040 1170
rect 974 1090 975 1154
rect 1039 1090 1040 1154
rect 974 1074 1040 1090
rect 974 1010 975 1074
rect 1039 1010 1040 1074
rect 974 994 1040 1010
rect 974 930 975 994
rect 1039 930 1040 994
rect 974 914 1040 930
rect 974 850 975 914
rect 1039 850 1040 914
rect 974 834 1040 850
rect 974 770 975 834
rect 1039 770 1040 834
rect 974 680 1040 770
rect 368 614 1040 616
rect 368 550 552 614
rect 616 550 632 614
rect 696 550 712 614
rect 776 550 792 614
rect 856 550 1040 614
rect 368 548 1040 550
<< via3 >>
rect 472 1710 536 1774
rect 552 1710 616 1774
rect 632 1710 696 1774
rect 712 1710 776 1774
rect 792 1710 856 1774
rect 872 1733 930 1774
rect 930 1733 936 1774
rect 872 1710 936 1733
rect 369 1490 433 1554
rect 369 1410 433 1474
rect 369 1330 433 1394
rect 369 1250 433 1314
rect 369 1170 433 1234
rect 369 1090 433 1154
rect 369 1010 433 1074
rect 369 930 433 994
rect 369 850 433 914
rect 369 770 433 834
rect 975 1490 1039 1554
rect 975 1410 1039 1474
rect 975 1330 1039 1394
rect 975 1250 1039 1314
rect 975 1170 1039 1234
rect 975 1090 1039 1154
rect 975 1010 1039 1074
rect 975 930 1039 994
rect 975 850 1039 914
rect 975 770 1039 834
rect 552 610 616 614
rect 552 554 556 610
rect 556 554 612 610
rect 612 554 616 610
rect 552 550 616 554
rect 632 610 696 614
rect 632 554 636 610
rect 636 554 692 610
rect 692 554 696 610
rect 632 550 696 554
rect 712 610 776 614
rect 712 554 716 610
rect 716 554 772 610
rect 772 554 776 610
rect 712 550 776 554
rect 792 610 856 614
rect 792 554 796 610
rect 796 554 852 610
rect 852 554 856 610
rect 792 550 856 554
<< metal4 >>
rect 368 1774 1040 1776
rect 368 1710 472 1774
rect 536 1710 552 1774
rect 616 1710 632 1774
rect 696 1710 712 1774
rect 776 1710 792 1774
rect 856 1710 872 1774
rect 936 1710 1040 1774
rect 368 1708 1040 1710
rect 368 1554 434 1708
rect 368 1490 369 1554
rect 433 1490 434 1554
rect 368 1474 434 1490
rect 368 1410 369 1474
rect 433 1410 434 1474
rect 368 1394 434 1410
rect 368 1330 369 1394
rect 433 1330 434 1394
rect 368 1314 434 1330
rect 368 1250 369 1314
rect 433 1250 434 1314
rect 368 1234 434 1250
rect 368 1170 369 1234
rect 433 1170 434 1234
rect 368 1154 434 1170
rect 368 1090 369 1154
rect 433 1090 434 1154
rect 368 1074 434 1090
rect 368 1010 369 1074
rect 433 1010 434 1074
rect 368 994 434 1010
rect 368 930 369 994
rect 433 930 434 994
rect 368 914 434 930
rect 368 850 369 914
rect 433 850 434 914
rect 368 834 434 850
rect 368 770 369 834
rect 433 770 434 834
rect 368 680 434 770
rect 494 616 554 1646
rect 614 676 674 1708
rect 734 616 794 1646
rect 854 676 914 1708
rect 974 1554 1040 1708
rect 974 1490 975 1554
rect 1039 1490 1040 1554
rect 974 1474 1040 1490
rect 974 1410 975 1474
rect 1039 1410 1040 1474
rect 974 1394 1040 1410
rect 974 1330 975 1394
rect 1039 1330 1040 1394
rect 974 1314 1040 1330
rect 974 1250 975 1314
rect 1039 1250 1040 1314
rect 974 1234 1040 1250
rect 974 1170 975 1234
rect 1039 1170 1040 1234
rect 974 1154 1040 1170
rect 974 1090 975 1154
rect 1039 1090 1040 1154
rect 974 1074 1040 1090
rect 974 1010 975 1074
rect 1039 1010 1040 1074
rect 974 994 1040 1010
rect 974 930 975 994
rect 1039 930 1040 994
rect 974 914 1040 930
rect 974 850 975 914
rect 1039 850 1040 914
rect 974 834 1040 850
rect 974 770 975 834
rect 1039 770 1040 834
rect 974 680 1040 770
rect 368 614 1040 616
rect 368 550 552 614
rect 616 550 632 614
rect 696 550 712 614
rect 776 550 792 614
rect 856 550 1040 614
rect 368 546 1040 550
<< labels >>
flabel metal1 929 1651 963 1685 0 FreeSans 320 0 0 0 SW
port 5 nsew
flabel ndiff 961 1723 1019 1807 0 FreeSans 320 0 0 0 delay_signal
port 7 nsew
flabel metal4 368 546 1040 614 0 FreeSans 320 0 0 0 CTOP
port 6 nsew
<< end >>
