* NGSPICE file created from hgu_clk_async_flat.ext - technology: sky130A

.subckt hgu_clk_async_RC async_clk_sar vdd vss sample_clk eob ready delay_offset     
+ async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[3]
+ async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[3]

X0 x4.x5[7].floating.t7 x4.x10.Y.t2 x4.x9.output_stack vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X1 x2.x9.output_stack async_setb_delay_ctrl_code[2].t0 x2.x4[3].floating vss.t42 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2 x4.x3[1].floating async_resetb_delay_ctrl_code[1].t0 x4.x9.output_stack vss.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X3 x10.Y x10.A vss.t38 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_1373_1841# eob.t0 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_2200_1841# sample_clk.t0 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 x4.x9.output_stack x4.x10.Y.t3 x4.x5[7].floating.t6 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X7 x9.Y x9.A vss.t45 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_n6207_n1487# ready.t0 a_n6295_n1487# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_n6207_n797# ready.t1 a_n6295_n935# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X10 a_n6182_1940# async_clk_sar.t2 a_n6270_2078# vdd.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X11 vss.t54 async_clk_sar.t3 a_n6207_n277# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X12 vss.t79 a_1771_1775# x3.X vss.t78 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_n397_1077# x4.x9.output_stack vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X14 x4.x9.output_stack async_resetb_delay_ctrl_code[2].t0 x4.x4[3].floating vss.t39 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X15 a_n6135_413# async_clk_sar.t4 a_n6207_413# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 vdd.t86 x9.Y a_1363_798# vdd.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X17 a_1307_1909# x3.X a_944_1775# vss.t28 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X18 a_818_1106# a_618_824# vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X19 a_618_824# x10.Y vss.t25 vss.t24 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X20 vss.t58 vdd.t96 a_2077_824# vss.t57 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X21 a_n397_736# x4.x9.output_stack x10.A vss.t62 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X22 a_2134_1909# x3.A0 a_1771_1775# vss.t77 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X23 a_1159_798# sample_clk.t1 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1403_1582# vss.t86 a_944_1775# vdd.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X25 a_n397_n2289# x9.A vss.t44 vdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X26 a_2230_1582# vss.t87 a_1771_1775# vdd.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X27 a_1094_1190# a_305_798# vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X28 a_1296_1190# a_1159_798# a_860_798# vdd.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 vss.t76 x9.Y a_724_824# vss.t75 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X30 vdd.t54 delay_offset.t0 x4.x6.SW vdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X31 a_618_824# x10.Y vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X32 a_n6207_n1# async_clk_sar.t5 a_n6295_n1# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X33 a_1363_798# a_1631_1008# a_1577_1106# vdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X34 x2.x4[3].floating async_setb_delay_ctrl_code[2].t1 x2.x9.output_stack vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X35 a_n6207_689# async_clk_sar.t6 a_n6295_551# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X36 vss.t6 a_944_1775# async_clk_sar.t0 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X37 a_n397_n1948# x2.x9.output_stack x9.A vss.t62 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X38 a_n6182_1664# async_clk_sar.t7 a_n6270_1526# vdd.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X39 a_210_798# a_305_798# vss.t17 vss.t16 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X40 a_n6182_n3152# ready.t2 a_n6270_n3014# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X41 a_944_1775# vss.t48 a_1086_1909# vss.t49 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X42 a_n397_1077# x10.A vss.t36 vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X43 a_n6135_n1073# ready.t3 a_n6207_n1073# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 vdd.t84 x9.Y a_305_798# vdd.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X45 x2.x4[3].floating async_setb_delay_ctrl_code[2].t2 x2.x9.output_stack vss.t40 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X46 a_n6207_n277# async_clk_sar.t8 a_n6295_n277# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X47 vss.t15 a_305_798# x27.Q_N vss.t14 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X48 a_n6135_n1349# ready.t4 a_n6207_n1349# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 x10.Y x10.A vdd.t35 vdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X50 vss.t43 x9.A a_n397_n2289# vdd.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X51 a_n6207_n1073# ready.t5 a_n6295_n1211# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X52 x2.x9.output_stack delay_offset.t1 x2.x7.floating vss.t59 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X53 x4.x10.Y.t0 async_resetb_delay_ctrl_code[3].t0 vss.t51 vss.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X54 a_210_798# a_305_798# vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X55 x4.x4[3].floating async_resetb_delay_ctrl_code[2].t1 x4.x9.output_stack vss.t40 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X56 x2.x9.output_stack ready.t6 a_n6270_n2738# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X57 vdd.t23 a_1373_1841# a_1403_1582# vdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X58 vdd.t13 a_305_798# x27.Q_N vdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X59 a_n6207_n1349# ready.t7 a_n6295_n1487# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X60 a_724_824# a_860_798# a_305_798# vss.t85 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X61 x4.x9.output_stack x4.x10.Y.t4 x4.x5[7].floating.t5 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X62 a_n397_n2289# x2.x9.output_stack vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X63 a_n6135_n139# async_clk_sar.t9 a_n6207_n139# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X64 a_2077_824# a_1159_798# a_1631_1008# vss.t21 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X65 a_n397_736# x4.x9.output_stack vss.t68 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X66 a_1159_798# sample_clk.t2 vss.t71 vss.t70 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 a_860_798# a_1159_798# a_1094_824# vss.t20 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X68 vss.t74 x9.Y a_1499_824# vss.t73 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X69 vss.t53 a_210_798# x3.A0 vss.t52 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X70 x2.x9.output_stack ready.t8 a_n6207_n1763# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X71 x4.x9.output_stack async_clk_sar.t10 a_n6207_689# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X72 a_1913_1909# sample_clk.t3 vss.t27 vss.t26 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X73 a_n6207_275# async_clk_sar.t11 a_n6295_275# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X74 a_2077_824# a_1158_1098# a_1631_1008# vdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 a_n6207_n1763# ready.t9 a_n6295_n1763# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X76 vss.t19 a_1159_798# a_1158_1098# vss.t18 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X77 a_305_798# a_618_824# a_724_824# vss.t30 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X78 a_n397_n1948# x2.x9.output_stack vss.t63 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X79 vss.t10 a_1363_798# a_1298_824# vss.t9 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X80 x4.x9.output_stack async_clk_sar.t12 a_n6270_1526# vdd.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X81 a_1086_1909# eob.t1 vss.t61 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X82 x4.x5[7].floating.t4 x4.x10.Y.t5 x4.x9.output_stack vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X83 x2.x9.output_stack x2.x6.SW x2.x6.floating vdd.t81 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X84 a_n6207_n139# async_clk_sar.t13 a_n6295_n277# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X85 x9.Y x9.A vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X86 vss.t56 delay_offset.t2 x4.x6.SW vss.t55 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X87 x4.x9.output_stack x4.x10.Y.t6 x4.x5[7].floating.t3 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X88 a_n6135_n1073# ready.t10 a_n6207_n935# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X89 vdd.t52 ready.t11 a_n6270_n3290# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X90 x2.x2.floating async_setb_delay_ctrl_code[0].t0 x2.x9.output_stack vss.t11 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X91 vdd.t93 a_1771_1775# x3.X vdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X92 a_1094_824# a_305_798# vss.t13 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X93 a_305_798# a_860_798# a_818_1106# vdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X94 x4.x9.output_stack x4.x6.SW x4.x6.floating vdd.t11 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X95 a_n6135_n139# async_clk_sar.t14 a_n6207_n1# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X96 vdd.t9 a_1363_798# a_1296_1190# vdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X97 vss.t81 delay_offset.t3 x2.x6.SW vss.t80 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X98 x2.x9.output_stack x2.x10.Y.t2 x2.x5[7].floating.t7 vdd.t63 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X99 a_n397_1077# x4.x9.output_stack x10.A vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X100 x4.x4[3].floating async_resetb_delay_ctrl_code[2].t2 x4.x9.output_stack vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X101 a_n397_n1948# x9.A vdd.t44 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X102 a_n6135_137# async_clk_sar.t15 a_n6207_275# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X103 a_n6182_1940# async_clk_sar.t16 a_n6270_1802# vdd.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X104 vdd.t3 a_2200_1841# a_2230_1582# vdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X105 a_1875_1190# a_1363_798# vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X106 x2.x9.output_stack x2.x10.Y.t3 x2.x5[7].floating.t6 vdd.t88 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X107 a_n6135_n1625# ready.t12 a_n6207_n1625# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X108 a_n6207_137# async_clk_sar.t17 a_n6295_n1# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X109 a_1577_1106# a_618_824# vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X110 vdd.t5 a_944_1775# async_clk_sar.t1 vdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X111 x4.x9.output_stack delay_offset.t4 x4.x7.floating vss.t59 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X112 x4.x9.output_stack async_resetb_delay_ctrl_code[1].t1 x4.x3[1].floating vss.t69 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X113 x2.x10.Y.t1 async_setb_delay_ctrl_code[3].t0 vss.t84 vss.t83 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X114 a_1298_824# a_1158_1098# a_860_798# vss.t65 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X115 a_n6182_n2876# ready.t13 a_n6270_n3014# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X116 a_n6207_n935# ready.t14 a_n6295_n935# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X117 a_1771_1775# x3.A0 a_1913_1582# vdd.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X118 a_n6207_n1625# ready.t15 a_n6295_n1763# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X119 vdd.t1 async_clk_sar.t18 a_n6270_2078# vdd.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X120 x2.x9.output_stack x2.x10.Y.t4 x2.x5[7].floating.t5 vdd.t40 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X121 a_1913_1582# sample_clk.t4 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X122 a_1499_824# a_1631_1008# a_1363_798# vss.t72 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X123 vdd.t43 x9.A a_n397_n1948# vss.t35 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X124 x4.x5[7].floating.t2 x4.x10.Y.t7 x4.x9.output_stack vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X125 x2.x9.output_stack x2.x10.Y.t5 x2.x5[7].floating.t4 vdd.t49 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X126 x4.x9.output_stack x4.x10.Y.t8 x4.x5[7].floating.t1 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X127 a_944_1775# x3.X a_1086_1582# vdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X128 a_n6207_551# async_clk_sar.t19 a_n6295_551# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X129 a_1086_1582# eob.t2 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X130 a_1363_798# a_618_824# a_1499_824# vss.t29 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X131 a_1631_1008# a_1159_798# a_1875_1190# vdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X132 a_n6135_137# async_clk_sar.t20 a_n6207_137# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X133 a_n6182_1664# async_clk_sar.t21 a_n6270_1802# vdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X134 a_n6135_n1349# ready.t16 a_n6207_n1211# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X135 a_1631_1008# a_1158_1098# a_1875_824# vss.t64 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X136 a_1875_824# a_1363_798# vss.t8 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X137 vdd.t34 x10.A a_n397_736# vss.t35 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X138 a_n6207_n1211# ready.t17 a_n6295_n1211# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X139 vdd.t19 a_1159_798# a_1158_1098# vdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X140 a_1373_1841# eob.t3 vss.t67 vss.t66 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X141 a_2200_1841# sample_clk.t5 vss.t32 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X142 a_n397_736# x10.A vdd.t33 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X143 a_n397_n2289# x2.x9.output_stack x9.A vdd.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X144 x4.x5[7].floating.t0 x4.x10.Y.t9 x4.x9.output_stack vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X145 x4.x9.output_stack async_resetb_delay_ctrl_code[2].t3 x4.x4[3].floating vss.t42 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X146 a_n6182_n2876# ready.t18 a_n6270_n2738# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X147 x2.x9.output_stack async_setb_delay_ctrl_code[1].t0 x2.x3[1].floating vss.t69 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X148 a_860_798# a_1158_1098# a_1094_1190# vdd.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X149 vdd.t90 delay_offset.t5 x2.x6.SW vdd.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X150 x2.x5[7].floating.t3 x2.x10.Y.t6 x2.x9.output_stack vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X151 a_n6135_413# async_clk_sar.t22 a_n6207_551# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X152 vss.t23 a_1373_1841# a_1307_1909# vss.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X153 a_1771_1775# vss.t46 a_1913_1909# vss.t47 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X154 vss.t4 a_2200_1841# a_2134_1909# vss.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X155 x2.x5[7].floating.t2 x2.x10.Y.t7 x2.x9.output_stack vdd.t78 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X156 x2.x5[7].floating.t1 x2.x10.Y.t8 x2.x9.output_stack vdd.t73 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X157 a_n6207_413# async_clk_sar.t23 a_n6295_275# vss.t0 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X158 x2.x10.Y.t0 async_setb_delay_ctrl_code[3].t1 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X159 vss.t82 ready.t19 a_n6207_n797# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 vdd.t50 a_210_798# x3.A0 vdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X161 vdd.t58 vdd.t56 a_2077_824# vdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X162 x2.x5[7].floating.t0 x2.x10.Y.t9 x2.x9.output_stack vdd.t94 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X163 x4.x2.floating async_resetb_delay_ctrl_code[0].t0 x4.x9.output_stack vss.t11 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X164 x4.x10.Y.t1 async_resetb_delay_ctrl_code[3].t1 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X165 a_n6182_n3152# ready.t20 a_n6270_n3290# vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X166 vss.t33 x10.A a_n397_1077# vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X167 x2.x9.output_stack async_setb_delay_ctrl_code[2].t3 x2.x4[3].floating vss.t39 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X168 x2.x3[1].floating async_setb_delay_ctrl_code[1].t1 x2.x9.output_stack vss.t2 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X169 a_n6135_n1625# ready.t21 a_n6207_n1487# vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
R0 x4.x10.Y x4.x10.Y.t9 154.847
R1 x4.x10.Y x4.x10.Y.t6 154.8
R2 x4.x10.Y x4.x10.Y.t5 154.8
R3 x4.x10.Y x4.x10.Y.t3 154.8
R4 x4.x10.Y x4.x10.Y.t2 154.8
R5 x4.x10.Y x4.x10.Y.t8 154.8
R6 x4.x10.Y x4.x10.Y.t7 154.8
R7 x4.x10.Y x4.x10.Y.t4 154.8
R8 x4.x10.Y.n0 x4.x10.Y 134.239
R9 x4.x10.Y x4.x10.Y.t0 106.635
R10 x4.x10.Y.n2 x4.x10.Y.t1 24.6567
R11 x4.x10.Y.n5 x4.x10.Y.n4 12.4089
R12 x4.x10.Y.n3 x4.x10.Y.n2 9.12522
R13 x4.x10.Y.n4 x4.x10.Y.n3 7.34048
R14 x4.x10.Y.n5 x4.x10.Y 2.22659
R15 x4.x10.Y.n2 x4.x10.Y.n1 1.93377
R16 x4.x10.Y x4.x10.Y.n5 1.55202
R17 x4.x10.Y.n3 x4.x10.Y.n0 0.69928
R18 x4.x5[7].floating.n154 x4.x5[7].floating.t5 68.0345
R19 x4.x5[7].floating.n142 x4.x5[7].floating.t2 68.0345
R20 x4.x5[7].floating.n12 x4.x5[7].floating.t1 68.0345
R21 x4.x5[7].floating.n24 x4.x5[7].floating.t7 68.0345
R22 x4.x5[7].floating.n54 x4.x5[7].floating.t4 68.0345
R23 x4.x5[7].floating.n72 x4.x5[7].floating.t3 68.0345
R24 x4.x5[7].floating.n84 x4.x5[7].floating.t0 68.0345
R25 x4.x5[7].floating.n42 x4.x5[7].floating.t6 68.0345
R26 x4.x5[7].floating.n103 x4.x5[7].floating.n65 0.660401
R27 x4.x5[7].floating.n112 x4.x5[7].floating.n50 0.660401
R28 x4.x5[7].floating.n121 x4.x5[7].floating.n35 0.660401
R29 x4.x5[7].floating.n130 x4.x5[7].floating.n20 0.660401
R30 x4.x5[7].floating.n139 x4.x5[7].floating.n5 0.660401
R31 x4.x5[7].floating.n90 x4.x5[7].floating.n89 0.320345
R32 x4.x5[7].floating.n160 x4.x5[7].floating.n159 0.308269
R33 x4.x5[7].floating.n161 x4.x5[7].floating.n160 0.173084
R34 x4.x5[7].floating.n91 x4.x5[7].floating.n90 0.162103
R35 x4.x5[7].floating.n160 x4.x5[7].floating 0.100688
R36 x4.x5[7].floating.n90 x4.x5[7].floating 0.0755007
R37 x4.x5[7].floating.n66 x4.x5[7].floating.n65 0.0716912
R38 x4.x5[7].floating.n65 x4.x5[7].floating.n64 0.0716912
R39 x4.x5[7].floating.n36 x4.x5[7].floating.n35 0.0716912
R40 x4.x5[7].floating.n35 x4.x5[7].floating.n34 0.0716912
R41 x4.x5[7].floating.n6 x4.x5[7].floating.n5 0.0716912
R42 x4.x5[7].floating.n5 x4.x5[7].floating.n4 0.0716912
R43 x4.x5[7].floating.n104 x4.x5[7].floating.n103 0.0716912
R44 x4.x5[7].floating.n122 x4.x5[7].floating.n121 0.0716912
R45 x4.x5[7].floating.n140 x4.x5[7].floating.n139 0.0716912
R46 x4.x5[7].floating.n70 x4.x5[7].floating.n69 0.0557941
R47 x4.x5[7].floating.n69 x4.x5[7].floating.n68 0.0557941
R48 x4.x5[7].floating.n68 x4.x5[7].floating.n67 0.0557941
R49 x4.x5[7].floating.n67 x4.x5[7].floating.n66 0.0557941
R50 x4.x5[7].floating.n64 x4.x5[7].floating.n63 0.0557941
R51 x4.x5[7].floating.n63 x4.x5[7].floating.n62 0.0557941
R52 x4.x5[7].floating.n62 x4.x5[7].floating.n61 0.0557941
R53 x4.x5[7].floating.n61 x4.x5[7].floating.n60 0.0557941
R54 x4.x5[7].floating.n40 x4.x5[7].floating.n39 0.0557941
R55 x4.x5[7].floating.n39 x4.x5[7].floating.n38 0.0557941
R56 x4.x5[7].floating.n38 x4.x5[7].floating.n37 0.0557941
R57 x4.x5[7].floating.n37 x4.x5[7].floating.n36 0.0557941
R58 x4.x5[7].floating.n34 x4.x5[7].floating.n33 0.0557941
R59 x4.x5[7].floating.n33 x4.x5[7].floating.n32 0.0557941
R60 x4.x5[7].floating.n32 x4.x5[7].floating.n31 0.0557941
R61 x4.x5[7].floating.n31 x4.x5[7].floating.n30 0.0557941
R62 x4.x5[7].floating.n10 x4.x5[7].floating.n9 0.0557941
R63 x4.x5[7].floating.n9 x4.x5[7].floating.n8 0.0557941
R64 x4.x5[7].floating.n8 x4.x5[7].floating.n7 0.0557941
R65 x4.x5[7].floating.n7 x4.x5[7].floating.n6 0.0557941
R66 x4.x5[7].floating.n4 x4.x5[7].floating.n3 0.0557941
R67 x4.x5[7].floating.n3 x4.x5[7].floating.n2 0.0557941
R68 x4.x5[7].floating.n2 x4.x5[7].floating.n1 0.0557941
R69 x4.x5[7].floating.n1 x4.x5[7].floating.n0 0.0557941
R70 x4.x5[7].floating.n99 x4.x5[7].floating.n98 0.0557941
R71 x4.x5[7].floating.n100 x4.x5[7].floating.n99 0.0557941
R72 x4.x5[7].floating.n101 x4.x5[7].floating.n100 0.0557941
R73 x4.x5[7].floating.n102 x4.x5[7].floating.n101 0.0557941
R74 x4.x5[7].floating.n106 x4.x5[7].floating.n105 0.0557941
R75 x4.x5[7].floating.n107 x4.x5[7].floating.n106 0.0557941
R76 x4.x5[7].floating.n108 x4.x5[7].floating.n107 0.0557941
R77 x4.x5[7].floating.n117 x4.x5[7].floating.n116 0.0557941
R78 x4.x5[7].floating.n118 x4.x5[7].floating.n117 0.0557941
R79 x4.x5[7].floating.n119 x4.x5[7].floating.n118 0.0557941
R80 x4.x5[7].floating.n120 x4.x5[7].floating.n119 0.0557941
R81 x4.x5[7].floating.n124 x4.x5[7].floating.n123 0.0557941
R82 x4.x5[7].floating.n125 x4.x5[7].floating.n124 0.0557941
R83 x4.x5[7].floating.n126 x4.x5[7].floating.n125 0.0557941
R84 x4.x5[7].floating.n135 x4.x5[7].floating.n134 0.0557941
R85 x4.x5[7].floating.n136 x4.x5[7].floating.n135 0.0557941
R86 x4.x5[7].floating.n137 x4.x5[7].floating.n136 0.0557941
R87 x4.x5[7].floating.n138 x4.x5[7].floating.n137 0.0557941
R88 x4.x5[7].floating.n171 x4.x5[7].floating.n170 0.0557941
R89 x4.x5[7].floating.n170 x4.x5[7].floating.n169 0.0557941
R90 x4.x5[7].floating.n169 x4.x5[7].floating.n168 0.0557941
R91 x4.x5[7].floating.n95 x4.x5[7].floating.n94 0.0537206
R92 x4.x5[7].floating.n113 x4.x5[7].floating.n112 0.0537206
R93 x4.x5[7].floating.n131 x4.x5[7].floating.n130 0.0537206
R94 x4.x5[7].floating.n164 x4.x5[7].floating.n163 0.0537206
R95 x4.x5[7].floating.n94 x4.x5[7].floating.n93 0.0530294
R96 x4.x5[7].floating.n112 x4.x5[7].floating.n111 0.0530294
R97 x4.x5[7].floating.n130 x4.x5[7].floating.n129 0.0530294
R98 x4.x5[7].floating.n165 x4.x5[7].floating.n164 0.0530294
R99 x4.x5[7].floating.n80 x4.x5[7].floating.n79 0.0529559
R100 x4.x5[7].floating.n50 x4.x5[7].floating.n49 0.0529559
R101 x4.x5[7].floating.n20 x4.x5[7].floating.n19 0.0529559
R102 x4.x5[7].floating.n151 x4.x5[7].floating.n150 0.0529559
R103 x4.x5[7].floating.n81 x4.x5[7].floating.n80 0.0524559
R104 x4.x5[7].floating.n51 x4.x5[7].floating.n50 0.0524559
R105 x4.x5[7].floating.n21 x4.x5[7].floating.n20 0.0524559
R106 x4.x5[7].floating.n150 x4.x5[7].floating.n149 0.0524559
R107 x4.x5[7].floating.n109 x4.x5[7].floating.n108 0.0523382
R108 x4.x5[7].floating.n127 x4.x5[7].floating.n126 0.0523382
R109 x4.x5[7].floating.n168 x4.x5[7].floating.n167 0.0523382
R110 x4.x5[7].floating.n98 x4.x5[7].floating.n97 0.0516471
R111 x4.x5[7].floating.n116 x4.x5[7].floating.n115 0.0516471
R112 x4.x5[7].floating.n134 x4.x5[7].floating.n133 0.0516471
R113 x4.x5[7].floating.n103 x4.x5[7].floating 0.0495735
R114 x4.x5[7].floating.n121 x4.x5[7].floating 0.0495735
R115 x4.x5[7].floating.n139 x4.x5[7].floating 0.0495735
R116 x4.x5[7].floating.n157 x4.x5[7].floating.n156 0.0408846
R117 x4.x5[7].floating.n15 x4.x5[7].floating.n14 0.0408846
R118 x4.x5[7].floating.n75 x4.x5[7].floating.n74 0.0408846
R119 x4.x5[7].floating.n45 x4.x5[7].floating.n44 0.0408846
R120 x4.x5[7].floating.n105 x4.x5[7].floating 0.0336765
R121 x4.x5[7].floating.n123 x4.x5[7].floating 0.0336765
R122 x4.x5[7].floating x4.x5[7].floating.n171 0.0336765
R123 x4.x5[7].floating.n60 x4.x5[7].floating.n59 0.0271618
R124 x4.x5[7].floating.n30 x4.x5[7].floating.n29 0.0271618
R125 x4.x5[7].floating.n71 x4.x5[7].floating.n70 0.0266618
R126 x4.x5[7].floating.n41 x4.x5[7].floating.n40 0.0266618
R127 x4.x5[7].floating.n11 x4.x5[7].floating.n10 0.0266618
R128 x4.x5[7].floating x4.x5[7].floating.n102 0.0226176
R129 x4.x5[7].floating x4.x5[7].floating.n104 0.0226176
R130 x4.x5[7].floating x4.x5[7].floating.n120 0.0226176
R131 x4.x5[7].floating x4.x5[7].floating.n122 0.0226176
R132 x4.x5[7].floating x4.x5[7].floating.n138 0.0226176
R133 x4.x5[7].floating x4.x5[7].floating.n140 0.0226176
R134 x4.x5[7].floating.n93 x4.x5[7].floating.n92 0.0191618
R135 x4.x5[7].floating.n111 x4.x5[7].floating.n110 0.0191618
R136 x4.x5[7].floating.n129 x4.x5[7].floating.n128 0.0191618
R137 x4.x5[7].floating.n166 x4.x5[7].floating.n165 0.0191618
R138 x4.x5[7].floating.n96 x4.x5[7].floating.n95 0.0184706
R139 x4.x5[7].floating.n114 x4.x5[7].floating.n113 0.0184706
R140 x4.x5[7].floating.n132 x4.x5[7].floating.n131 0.0184706
R141 x4.x5[7].floating.n163 x4.x5[7].floating.n162 0.0184706
R142 x4.x5[7].floating.n82 x4.x5[7].floating.n81 0.014
R143 x4.x5[7].floating.n76 x4.x5[7].floating.n71 0.014
R144 x4.x5[7].floating.n52 x4.x5[7].floating.n51 0.014
R145 x4.x5[7].floating.n46 x4.x5[7].floating.n41 0.014
R146 x4.x5[7].floating.n22 x4.x5[7].floating.n21 0.014
R147 x4.x5[7].floating.n16 x4.x5[7].floating.n11 0.014
R148 x4.x5[7].floating.n149 x4.x5[7].floating.n148 0.014
R149 x4.x5[7].floating.n159 x4.x5[7].floating.n158 0.014
R150 x4.x5[7].floating.n89 x4.x5[7].floating.n88 0.0135
R151 x4.x5[7].floating.n79 x4.x5[7].floating.n78 0.0135
R152 x4.x5[7].floating.n59 x4.x5[7].floating.n58 0.0135
R153 x4.x5[7].floating.n49 x4.x5[7].floating.n48 0.0135
R154 x4.x5[7].floating.n29 x4.x5[7].floating.n28 0.0135
R155 x4.x5[7].floating.n19 x4.x5[7].floating.n18 0.0135
R156 x4.x5[7].floating.n146 x4.x5[7].floating.n141 0.0135
R157 x4.x5[7].floating.n152 x4.x5[7].floating.n151 0.0135
R158 x4.x5[7].floating.n145 x4.x5[7].floating.n144 0.0120385
R159 x4.x5[7].floating.n27 x4.x5[7].floating.n26 0.0120385
R160 x4.x5[7].floating.n57 x4.x5[7].floating.n56 0.0120385
R161 x4.x5[7].floating.n87 x4.x5[7].floating.n86 0.0120385
R162 x4.x5[7].floating.n97 x4.x5[7].floating.n96 0.00464706
R163 x4.x5[7].floating.n115 x4.x5[7].floating.n114 0.00464706
R164 x4.x5[7].floating.n133 x4.x5[7].floating.n132 0.00464706
R165 x4.x5[7].floating.n162 x4.x5[7].floating.n161 0.00464706
R166 x4.x5[7].floating.n92 x4.x5[7].floating.n91 0.00395588
R167 x4.x5[7].floating.n110 x4.x5[7].floating.n109 0.00395588
R168 x4.x5[7].floating.n128 x4.x5[7].floating.n127 0.00395588
R169 x4.x5[7].floating.n167 x4.x5[7].floating.n166 0.00395588
R170 x4.x5[7].floating.n143 x4.x5[7].floating.n142 0.00359614
R171 x4.x5[7].floating.n25 x4.x5[7].floating.n24 0.00359614
R172 x4.x5[7].floating.n55 x4.x5[7].floating.n54 0.00359614
R173 x4.x5[7].floating.n85 x4.x5[7].floating.n84 0.00359614
R174 x4.x5[7].floating.n88 x4.x5[7].floating.n83 0.0035
R175 x4.x5[7].floating.n78 x4.x5[7].floating.n77 0.0035
R176 x4.x5[7].floating.n58 x4.x5[7].floating.n53 0.0035
R177 x4.x5[7].floating.n48 x4.x5[7].floating.n47 0.0035
R178 x4.x5[7].floating.n28 x4.x5[7].floating.n23 0.0035
R179 x4.x5[7].floating.n18 x4.x5[7].floating.n17 0.0035
R180 x4.x5[7].floating.n147 x4.x5[7].floating.n146 0.0035
R181 x4.x5[7].floating.n153 x4.x5[7].floating.n152 0.0035
R182 x4.x5[7].floating.n83 x4.x5[7].floating.n82 0.003
R183 x4.x5[7].floating.n77 x4.x5[7].floating.n76 0.003
R184 x4.x5[7].floating.n53 x4.x5[7].floating.n52 0.003
R185 x4.x5[7].floating.n47 x4.x5[7].floating.n46 0.003
R186 x4.x5[7].floating.n23 x4.x5[7].floating.n22 0.003
R187 x4.x5[7].floating.n17 x4.x5[7].floating.n16 0.003
R188 x4.x5[7].floating.n148 x4.x5[7].floating.n147 0.003
R189 x4.x5[7].floating.n158 x4.x5[7].floating.n153 0.003
R190 x4.x5[7].floating.n155 x4.x5[7].floating.n154 0.00277942
R191 x4.x5[7].floating.n43 x4.x5[7].floating.n42 0.0023396
R192 x4.x5[7].floating.n13 x4.x5[7].floating.n12 0.0023396
R193 x4.x5[7].floating.n73 x4.x5[7].floating.n72 0.0023396
R194 x4.x5[7].floating.n157 x4.x5[7].floating.n155 0.00233747
R195 x4.x5[7].floating.n15 x4.x5[7].floating.n13 0.00200689
R196 x4.x5[7].floating.n75 x4.x5[7].floating.n73 0.00200689
R197 x4.x5[7].floating.n45 x4.x5[7].floating.n43 0.00200689
R198 x4.x5[7].floating.n145 x4.x5[7].floating.n143 0.0010233
R199 x4.x5[7].floating.n27 x4.x5[7].floating.n25 0.0010233
R200 x4.x5[7].floating.n57 x4.x5[7].floating.n55 0.0010233
R201 x4.x5[7].floating.n87 x4.x5[7].floating.n85 0.0010233
R202 x4.x5[7].floating.n88 x4.x5[7].floating.n87 0.00053972
R203 x4.x5[7].floating.n76 x4.x5[7].floating.n75 0.00053972
R204 x4.x5[7].floating.n58 x4.x5[7].floating.n57 0.00053972
R205 x4.x5[7].floating.n28 x4.x5[7].floating.n27 0.00053972
R206 x4.x5[7].floating.n16 x4.x5[7].floating.n15 0.00053972
R207 x4.x5[7].floating.n146 x4.x5[7].floating.n145 0.00053972
R208 x4.x5[7].floating.n158 x4.x5[7].floating.n157 0.00053972
R209 x4.x5[7].floating.n46 x4.x5[7].floating.n45 0.00053972
R210 vdd.n2677 vdd.n2508 13300
R211 vdd.t32 vdd 6325.98
R212 vdd.n2812 vdd.n2508 3575.45
R213 vdd vdd.n2508 1986.36
R214 vdd.n696 vdd.t48 1761.46
R215 vdd.n2604 vdd.n2572 556.851
R216 vdd.n2524 vdd.t30 500.865
R217 vdd.n2713 vdd.n2528 440.25
R218 vdd.n2807 vdd.n2755 426
R219 vdd.n2577 vdd.t58 371
R220 vdd.n669 vdd.t45 361.541
R221 vdd.n2793 vdd.n2790 351
R222 vdd.n2575 vdd.n2574 337.3
R223 vdd.n2635 vdd.n2631 337.3
R224 vdd.t56 vdd.n2591 331.51
R225 vdd.t51 vdd 325.205
R226 vdd.n2585 vdd.n2579 308.598
R227 vdd.n2568 vdd.n2567 304.122
R228 vdd.n2667 vdd.n2666 302.438
R229 vdd.n1829 vdd.t89 258.856
R230 vdd.t53 vdd.n2808 258.856
R231 vdd.n2810 vdd 242.981
R232 vdd.n2721 vdd.n2519 233.143
R233 vdd.n2534 vdd.t14 212.315
R234 vdd.n2592 vdd.t56 210.692
R235 vdd.n2591 vdd.t96 209.403
R236 vdd.n2705 vdd.n2519 202.286
R237 vdd.n1676 vdd.n77 198.234
R238 vdd.n699 vdd.n698 198.234
R239 vdd.n3482 vdd.n3481 198.118
R240 vdd.n3256 vdd.n3255 198.118
R241 vdd.n3030 vdd.n3029 198.118
R242 vdd.n2482 vdd.n2481 198.118
R243 vdd.n3032 vdd.n3031 198.118
R244 vdd.n3258 vdd.n3257 198.118
R245 vdd.n3484 vdd.n3483 198.118
R246 vdd.n1827 vdd.t64 188.965
R247 vdd.t66 vdd.n2791 188.965
R248 vdd.n1701 vdd.n64 185
R249 vdd.n1705 vdd.n64 185
R250 vdd.n50 vdd.n49 185
R251 vdd.n49 vdd.n48 185
R252 vdd.n1731 vdd.n1730 185
R253 vdd.n1730 vdd.n1729 185
R254 vdd.n29 vdd.n28 185
R255 vdd.n1760 vdd.n29 185
R256 vdd.n1783 vdd.n1782 185
R257 vdd.n1784 vdd.n1783 185
R258 vdd.n1781 vdd.n15 185
R259 vdd.n1785 vdd.n15 185
R260 vdd.n1763 vdd.n1762 185
R261 vdd.n1762 vdd.n1761 185
R262 vdd.n1732 vdd.n31 185
R263 vdd.n31 vdd.n30 185
R264 vdd.n1726 vdd.n1725 185
R265 vdd.n1727 vdd.n1726 185
R266 vdd.n1846 vdd.n1845 185
R267 vdd.n1847 vdd.n1846 185
R268 vdd.n16 vdd.n14 185
R269 vdd.n1848 vdd.n16 185
R270 vdd.n1703 vdd.n1702 185
R271 vdd.n1704 vdd.n1703 185
R272 vdd.n594 vdd.n592 185
R273 vdd.n724 vdd.n594 185
R274 vdd.n747 vdd.n746 185
R275 vdd.n748 vdd.n747 185
R276 vdd.n566 vdd.n565 185
R277 vdd.n565 vdd.n564 185
R278 vdd.n781 vdd.n780 185
R279 vdd.n780 vdd.n779 185
R280 vdd.n801 vdd.n800 185
R281 vdd.n802 vdd.n801 185
R282 vdd.n838 vdd.n529 185
R283 vdd.n842 vdd.n529 185
R284 vdd.n516 vdd.n515 185
R285 vdd.n515 vdd.n514 185
R286 vdd.n868 vdd.n867 185
R287 vdd.n867 vdd.n866 185
R288 vdd.n500 vdd.n499 185
R289 vdd.n887 vdd.n500 185
R290 vdd.n937 vdd.n936 185
R291 vdd.n938 vdd.n937 185
R292 vdd.n475 vdd.n474 185
R293 vdd.n947 vdd.n475 185
R294 vdd.n460 vdd.n458 185
R295 vdd.n975 vdd.n460 185
R296 vdd.n998 vdd.n997 185
R297 vdd.n999 vdd.n998 185
R298 vdd.n432 vdd.n431 185
R299 vdd.n431 vdd.n430 185
R300 vdd.n1032 vdd.n1031 185
R301 vdd.n1031 vdd.n1030 185
R302 vdd.n1052 vdd.n1051 185
R303 vdd.n1053 vdd.n1052 185
R304 vdd.n1089 vdd.n395 185
R305 vdd.n1093 vdd.n395 185
R306 vdd.n382 vdd.n381 185
R307 vdd.n381 vdd.n380 185
R308 vdd.n1119 vdd.n1118 185
R309 vdd.n1118 vdd.n1117 185
R310 vdd.n366 vdd.n365 185
R311 vdd.n1138 vdd.n366 185
R312 vdd.n1188 vdd.n1187 185
R313 vdd.n1189 vdd.n1188 185
R314 vdd.n341 vdd.n340 185
R315 vdd.n1198 vdd.n341 185
R316 vdd.n326 vdd.n324 185
R317 vdd.n1226 vdd.n326 185
R318 vdd.n1249 vdd.n1248 185
R319 vdd.n1250 vdd.n1249 185
R320 vdd.n298 vdd.n297 185
R321 vdd.n297 vdd.n296 185
R322 vdd.n1283 vdd.n1282 185
R323 vdd.n1282 vdd.n1281 185
R324 vdd.n1303 vdd.n1302 185
R325 vdd.n1304 vdd.n1303 185
R326 vdd.n1340 vdd.n261 185
R327 vdd.n1344 vdd.n261 185
R328 vdd.n248 vdd.n247 185
R329 vdd.n247 vdd.n246 185
R330 vdd.n1370 vdd.n1369 185
R331 vdd.n1369 vdd.n1368 185
R332 vdd.n232 vdd.n231 185
R333 vdd.n1389 vdd.n232 185
R334 vdd.n1439 vdd.n1438 185
R335 vdd.n1440 vdd.n1439 185
R336 vdd.n207 vdd.n206 185
R337 vdd.n1449 vdd.n207 185
R338 vdd.n192 vdd.n190 185
R339 vdd.n1477 vdd.n192 185
R340 vdd.n1500 vdd.n1499 185
R341 vdd.n1501 vdd.n1500 185
R342 vdd.n164 vdd.n163 185
R343 vdd.n163 vdd.n162 185
R344 vdd.n1534 vdd.n1533 185
R345 vdd.n1533 vdd.n1532 185
R346 vdd.n1554 vdd.n1553 185
R347 vdd.n1555 vdd.n1554 185
R348 vdd.n1586 vdd.n128 185
R349 vdd.n1590 vdd.n128 185
R350 vdd.n114 vdd.n113 185
R351 vdd.n113 vdd.n112 185
R352 vdd.n1616 vdd.n1615 185
R353 vdd.n1615 vdd.n1614 185
R354 vdd.n93 vdd.n92 185
R355 vdd.n1645 vdd.n93 185
R356 vdd.n1673 vdd.n1672 185
R357 vdd.n1674 vdd.n1673 185
R358 vdd.n1671 vdd.n78 185
R359 vdd.n1675 vdd.n78 185
R360 vdd.n1648 vdd.n1647 185
R361 vdd.n1647 vdd.n1646 185
R362 vdd.n1617 vdd.n95 185
R363 vdd.n95 vdd.n94 185
R364 vdd.n1611 vdd.n1610 185
R365 vdd.n1612 vdd.n1611 185
R366 vdd.n1677 vdd.n79 185
R367 vdd.n1588 vdd.n1587 185
R368 vdd.n1589 vdd.n1588 185
R369 vdd.n161 vdd.n160 185
R370 vdd.n1531 vdd.n161 185
R371 vdd.n1505 vdd.n1504 185
R372 vdd.n1504 vdd.n1503 185
R373 vdd.n181 vdd.n180 185
R374 vdd.n180 vdd.n179 185
R375 vdd.n1475 vdd.n1474 185
R376 vdd.n1476 vdd.n1475 185
R377 vdd.n147 vdd.n146 185
R378 vdd.n1556 vdd.n147 185
R379 vdd.n1452 vdd.n1451 185
R380 vdd.n1451 vdd.n1450 185
R381 vdd.n1437 vdd.n212 185
R382 vdd.n1441 vdd.n212 185
R383 vdd.n1392 vdd.n1391 185
R384 vdd.n1391 vdd.n1390 185
R385 vdd.n1371 vdd.n234 185
R386 vdd.n234 vdd.n233 185
R387 vdd.n1365 vdd.n1364 185
R388 vdd.n1366 vdd.n1365 185
R389 vdd.n1447 vdd.n1446 185
R390 vdd.n1448 vdd.n1447 185
R391 vdd.n1445 vdd.n209 185
R392 vdd.n209 vdd.n208 185
R393 vdd.n1342 vdd.n1341 185
R394 vdd.n1343 vdd.n1342 185
R395 vdd.n295 vdd.n294 185
R396 vdd.n1280 vdd.n295 185
R397 vdd.n1254 vdd.n1253 185
R398 vdd.n1253 vdd.n1252 185
R399 vdd.n315 vdd.n314 185
R400 vdd.n314 vdd.n313 185
R401 vdd.n1224 vdd.n1223 185
R402 vdd.n1225 vdd.n1224 185
R403 vdd.n281 vdd.n280 185
R404 vdd.n1305 vdd.n281 185
R405 vdd.n1201 vdd.n1200 185
R406 vdd.n1200 vdd.n1199 185
R407 vdd.n1186 vdd.n346 185
R408 vdd.n1190 vdd.n346 185
R409 vdd.n1141 vdd.n1140 185
R410 vdd.n1140 vdd.n1139 185
R411 vdd.n1120 vdd.n368 185
R412 vdd.n368 vdd.n367 185
R413 vdd.n1114 vdd.n1113 185
R414 vdd.n1115 vdd.n1114 185
R415 vdd.n1196 vdd.n1195 185
R416 vdd.n1197 vdd.n1196 185
R417 vdd.n1194 vdd.n343 185
R418 vdd.n343 vdd.n342 185
R419 vdd.n1091 vdd.n1090 185
R420 vdd.n1092 vdd.n1091 185
R421 vdd.n429 vdd.n428 185
R422 vdd.n1029 vdd.n429 185
R423 vdd.n1003 vdd.n1002 185
R424 vdd.n1002 vdd.n1001 185
R425 vdd.n449 vdd.n448 185
R426 vdd.n448 vdd.n447 185
R427 vdd.n973 vdd.n972 185
R428 vdd.n974 vdd.n973 185
R429 vdd.n415 vdd.n414 185
R430 vdd.n1054 vdd.n415 185
R431 vdd.n950 vdd.n949 185
R432 vdd.n949 vdd.n948 185
R433 vdd.n935 vdd.n480 185
R434 vdd.n939 vdd.n480 185
R435 vdd.n890 vdd.n889 185
R436 vdd.n889 vdd.n888 185
R437 vdd.n869 vdd.n502 185
R438 vdd.n502 vdd.n501 185
R439 vdd.n863 vdd.n862 185
R440 vdd.n864 vdd.n863 185
R441 vdd.n945 vdd.n944 185
R442 vdd.n946 vdd.n945 185
R443 vdd.n943 vdd.n477 185
R444 vdd.n477 vdd.n476 185
R445 vdd.n840 vdd.n839 185
R446 vdd.n841 vdd.n840 185
R447 vdd.n563 vdd.n562 185
R448 vdd.n778 vdd.n563 185
R449 vdd.n752 vdd.n751 185
R450 vdd.n751 vdd.n750 185
R451 vdd.n722 vdd.n721 185
R452 vdd.n723 vdd.n722 185
R453 vdd.n583 vdd.n582 185
R454 vdd.n582 vdd.n581 185
R455 vdd.n549 vdd.n548 185
R456 vdd.n803 vdd.n549 185
R457 vdd.n697 vdd.n608 185
R458 vdd.n3737 vdd.n3736 185
R459 vdd.n1921 vdd.n1920 185
R460 vdd.n1910 vdd.n1909 185
R461 vdd.n1899 vdd.n1898 185
R462 vdd.n1888 vdd.n1887 185
R463 vdd.n3756 vdd.n3755 185
R464 vdd.n3756 vdd.n1886 185
R465 vdd.n3775 vdd.n3774 185
R466 vdd.n3775 vdd.n1886 185
R467 vdd.n3794 vdd.n3793 185
R468 vdd.n3794 vdd.n1886 185
R469 vdd.n3813 vdd.n3812 185
R470 vdd.n1885 vdd.n1884 185
R471 vdd.n3719 vdd.n1932 185
R472 vdd.n2835 vdd.n2834 185
R473 vdd.n2438 vdd.n2437 185
R474 vdd.n2884 vdd.n2883 185
R475 vdd.n2903 vdd.n2425 185
R476 vdd.n2921 vdd.n2920 185
R477 vdd.n2940 vdd.n2390 185
R478 vdd.n2939 vdd.n2393 185
R479 vdd.n2943 vdd.n2392 185
R480 vdd.n2391 vdd.n2376 185
R481 vdd.n2979 vdd.n2978 185
R482 vdd.n2976 vdd.n2375 185
R483 vdd.n3006 vdd.n3005 185
R484 vdd.n3008 vdd.n2357 185
R485 vdd.n3027 vdd.n3026 185
R486 vdd.n2347 vdd.n2346 185
R487 vdd.n3033 vdd.n2345 185
R488 vdd.n2319 vdd.n2318 185
R489 vdd.n2304 vdd.n2303 185
R490 vdd.n3110 vdd.n3109 185
R491 vdd.n3129 vdd.n2291 185
R492 vdd.n3147 vdd.n3146 185
R493 vdd.n3166 vdd.n2256 185
R494 vdd.n3165 vdd.n2259 185
R495 vdd.n3169 vdd.n2258 185
R496 vdd.n2257 vdd.n2242 185
R497 vdd.n3205 vdd.n3204 185
R498 vdd.n3202 vdd.n2241 185
R499 vdd.n3232 vdd.n3231 185
R500 vdd.n3234 vdd.n2223 185
R501 vdd.n3253 vdd.n3252 185
R502 vdd.n2213 vdd.n2212 185
R503 vdd.n3259 vdd.n2211 185
R504 vdd.n2185 vdd.n2184 185
R505 vdd.n2170 vdd.n2169 185
R506 vdd.n3336 vdd.n3335 185
R507 vdd.n3355 vdd.n2157 185
R508 vdd.n3373 vdd.n3372 185
R509 vdd.n3392 vdd.n2122 185
R510 vdd.n3391 vdd.n2125 185
R511 vdd.n3395 vdd.n2124 185
R512 vdd.n2123 vdd.n2108 185
R513 vdd.n3431 vdd.n3430 185
R514 vdd.n3428 vdd.n2107 185
R515 vdd.n3458 vdd.n3457 185
R516 vdd.n3460 vdd.n2089 185
R517 vdd.n3479 vdd.n3478 185
R518 vdd.n2079 vdd.n2078 185
R519 vdd.n3485 vdd.n2077 185
R520 vdd.n2051 vdd.n2050 185
R521 vdd.n2036 vdd.n2035 185
R522 vdd.n3562 vdd.n3561 185
R523 vdd.n3581 vdd.n2023 185
R524 vdd.n3599 vdd.n3598 185
R525 vdd.n3618 vdd.n1988 185
R526 vdd.n3617 vdd.n1991 185
R527 vdd.n3621 vdd.n1990 185
R528 vdd.n1989 vdd.n1974 185
R529 vdd.n3657 vdd.n3656 185
R530 vdd.n3654 vdd.n1973 185
R531 vdd.n3684 vdd.n3683 185
R532 vdd.n3686 vdd.n1955 185
R533 vdd.n3710 vdd.n3709 185
R534 vdd.n1944 vdd.n1943 185
R535 vdd.n3579 vdd.n3578 185
R536 vdd.n3559 vdd.n2034 185
R537 vdd.n3534 vdd.n3533 185
R538 vdd.n3513 vdd.n3512 185
R539 vdd.n3600 vdd.n2003 185
R540 vdd.n2062 vdd.n2061 185
R541 vdd.n3353 vdd.n3352 185
R542 vdd.n3333 vdd.n2168 185
R543 vdd.n3308 vdd.n3307 185
R544 vdd.n3287 vdd.n3286 185
R545 vdd.n3374 vdd.n2137 185
R546 vdd.n2196 vdd.n2195 185
R547 vdd.n3127 vdd.n3126 185
R548 vdd.n3107 vdd.n2302 185
R549 vdd.n3082 vdd.n3081 185
R550 vdd.n3061 vdd.n3060 185
R551 vdd.n3148 vdd.n2271 185
R552 vdd.n2330 vdd.n2329 185
R553 vdd.n2901 vdd.n2900 185
R554 vdd.n2881 vdd.n2436 185
R555 vdd.n2856 vdd.n2855 185
R556 vdd.n2922 vdd.n2405 185
R557 vdd.n2833 vdd.n2453 185
R558 vdd.n2790 vdd.n2789 185
R559 vdd.n2791 vdd.n2790 185
R560 vdd.n2533 vdd.n2523 174.857
R561 vdd.n2625 vdd.n2552 173.143
R562 vdd.n672 vdd.n671 172.5
R563 vdd.n2609 vdd.n2572 168
R564 vdd.n2604 vdd.n2573 168
R565 vdd.n2620 vdd.n2564 166.286
R566 vdd.n2719 vdd.n2522 166.286
R567 vdd.n2538 vdd.n2537 165.252
R568 vdd.n2647 vdd.n2565 164.571
R569 vdd.n2634 vdd.n2632 160.918
R570 vdd.n1788 vdd 160.49
R571 vdd.n2792 vdd 160.49
R572 vdd.n2643 vdd.n2565 159.429
R573 vdd.n2674 vdd.n2551 157.714
R574 vdd.n2679 vdd.n2551 157.714
R575 vdd.n2609 vdd.n2566 154.286
R576 vdd.n2518 vdd.t35 152.88
R577 vdd.n2795 vdd.t67 152.88
R578 vdd.n666 vdd.t46 152.879
R579 vdd.n1786 vdd.t90 152.879
R580 vdd.n1791 vdd.t65 152.879
R581 vdd.n2772 vdd.t54 152.879
R582 vdd.n2647 vdd.n2564 152.571
R583 vdd.n2719 vdd.n2523 152.571
R584 vdd.n2643 vdd.n2625 150.857
R585 vdd.n2674 vdd.n2552 150.857
R586 vdd.n2679 vdd.n2522 147.429
R587 vdd.n2536 vdd.n2533 145.714
R588 vdd.n2620 vdd.n2566 144
R589 vdd.n2582 vdd.n2573 142.286
R590 vdd.n698 vdd.t68 141.692
R591 vdd.n2613 vdd.n2612 137.606
R592 vdd.n2550 vdd.n2549 137.606
R593 vdd.n667 vdd.n664 137.135
R594 vdd.n2707 vdd.n2536 128.571
R595 vdd.n2622 vdd.n2621 123.692
R596 vdd.n2612 vdd.t37 123.496
R597 vdd.n2549 vdd.t72 123.496
R598 vdd.t75 vdd.t57 118.591
R599 vdd vdd.t81 116.731
R600 vdd vdd.n669 115.751
R601 vdd.n2792 vdd.t66 113.897
R602 vdd.t76 vdd.n2645 112.216
R603 vdd.n2644 vdd.n2624 112.216
R604 vdd.n1592 vdd.n128 111.177
R605 vdd.n1611 vdd.n111 111.177
R606 vdd.n1643 vdd.n95 111.177
R607 vdd.n1647 vdd.n81 111.177
R608 vdd.n1679 vdd.n78 111.177
R609 vdd.n1475 vdd.n194 111.177
R610 vdd.n1479 vdd.n180 111.177
R611 vdd.n1504 vdd.n178 111.177
R612 vdd.n1529 vdd.n161 111.177
R613 vdd.n1554 vdd.n149 111.177
R614 vdd.n1346 vdd.n261 111.177
R615 vdd.n1365 vdd.n245 111.177
R616 vdd.n1387 vdd.n234 111.177
R617 vdd.n1391 vdd.n214 111.177
R618 vdd.n1443 vdd.n212 111.177
R619 vdd.n1224 vdd.n328 111.177
R620 vdd.n1228 vdd.n314 111.177
R621 vdd.n1253 vdd.n312 111.177
R622 vdd.n1278 vdd.n295 111.177
R623 vdd.n1303 vdd.n283 111.177
R624 vdd.n1095 vdd.n395 111.177
R625 vdd.n1114 vdd.n379 111.177
R626 vdd.n1136 vdd.n368 111.177
R627 vdd.n1140 vdd.n348 111.177
R628 vdd.n1192 vdd.n346 111.177
R629 vdd.n973 vdd.n462 111.177
R630 vdd.n977 vdd.n448 111.177
R631 vdd.n1002 vdd.n446 111.177
R632 vdd.n1027 vdd.n429 111.177
R633 vdd.n1052 vdd.n417 111.177
R634 vdd.n844 vdd.n529 111.177
R635 vdd.n863 vdd.n513 111.177
R636 vdd.n885 vdd.n502 111.177
R637 vdd.n889 vdd.n482 111.177
R638 vdd.n941 vdd.n480 111.177
R639 vdd.n722 vdd.n596 111.177
R640 vdd.n726 vdd.n582 111.177
R641 vdd.n751 vdd.n580 111.177
R642 vdd.n776 vdd.n563 111.177
R643 vdd.n801 vdd.n551 111.177
R644 vdd.n1707 vdd.n64 111.177
R645 vdd.n1726 vdd.n47 111.177
R646 vdd.n1758 vdd.n31 111.177
R647 vdd.n1762 vdd.n18 111.177
R648 vdd.n1850 vdd.n15 111.177
R649 vdd.n3652 vdd.n1974 111.177
R650 vdd.n3688 vdd.n3686 111.177
R651 vdd.n3512 vdd.n3510 111.177
R652 vdd.n3533 vdd.n3531 111.177
R653 vdd.n3559 vdd.n3558 111.177
R654 vdd.n3579 vdd.n2024 111.177
R655 vdd.n3426 vdd.n2108 111.177
R656 vdd.n3462 vdd.n3460 111.177
R657 vdd.n3286 vdd.n3284 111.177
R658 vdd.n3307 vdd.n3305 111.177
R659 vdd.n3333 vdd.n3332 111.177
R660 vdd.n3353 vdd.n2158 111.177
R661 vdd.n3200 vdd.n2242 111.177
R662 vdd.n3236 vdd.n3234 111.177
R663 vdd.n3060 vdd.n3058 111.177
R664 vdd.n3081 vdd.n3079 111.177
R665 vdd.n3107 vdd.n3106 111.177
R666 vdd.n3127 vdd.n2292 111.177
R667 vdd.n2974 vdd.n2376 111.177
R668 vdd.n3010 vdd.n3008 111.177
R669 vdd.n2855 vdd.n2853 111.177
R670 vdd.n2881 vdd.n2880 111.177
R671 vdd.n2901 vdd.n2426 111.177
R672 vdd.n3739 vdd.n3737 111.177
R673 vdd.n3758 vdd.n3756 111.177
R674 vdd.n3777 vdd.n3775 111.177
R675 vdd.n3796 vdd.n3794 111.177
R676 vdd.n2809 vdd.t53 108.719
R677 vdd.t21 vdd.t74 107.115
R678 vdd.n2646 vdd.t82 104.564
R679 vdd.n2675 vdd.t26 96.9133
R680 vdd.n671 vdd.n668 92.5005
R681 vdd.n671 vdd.n670 92.5005
R682 vdd.n673 vdd.n672 92.5005
R683 vdd.n1839 vdd.n1838 92.5005
R684 vdd.n1840 vdd.n1839 92.5005
R685 vdd.n1790 vdd.n1789 92.5005
R686 vdd.n1789 vdd.n1788 92.5005
R687 vdd.n2584 vdd.n2573 92.5005
R688 vdd.n2580 vdd.n2573 92.5005
R689 vdd.n2553 vdd.n2552 92.5005
R690 vdd.n2623 vdd.n2552 92.5005
R691 vdd.n2627 vdd.n2625 92.5005
R692 vdd.n2625 vdd.n2624 92.5005
R693 vdd.n2643 vdd.n2642 92.5005
R694 vdd.n2644 vdd.n2643 92.5005
R695 vdd.n2636 vdd.n2565 92.5005
R696 vdd.n2645 vdd.n2565 92.5005
R697 vdd.n2648 vdd.n2647 92.5005
R698 vdd.n2647 vdd.n2646 92.5005
R699 vdd.n2564 vdd.n2562 92.5005
R700 vdd.n2622 vdd.n2564 92.5005
R701 vdd.n2611 vdd.n2566 92.5005
R702 vdd.n2607 vdd.n2566 92.5005
R703 vdd.n2610 vdd.n2609 92.5005
R704 vdd.n2609 vdd.n2608 92.5005
R705 vdd.n2598 vdd.n2572 92.5005
R706 vdd.n2606 vdd.n2572 92.5005
R707 vdd.n2583 vdd.n2582 92.5005
R708 vdd.n2582 vdd.n2581 92.5005
R709 vdd.n2604 vdd.n2603 92.5005
R710 vdd.n2605 vdd.n2604 92.5005
R711 vdd.n2620 vdd.n2619 92.5005
R712 vdd.n2621 vdd.n2620 92.5005
R713 vdd.n2674 vdd.n2673 92.5005
R714 vdd.n2675 vdd.n2674 92.5005
R715 vdd.n2669 vdd.n2551 92.5005
R716 vdd.n2676 vdd.n2551 92.5005
R717 vdd.n2680 vdd.n2679 92.5005
R718 vdd.n2679 vdd.n2678 92.5005
R719 vdd.n2682 vdd.n2522 92.5005
R720 vdd.n2534 vdd.n2522 92.5005
R721 vdd.n2533 vdd.n2529 92.5005
R722 vdd.n2534 vdd.n2533 92.5005
R723 vdd.n2536 vdd.n2531 92.5005
R724 vdd.n2536 vdd.n2535 92.5005
R725 vdd.n2539 vdd.n2519 92.5005
R726 vdd.n2535 vdd.n2519 92.5005
R727 vdd.n2708 vdd.n2707 92.5005
R728 vdd.n2705 vdd.n2704 92.5005
R729 vdd.n2722 vdd.n2721 92.5005
R730 vdd.n2721 vdd.n2720 92.5005
R731 vdd.n2719 vdd.n2718 92.5005
R732 vdd.n2720 vdd.n2719 92.5005
R733 vdd.n2525 vdd.n2523 92.5005
R734 vdd.n2523 vdd.n2520 92.5005
R735 vdd.n2794 vdd.n2793 92.5005
R736 vdd.n2793 vdd.n2792 92.5005
R737 vdd.n2773 vdd.n2755 92.5005
R738 vdd.n2809 vdd.n2755 92.5005
R739 vdd.n2759 vdd.n2757 92.5005
R740 vdd.n2757 vdd.n2756 92.5005
R741 vdd.t31 vdd.t2 91.8126
R742 vdd.n2666 vdd.t17 91.4648
R743 vdd.n2666 vdd.t84 91.4648
R744 vdd.n2567 vdd.t86 91.4648
R745 vdd.n700 vdd.n699 86.9025
R746 vdd.n1680 vdd.n77 86.9025
R747 vdd.n2574 vdd.t3 86.7743
R748 vdd.n2631 vdd.t23 86.7743
R749 vdd.n2632 vdd.t9 86.7743
R750 vdd.n2567 vdd.t7 86.7743
R751 vdd.n1931 vdd.n1886 85.9427
R752 vdd.n2481 vdd.n1886 85.9427
R753 vdd.n2854 vdd.n1942 85.9427
R754 vdd.n2882 vdd.n1942 85.9427
R755 vdd.n2902 vdd.n1942 85.9427
R756 vdd.n2942 vdd.n1942 85.9427
R757 vdd.n3007 vdd.n1942 85.9427
R758 vdd.n3032 vdd.n1942 85.9427
R759 vdd.n3029 vdd.n1942 85.9427
R760 vdd.n3059 vdd.n1942 85.9427
R761 vdd.n3080 vdd.n1942 85.9427
R762 vdd.n3108 vdd.n1942 85.9427
R763 vdd.n3128 vdd.n1942 85.9427
R764 vdd.n3168 vdd.n1942 85.9427
R765 vdd.n3233 vdd.n1942 85.9427
R766 vdd.n3258 vdd.n1942 85.9427
R767 vdd.n3255 vdd.n1942 85.9427
R768 vdd.n3285 vdd.n1942 85.9427
R769 vdd.n3306 vdd.n1942 85.9427
R770 vdd.n3334 vdd.n1942 85.9427
R771 vdd.n3354 vdd.n1942 85.9427
R772 vdd.n3394 vdd.n1942 85.9427
R773 vdd.n3459 vdd.n1942 85.9427
R774 vdd.n3484 vdd.n1942 85.9427
R775 vdd.n3481 vdd.n1942 85.9427
R776 vdd.n3511 vdd.n1942 85.9427
R777 vdd.n3532 vdd.n1942 85.9427
R778 vdd.n3560 vdd.n1942 85.9427
R779 vdd.n3580 vdd.n1942 85.9427
R780 vdd.n3620 vdd.n1942 85.9427
R781 vdd.n3685 vdd.n1942 85.9427
R782 vdd vdd.n946 85.8969
R783 vdd vdd.n1197 85.8969
R784 vdd vdd.n1448 85.8969
R785 vdd.n1676 vdd 85.8969
R786 vdd.n2676 vdd.t71 82.8864
R787 vdd vdd.n1840 77.6572
R788 vdd vdd.n2809 77.6572
R789 vdd.n2591 vdd.n2590 76.0005
R790 vdd.n669 vdd.t48 74.7864
R791 vdd.t57 vdd.t31 73.9602
R792 vdd.n1841 vdd 73.4163
R793 vdd.n2608 vdd.t20 71.4099
R794 vdd.n2743 vdd.t80 70.3949
R795 vdd.n649 vdd.t69 70.3649
R796 vdd.n1843 vdd.t52 68.0287
R797 vdd.n2484 vdd.t1 68.0287
R798 vdd.n2574 vdd.t60 68.0124
R799 vdd.n2631 vdd.t77 68.0124
R800 vdd.t94 vdd.n804 67.9081
R801 vdd.t78 vdd.n1055 67.9081
R802 vdd.t42 vdd.n1306 67.9081
R803 vdd.t73 vdd.n1557 67.9081
R804 vdd.n2834 vdd.n2832 67.5405
R805 vdd.n3711 vdd.n3710 67.5405
R806 vdd.n3599 vdd.n2013 67.3307
R807 vdd.n3373 vdd.n2147 67.3307
R808 vdd.n3147 vdd.n2281 67.3307
R809 vdd.n2921 vdd.n2415 67.3307
R810 vdd.n3814 vdd.n3813 67.3307
R811 vdd.n2941 vdd.n2940 67.3307
R812 vdd.n2978 vdd.n2977 67.3307
R813 vdd.n3028 vdd.n3027 67.3307
R814 vdd.n3167 vdd.n3166 67.3307
R815 vdd.n3204 vdd.n3203 67.3307
R816 vdd.n3254 vdd.n3253 67.3307
R817 vdd.n3393 vdd.n3392 67.3307
R818 vdd.n3430 vdd.n3429 67.3307
R819 vdd.n3480 vdd.n3479 67.3307
R820 vdd.n3619 vdd.n3618 67.3307
R821 vdd.n3656 vdd.n3655 67.3307
R822 vdd.n2605 vdd.t18 66.3092
R823 vdd.t68 vdd.t47 65.1272
R824 vdd.n2528 vdd.t25 63.1021
R825 vdd.n670 vdd 58.5621
R826 vdd.n2537 vdd.t15 58.4849
R827 vdd.n2607 vdd.t92 57.383
R828 vdd.t95 vdd.n2677 57.383
R829 vdd.n2606 vdd.t75 53.5575
R830 vdd.n2707 vdd.n2706 52.7184
R831 vdd.n2706 vdd.n2705 52.7178
R832 vdd.n2678 vdd.t95 49.732
R833 vdd.t38 vdd.n2580 48.4569
R834 vdd.t59 vdd.t18 48.4569
R835 vdd.t36 vdd.t6 48.4569
R836 vdd.t55 vdd.t79 47.6077
R837 vdd.t8 vdd.t41 47.1817
R838 vdd.n656 vdd.t44 47.1434
R839 vdd.n656 vdd.t43 47.1434
R840 vdd.n2735 vdd.t33 47.1434
R841 vdd.n2735 vdd.t34 47.1434
R842 vdd.n723 vdd.n595 46.2524
R843 vdd.n725 vdd.n581 46.2524
R844 vdd.n750 vdd.n749 46.2524
R845 vdd.n778 vdd.n777 46.2524
R846 vdd.n802 vdd.n550 46.2524
R847 vdd.n843 vdd.n842 46.2524
R848 vdd.n865 vdd.n864 46.2524
R849 vdd.n886 vdd.n501 46.2524
R850 vdd.n888 vdd.n481 46.2524
R851 vdd.n940 vdd.n939 46.2524
R852 vdd.n974 vdd.n461 46.2524
R853 vdd.n976 vdd.n447 46.2524
R854 vdd.n1001 vdd.n1000 46.2524
R855 vdd.n1029 vdd.n1028 46.2524
R856 vdd.n1053 vdd.n416 46.2524
R857 vdd.n1094 vdd.n1093 46.2524
R858 vdd.n1116 vdd.n1115 46.2524
R859 vdd.n1137 vdd.n367 46.2524
R860 vdd.n1139 vdd.n347 46.2524
R861 vdd.n1191 vdd.n1190 46.2524
R862 vdd.n1225 vdd.n327 46.2524
R863 vdd.n1227 vdd.n313 46.2524
R864 vdd.n1252 vdd.n1251 46.2524
R865 vdd.n1280 vdd.n1279 46.2524
R866 vdd.n1304 vdd.n282 46.2524
R867 vdd.n1345 vdd.n1344 46.2524
R868 vdd.n1367 vdd.n1366 46.2524
R869 vdd.n1388 vdd.n233 46.2524
R870 vdd.n1390 vdd.n213 46.2524
R871 vdd.n1442 vdd.n1441 46.2524
R872 vdd.n1476 vdd.n193 46.2524
R873 vdd.n1478 vdd.n179 46.2524
R874 vdd.n1503 vdd.n1502 46.2524
R875 vdd.n1531 vdd.n1530 46.2524
R876 vdd.n1555 vdd.n148 46.2524
R877 vdd.n1591 vdd.n1590 46.2524
R878 vdd.n1613 vdd.n1612 46.2524
R879 vdd.n1644 vdd.n94 46.2524
R880 vdd.n1646 vdd.n80 46.2524
R881 vdd.n1678 vdd.n1675 46.2524
R882 vdd.n1706 vdd.n1705 46.2524
R883 vdd.n1728 vdd.n1727 46.2524
R884 vdd.n1759 vdd.n30 46.2524
R885 vdd.n1761 vdd.n17 46.2524
R886 vdd.n1849 vdd.n1785 46.2524
R887 vdd.n672 vdd.n667 44.6345
R888 vdd.t22 vdd.t8 44.6314
R889 vdd.t83 vdd.n2676 44.6314
R890 vdd.n947 vdd 41.8475
R891 vdd.n1198 vdd 41.8475
R892 vdd.n1449 vdd 41.8475
R893 vdd.n2579 vdd.t39 41.5552
R894 vdd.n2579 vdd.t19 41.5552
R895 vdd.n1826 vdd.n1825 39.0005
R896 vdd.n2790 vdd.n2757 39.0005
R897 vdd.n2632 vdd.t28 38.6969
R898 vdd vdd.t38 38.2555
R899 vdd.n635 vdd.t48 37.4425
R900 vdd.n2678 vdd 35.7052
R901 vdd.t12 vdd.t24 34.6641
R902 vdd.n944 vdd.n474 33.746
R903 vdd.n1195 vdd.n340 33.746
R904 vdd.n1446 vdd.n206 33.746
R905 vdd.n3031 vdd.n3030 33.746
R906 vdd.n3257 vdd.n3256 33.746
R907 vdd.n3483 vdd.n3482 33.746
R908 vdd.n1828 vdd.n1827 33.6517
R909 vdd.n2791 vdd.n2756 33.6517
R910 vdd.n2608 vdd.t36 33.1549
R911 vdd.t6 vdd.n2607 33.1549
R912 vdd.n816 vdd.n815 32.9702
R913 vdd.n1067 vdd.n1066 32.9702
R914 vdd.n1318 vdd.n1317 32.9702
R915 vdd.n1569 vdd.n1568 32.9702
R916 vdd.n2413 vdd.n2406 32.9702
R917 vdd.n2279 vdd.n2272 32.9702
R918 vdd.n2145 vdd.n2138 32.9702
R919 vdd.n2011 vdd.n2004 32.9702
R920 vdd.n2537 vdd.t50 31.831
R921 vdd.n2490 vdd.n2485 29.4128
R922 vdd.n1844 vdd.n1841 29.2586
R923 vdd.n2612 vdd.t93 28.7575
R924 vdd.n2549 vdd.t5 28.7575
R925 vdd.n805 vdd.t94 28.6326
R926 vdd.t49 vdd.n530 28.6326
R927 vdd.n1056 vdd.t78 28.6326
R928 vdd.t40 vdd.n396 28.6326
R929 vdd.n1307 vdd.t42 28.6326
R930 vdd.t88 vdd.n262 28.6326
R931 vdd.n1558 vdd.t73 28.6326
R932 vdd.t63 vdd.n129 28.6326
R933 vdd.t81 vdd.n65 28.6326
R934 vdd.n1588 vdd.n128 28.2358
R935 vdd.n1611 vdd.n113 28.2358
R936 vdd.n1615 vdd.n95 28.2358
R937 vdd.n1647 vdd.n93 28.2358
R938 vdd.n1673 vdd.n78 28.2358
R939 vdd.n1451 vdd.n207 28.2358
R940 vdd.n1475 vdd.n192 28.2358
R941 vdd.n1500 vdd.n180 28.2358
R942 vdd.n1504 vdd.n163 28.2358
R943 vdd.n1533 vdd.n161 28.2358
R944 vdd.n1554 vdd.n147 28.2358
R945 vdd.n1342 vdd.n261 28.2358
R946 vdd.n1365 vdd.n247 28.2358
R947 vdd.n1369 vdd.n234 28.2358
R948 vdd.n1391 vdd.n232 28.2358
R949 vdd.n1439 vdd.n212 28.2358
R950 vdd.n1447 vdd.n209 28.2358
R951 vdd.n1200 vdd.n341 28.2358
R952 vdd.n1224 vdd.n326 28.2358
R953 vdd.n1249 vdd.n314 28.2358
R954 vdd.n1253 vdd.n297 28.2358
R955 vdd.n1282 vdd.n295 28.2358
R956 vdd.n1303 vdd.n281 28.2358
R957 vdd.n1091 vdd.n395 28.2358
R958 vdd.n1114 vdd.n381 28.2358
R959 vdd.n1118 vdd.n368 28.2358
R960 vdd.n1140 vdd.n366 28.2358
R961 vdd.n1188 vdd.n346 28.2358
R962 vdd.n1196 vdd.n343 28.2358
R963 vdd.n949 vdd.n475 28.2358
R964 vdd.n973 vdd.n460 28.2358
R965 vdd.n998 vdd.n448 28.2358
R966 vdd.n1002 vdd.n431 28.2358
R967 vdd.n1031 vdd.n429 28.2358
R968 vdd.n1052 vdd.n415 28.2358
R969 vdd.n840 vdd.n529 28.2358
R970 vdd.n863 vdd.n515 28.2358
R971 vdd.n867 vdd.n502 28.2358
R972 vdd.n889 vdd.n500 28.2358
R973 vdd.n937 vdd.n480 28.2358
R974 vdd.n945 vdd.n477 28.2358
R975 vdd.n722 vdd.n594 28.2358
R976 vdd.n747 vdd.n582 28.2358
R977 vdd.n751 vdd.n565 28.2358
R978 vdd.n780 vdd.n563 28.2358
R979 vdd.n801 vdd.n549 28.2358
R980 vdd.n1703 vdd.n64 28.2358
R981 vdd.n1726 vdd.n49 28.2358
R982 vdd.n1730 vdd.n31 28.2358
R983 vdd.n1762 vdd.n29 28.2358
R984 vdd.n1783 vdd.n15 28.2358
R985 vdd.n1846 vdd.n16 28.2358
R986 vdd.n3618 vdd.n3617 28.2358
R987 vdd.n3656 vdd.n3654 28.2358
R988 vdd.n3710 vdd.n1943 28.2358
R989 vdd.n3600 vdd.n3599 28.2358
R990 vdd.n3392 vdd.n3391 28.2358
R991 vdd.n3430 vdd.n3428 28.2358
R992 vdd.n3479 vdd.n2078 28.2358
R993 vdd.n3374 vdd.n3373 28.2358
R994 vdd.n3166 vdd.n3165 28.2358
R995 vdd.n3204 vdd.n3202 28.2358
R996 vdd.n3253 vdd.n2212 28.2358
R997 vdd.n3148 vdd.n3147 28.2358
R998 vdd.n2940 vdd.n2939 28.2358
R999 vdd.n2978 vdd.n2976 28.2358
R1000 vdd.n3027 vdd.n2346 28.2358
R1001 vdd.n2834 vdd.n2833 28.2358
R1002 vdd.n2922 vdd.n2921 28.2358
R1003 vdd.n3756 vdd.n1920 28.2358
R1004 vdd.n3775 vdd.n1909 28.2358
R1005 vdd.n3794 vdd.n1898 28.2358
R1006 vdd.n3813 vdd.n1887 28.2358
R1007 vdd.n2528 vdd.t13 28.0332
R1008 vdd.n2775 vdd.n2774 27.3454
R1009 vdd.n670 vdd.n667 27.1882
R1010 vdd.t91 vdd.n2606 26.779
R1011 vdd.t20 vdd.t91 26.779
R1012 vdd.t92 vdd 25.5039
R1013 vdd vdd.t4 25.5039
R1014 vdd.t16 vdd.n2675 24.2287
R1015 vdd.n696 vdd.n695 23.4935
R1016 vdd.n2789 vdd.n2788 22.8875
R1017 vdd.t79 vdd.t32 21.1252
R1018 vdd.n622 vdd.n609 20.7428
R1019 vdd.n635 vdd.n634 20.7428
R1020 vdd.n637 vdd.n635 20.7428
R1021 vdd.n644 vdd.n609 20.7428
R1022 vdd.n695 vdd.n694 20.7428
R1023 vdd.n2493 vdd.n2491 20.7428
R1024 vdd.n2489 vdd.n2488 20.7428
R1025 vdd.n2507 vdd.n2506 20.7428
R1026 vdd.n2815 vdd.n2813 20.7428
R1027 vdd.n2811 vdd.n2753 20.7428
R1028 vdd.n804 vdd.t49 20.3031
R1029 vdd.n1055 vdd.t40 20.3031
R1030 vdd.n1306 vdd.t88 20.3031
R1031 vdd.n1557 vdd.t63 20.3031
R1032 vdd.n2706 vdd.n2521 19.8929
R1033 vdd vdd.t51 19.8228
R1034 vdd.n2581 vdd 19.128
R1035 vdd vdd.t85 19.128
R1036 vdd.n2489 vdd.t87 18.5229
R1037 vdd.t29 vdd.t12 17.3323
R1038 vdd.t41 vdd.n2644 16.5777
R1039 vdd vdd.t61 16.5329
R1040 vdd.t10 vdd.n2507 16.3798
R1041 vdd.n1792 vdd.n1791 15.4666
R1042 vdd.n2796 vdd.n2795 15.4666
R1043 vdd.n2623 vdd.t26 15.3025
R1044 vdd vdd.n1786 15.1421
R1045 vdd.n2772 vdd 15.1421
R1046 vdd.t74 vdd.n2623 14.0273
R1047 vdd.n1844 vdd.n1843 13.6721
R1048 vdd.n2485 vdd.n2484 13.3673
R1049 vdd.n3621 vdd.n3620 13.1177
R1050 vdd.n3685 vdd.n3684 13.1177
R1051 vdd.n3511 vdd.n2050 13.1177
R1052 vdd.n3532 vdd.n2035 13.1177
R1053 vdd.n3561 vdd.n3560 13.1177
R1054 vdd.n3581 vdd.n3580 13.1177
R1055 vdd.n3395 vdd.n3394 13.1177
R1056 vdd.n3459 vdd.n3458 13.1177
R1057 vdd.n3485 vdd.n3484 13.1177
R1058 vdd.n3285 vdd.n2184 13.1177
R1059 vdd.n3306 vdd.n2169 13.1177
R1060 vdd.n3335 vdd.n3334 13.1177
R1061 vdd.n3355 vdd.n3354 13.1177
R1062 vdd.n3169 vdd.n3168 13.1177
R1063 vdd.n3233 vdd.n3232 13.1177
R1064 vdd.n3259 vdd.n3258 13.1177
R1065 vdd.n3059 vdd.n2318 13.1177
R1066 vdd.n3080 vdd.n2303 13.1177
R1067 vdd.n3109 vdd.n3108 13.1177
R1068 vdd.n3129 vdd.n3128 13.1177
R1069 vdd.n2943 vdd.n2942 13.1177
R1070 vdd.n3007 vdd.n3006 13.1177
R1071 vdd.n3033 vdd.n3032 13.1177
R1072 vdd.n2854 vdd.n2437 13.1177
R1073 vdd.n2883 vdd.n2882 13.1177
R1074 vdd.n2903 vdd.n2902 13.1177
R1075 vdd.n3737 vdd.n1931 13.1177
R1076 vdd.n2481 vdd.n1885 13.1177
R1077 vdd.n3719 vdd.n1931 13.1177
R1078 vdd.n2942 vdd.n2376 13.1177
R1079 vdd.n3008 vdd.n3007 13.1177
R1080 vdd.n3168 vdd.n2242 13.1177
R1081 vdd.n3234 vdd.n3233 13.1177
R1082 vdd.n3394 vdd.n2108 13.1177
R1083 vdd.n3460 vdd.n3459 13.1177
R1084 vdd.n3620 vdd.n1974 13.1177
R1085 vdd.n3686 vdd.n3685 13.1177
R1086 vdd.n3580 vdd.n3579 13.1177
R1087 vdd.n3560 vdd.n3559 13.1177
R1088 vdd.n3533 vdd.n3532 13.1177
R1089 vdd.n3512 vdd.n3511 13.1177
R1090 vdd.n3481 vdd.n2061 13.1177
R1091 vdd.n3354 vdd.n3353 13.1177
R1092 vdd.n3334 vdd.n3333 13.1177
R1093 vdd.n3307 vdd.n3306 13.1177
R1094 vdd.n3286 vdd.n3285 13.1177
R1095 vdd.n3255 vdd.n2195 13.1177
R1096 vdd.n3128 vdd.n3127 13.1177
R1097 vdd.n3108 vdd.n3107 13.1177
R1098 vdd.n3081 vdd.n3080 13.1177
R1099 vdd.n3060 vdd.n3059 13.1177
R1100 vdd.n3029 vdd.n2329 13.1177
R1101 vdd.n2902 vdd.n2901 13.1177
R1102 vdd.n2882 vdd.n2881 13.1177
R1103 vdd.n2855 vdd.n2854 13.1177
R1104 vdd.n79 vdd.n77 13.0163
R1105 vdd.n699 vdd.n608 13.0163
R1106 vdd.n673 vdd.n664 12.5282
R1107 vdd.n1847 vdd.n1841 12.4812
R1108 vdd.t70 vdd.n2812 12.2467
R1109 vdd.n1830 vdd.n1826 12.0005
R1110 vdd.n2807 vdd.n2757 12.0005
R1111 vdd.n2794 vdd.n2788 11.9758
R1112 vdd.n698 vdd.n697 11.747
R1113 vdd.n724 vdd.n723 11.747
R1114 vdd.n748 vdd.n581 11.747
R1115 vdd.n750 vdd.n564 11.747
R1116 vdd.n779 vdd.n778 11.747
R1117 vdd.n803 vdd.n802 11.747
R1118 vdd.n842 vdd.n841 11.747
R1119 vdd.n864 vdd.n514 11.747
R1120 vdd.n866 vdd.n501 11.747
R1121 vdd.n888 vdd.n887 11.747
R1122 vdd.n939 vdd.n938 11.747
R1123 vdd.n946 vdd.n476 11.747
R1124 vdd.n948 vdd.n947 11.747
R1125 vdd.n975 vdd.n974 11.747
R1126 vdd.n999 vdd.n447 11.747
R1127 vdd.n1001 vdd.n430 11.747
R1128 vdd.n1030 vdd.n1029 11.747
R1129 vdd.n1054 vdd.n1053 11.747
R1130 vdd.n1093 vdd.n1092 11.747
R1131 vdd.n1115 vdd.n380 11.747
R1132 vdd.n1117 vdd.n367 11.747
R1133 vdd.n1139 vdd.n1138 11.747
R1134 vdd.n1190 vdd.n1189 11.747
R1135 vdd.n1197 vdd.n342 11.747
R1136 vdd.n1199 vdd.n1198 11.747
R1137 vdd.n1226 vdd.n1225 11.747
R1138 vdd.n1250 vdd.n313 11.747
R1139 vdd.n1252 vdd.n296 11.747
R1140 vdd.n1281 vdd.n1280 11.747
R1141 vdd.n1305 vdd.n1304 11.747
R1142 vdd.n1344 vdd.n1343 11.747
R1143 vdd.n1366 vdd.n246 11.747
R1144 vdd.n1368 vdd.n233 11.747
R1145 vdd.n1390 vdd.n1389 11.747
R1146 vdd.n1441 vdd.n1440 11.747
R1147 vdd.n1448 vdd.n208 11.747
R1148 vdd.n1450 vdd.n1449 11.747
R1149 vdd.n1477 vdd.n1476 11.747
R1150 vdd.n1501 vdd.n179 11.747
R1151 vdd.n1503 vdd.n162 11.747
R1152 vdd.n1532 vdd.n1531 11.747
R1153 vdd.n1556 vdd.n1555 11.747
R1154 vdd.n1590 vdd.n1589 11.747
R1155 vdd.n1612 vdd.n112 11.747
R1156 vdd.n1614 vdd.n94 11.747
R1157 vdd.n1646 vdd.n1645 11.747
R1158 vdd.n1675 vdd.n1674 11.747
R1159 vdd.n1677 vdd.n1676 11.747
R1160 vdd.n1705 vdd.n1704 11.747
R1161 vdd.n1727 vdd.n48 11.747
R1162 vdd.n1729 vdd.n30 11.747
R1163 vdd.n1761 vdd.n1760 11.747
R1164 vdd.n1785 vdd.n1784 11.747
R1165 vdd.n1848 vdd.n1847 11.747
R1166 vdd.n3712 vdd.n3711 11.5452
R1167 vdd.n2832 vdd.n2831 11.5452
R1168 vdd.n2813 vdd.t70 11.4813
R1169 vdd.t4 vdd.t83 11.477
R1170 vdd.n1838 vdd.n1837 11.2229
R1171 vdd.n2774 vdd.n2773 11.2229
R1172 vdd.n1829 vdd.n1828 10.3547
R1173 vdd.n2808 vdd.n2756 10.3547
R1174 vdd.n2580 vdd.t59 10.2018
R1175 vdd.n2645 vdd.t22 10.2018
R1176 vdd.t71 vdd.t16 10.2018
R1177 vdd.n2813 vdd.t10 9.64439
R1178 vdd.n3616 vdd.n3615 9.38471
R1179 vdd.n3602 vdd.n3601 9.38471
R1180 vdd.n3390 vdd.n3389 9.38471
R1181 vdd.n3376 vdd.n3375 9.38471
R1182 vdd.n3164 vdd.n3163 9.38471
R1183 vdd.n3150 vdd.n3149 9.38471
R1184 vdd.n2938 vdd.n2937 9.38471
R1185 vdd.n2924 vdd.n2923 9.38471
R1186 vdd.n815 vdd.n814 9.3005
R1187 vdd.n816 vdd.n541 9.3005
R1188 vdd.n934 vdd.n933 9.3005
R1189 vdd.n1066 vdd.n1065 9.3005
R1190 vdd.n1067 vdd.n407 9.3005
R1191 vdd.n1185 vdd.n1184 9.3005
R1192 vdd.n1317 vdd.n1316 9.3005
R1193 vdd.n1318 vdd.n273 9.3005
R1194 vdd.n1436 vdd.n1435 9.3005
R1195 vdd.n1568 vdd.n1567 9.3005
R1196 vdd.n1569 vdd.n139 9.3005
R1197 vdd.n1670 vdd.n1669 9.3005
R1198 vdd.n1649 vdd.n91 9.3005
R1199 vdd.n1619 vdd.n1618 9.3005
R1200 vdd.n1609 vdd.n1608 9.3005
R1201 vdd.n1585 vdd.n1584 9.3005
R1202 vdd.n1552 vdd.n1551 9.3005
R1203 vdd.n169 vdd.n168 9.3005
R1204 vdd.n1507 vdd.n1506 9.3005
R1205 vdd.n1483 vdd.n1482 9.3005
R1206 vdd.n1473 vdd.n1472 9.3005
R1207 vdd.n1395 vdd.n1394 9.3005
R1208 vdd.n1373 vdd.n1372 9.3005
R1209 vdd.n1363 vdd.n1362 9.3005
R1210 vdd.n1339 vdd.n1338 9.3005
R1211 vdd.n1301 vdd.n1300 9.3005
R1212 vdd.n303 vdd.n302 9.3005
R1213 vdd.n1256 vdd.n1255 9.3005
R1214 vdd.n1232 vdd.n1231 9.3005
R1215 vdd.n1222 vdd.n1221 9.3005
R1216 vdd.n1144 vdd.n1143 9.3005
R1217 vdd.n1122 vdd.n1121 9.3005
R1218 vdd.n1112 vdd.n1111 9.3005
R1219 vdd.n1088 vdd.n1087 9.3005
R1220 vdd.n1050 vdd.n1049 9.3005
R1221 vdd.n437 vdd.n436 9.3005
R1222 vdd.n1005 vdd.n1004 9.3005
R1223 vdd.n981 vdd.n980 9.3005
R1224 vdd.n971 vdd.n970 9.3005
R1225 vdd.n893 vdd.n892 9.3005
R1226 vdd.n871 vdd.n870 9.3005
R1227 vdd.n861 vdd.n860 9.3005
R1228 vdd.n837 vdd.n836 9.3005
R1229 vdd.n799 vdd.n798 9.3005
R1230 vdd.n571 vdd.n570 9.3005
R1231 vdd.n730 vdd.n729 9.3005
R1232 vdd.n754 vdd.n753 9.3005
R1233 vdd.n720 vdd.n719 9.3005
R1234 vdd.n1780 vdd.n1779 9.3005
R1235 vdd.n1764 vdd.n27 9.3005
R1236 vdd.n1734 vdd.n1733 9.3005
R1237 vdd.n1700 vdd.n1699 9.3005
R1238 vdd.n1724 vdd.n1723 9.3005
R1239 vdd.n1767 vdd.n19 9.3005
R1240 vdd.n19 vdd.n18 9.3005
R1241 vdd.n18 vdd.n17 9.3005
R1242 vdd.n1757 vdd.n1756 9.3005
R1243 vdd.n1758 vdd.n1757 9.3005
R1244 vdd.n1759 vdd.n1758 9.3005
R1245 vdd.n1709 vdd.n1708 9.3005
R1246 vdd.n1708 vdd.n1707 9.3005
R1247 vdd.n1707 vdd.n1706 9.3005
R1248 vdd.n46 vdd.n45 9.3005
R1249 vdd.n47 vdd.n46 9.3005
R1250 vdd.n1728 vdd.n47 9.3005
R1251 vdd.n1852 vdd.n1851 9.3005
R1252 vdd.n1851 vdd.n1850 9.3005
R1253 vdd.n1850 vdd.n1849 9.3005
R1254 vdd.n67 vdd.n66 9.3005
R1255 vdd.n66 vdd.n65 9.3005
R1256 vdd.n1652 vdd.n82 9.3005
R1257 vdd.n82 vdd.n81 9.3005
R1258 vdd.n81 vdd.n80 9.3005
R1259 vdd.n1642 vdd.n1641 9.3005
R1260 vdd.n1643 vdd.n1642 9.3005
R1261 vdd.n1644 vdd.n1643 9.3005
R1262 vdd.n110 vdd.n109 9.3005
R1263 vdd.n111 vdd.n110 9.3005
R1264 vdd.n1613 vdd.n111 9.3005
R1265 vdd.n1594 vdd.n1593 9.3005
R1266 vdd.n1593 vdd.n1592 9.3005
R1267 vdd.n1592 vdd.n1591 9.3005
R1268 vdd.n1681 vdd.n1680 9.3005
R1269 vdd.n1680 vdd.n1679 9.3005
R1270 vdd.n1679 vdd.n1678 9.3005
R1271 vdd.n1572 vdd.n131 9.3005
R1272 vdd.n131 vdd.n130 9.3005
R1273 vdd.n130 vdd.n129 9.3005
R1274 vdd.n1536 vdd.n1535 9.3005
R1275 vdd.n1535 vdd.n149 9.3005
R1276 vdd.n149 vdd.n148 9.3005
R1277 vdd.n1528 vdd.n1527 9.3005
R1278 vdd.n1529 vdd.n1528 9.3005
R1279 vdd.n1530 vdd.n1529 9.3005
R1280 vdd.n1498 vdd.n1497 9.3005
R1281 vdd.n1498 vdd.n178 9.3005
R1282 vdd.n1502 vdd.n178 9.3005
R1283 vdd.n1480 vdd.n191 9.3005
R1284 vdd.n1480 vdd.n1479 9.3005
R1285 vdd.n1479 vdd.n1478 9.3005
R1286 vdd.n1561 vdd.n1560 9.3005
R1287 vdd.n1560 vdd.n1559 9.3005
R1288 vdd.n1559 vdd.n1558 9.3005
R1289 vdd.n1454 vdd.n1453 9.3005
R1290 vdd.n1453 vdd.n194 9.3005
R1291 vdd.n194 vdd.n193 9.3005
R1292 vdd.n1407 vdd.n215 9.3005
R1293 vdd.n215 vdd.n214 9.3005
R1294 vdd.n214 vdd.n213 9.3005
R1295 vdd.n1386 vdd.n1385 9.3005
R1296 vdd.n1387 vdd.n1386 9.3005
R1297 vdd.n1388 vdd.n1387 9.3005
R1298 vdd.n251 vdd.n244 9.3005
R1299 vdd.n245 vdd.n244 9.3005
R1300 vdd.n1367 vdd.n245 9.3005
R1301 vdd.n1348 vdd.n1347 9.3005
R1302 vdd.n1347 vdd.n1346 9.3005
R1303 vdd.n1346 vdd.n1345 9.3005
R1304 vdd.n1444 vdd.n211 9.3005
R1305 vdd.n1444 vdd.n1443 9.3005
R1306 vdd.n1443 vdd.n1442 9.3005
R1307 vdd.n1321 vdd.n264 9.3005
R1308 vdd.n264 vdd.n263 9.3005
R1309 vdd.n263 vdd.n262 9.3005
R1310 vdd.n1285 vdd.n1284 9.3005
R1311 vdd.n1284 vdd.n283 9.3005
R1312 vdd.n283 vdd.n282 9.3005
R1313 vdd.n1277 vdd.n1276 9.3005
R1314 vdd.n1278 vdd.n1277 9.3005
R1315 vdd.n1279 vdd.n1278 9.3005
R1316 vdd.n1247 vdd.n1246 9.3005
R1317 vdd.n1247 vdd.n312 9.3005
R1318 vdd.n1251 vdd.n312 9.3005
R1319 vdd.n1229 vdd.n325 9.3005
R1320 vdd.n1229 vdd.n1228 9.3005
R1321 vdd.n1228 vdd.n1227 9.3005
R1322 vdd.n1310 vdd.n1309 9.3005
R1323 vdd.n1309 vdd.n1308 9.3005
R1324 vdd.n1308 vdd.n1307 9.3005
R1325 vdd.n1203 vdd.n1202 9.3005
R1326 vdd.n1202 vdd.n328 9.3005
R1327 vdd.n328 vdd.n327 9.3005
R1328 vdd.n1156 vdd.n349 9.3005
R1329 vdd.n349 vdd.n348 9.3005
R1330 vdd.n348 vdd.n347 9.3005
R1331 vdd.n1135 vdd.n1134 9.3005
R1332 vdd.n1136 vdd.n1135 9.3005
R1333 vdd.n1137 vdd.n1136 9.3005
R1334 vdd.n385 vdd.n378 9.3005
R1335 vdd.n379 vdd.n378 9.3005
R1336 vdd.n1116 vdd.n379 9.3005
R1337 vdd.n1097 vdd.n1096 9.3005
R1338 vdd.n1096 vdd.n1095 9.3005
R1339 vdd.n1095 vdd.n1094 9.3005
R1340 vdd.n1193 vdd.n345 9.3005
R1341 vdd.n1193 vdd.n1192 9.3005
R1342 vdd.n1192 vdd.n1191 9.3005
R1343 vdd.n1070 vdd.n398 9.3005
R1344 vdd.n398 vdd.n397 9.3005
R1345 vdd.n397 vdd.n396 9.3005
R1346 vdd.n1034 vdd.n1033 9.3005
R1347 vdd.n1033 vdd.n417 9.3005
R1348 vdd.n417 vdd.n416 9.3005
R1349 vdd.n1026 vdd.n1025 9.3005
R1350 vdd.n1027 vdd.n1026 9.3005
R1351 vdd.n1028 vdd.n1027 9.3005
R1352 vdd.n996 vdd.n995 9.3005
R1353 vdd.n996 vdd.n446 9.3005
R1354 vdd.n1000 vdd.n446 9.3005
R1355 vdd.n978 vdd.n459 9.3005
R1356 vdd.n978 vdd.n977 9.3005
R1357 vdd.n977 vdd.n976 9.3005
R1358 vdd.n1059 vdd.n1058 9.3005
R1359 vdd.n1058 vdd.n1057 9.3005
R1360 vdd.n1057 vdd.n1056 9.3005
R1361 vdd.n952 vdd.n951 9.3005
R1362 vdd.n951 vdd.n462 9.3005
R1363 vdd.n462 vdd.n461 9.3005
R1364 vdd.n905 vdd.n483 9.3005
R1365 vdd.n483 vdd.n482 9.3005
R1366 vdd.n482 vdd.n481 9.3005
R1367 vdd.n884 vdd.n883 9.3005
R1368 vdd.n885 vdd.n884 9.3005
R1369 vdd.n886 vdd.n885 9.3005
R1370 vdd.n519 vdd.n512 9.3005
R1371 vdd.n513 vdd.n512 9.3005
R1372 vdd.n865 vdd.n513 9.3005
R1373 vdd.n846 vdd.n845 9.3005
R1374 vdd.n845 vdd.n844 9.3005
R1375 vdd.n844 vdd.n843 9.3005
R1376 vdd.n942 vdd.n479 9.3005
R1377 vdd.n942 vdd.n941 9.3005
R1378 vdd.n941 vdd.n940 9.3005
R1379 vdd.n819 vdd.n532 9.3005
R1380 vdd.n532 vdd.n531 9.3005
R1381 vdd.n531 vdd.n530 9.3005
R1382 vdd.n783 vdd.n782 9.3005
R1383 vdd.n782 vdd.n551 9.3005
R1384 vdd.n551 vdd.n550 9.3005
R1385 vdd.n775 vdd.n774 9.3005
R1386 vdd.n776 vdd.n775 9.3005
R1387 vdd.n777 vdd.n776 9.3005
R1388 vdd.n727 vdd.n593 9.3005
R1389 vdd.n727 vdd.n726 9.3005
R1390 vdd.n726 vdd.n725 9.3005
R1391 vdd.n745 vdd.n744 9.3005
R1392 vdd.n745 vdd.n580 9.3005
R1393 vdd.n749 vdd.n580 9.3005
R1394 vdd.n808 vdd.n807 9.3005
R1395 vdd.n807 vdd.n806 9.3005
R1396 vdd.n806 vdd.n805 9.3005
R1397 vdd.n701 vdd.n700 9.3005
R1398 vdd.n700 vdd.n596 9.3005
R1399 vdd.n596 vdd.n595 9.3005
R1400 vdd.n1831 vdd.n1830 9.3005
R1401 vdd.n1830 vdd.n1829 9.3005
R1402 vdd.n2413 vdd.n2412 9.3005
R1403 vdd.n3025 vdd.n3024 9.3005
R1404 vdd.n2981 vdd.n2980 9.3005
R1405 vdd.n2948 vdd.n2947 9.3005
R1406 vdd.n2407 vdd.n2406 9.3005
R1407 vdd.n2378 vdd.n2377 9.3005
R1408 vdd.n2363 vdd.n2362 9.3005
R1409 vdd.n2279 vdd.n2278 9.3005
R1410 vdd.n3251 vdd.n3250 9.3005
R1411 vdd.n3207 vdd.n3206 9.3005
R1412 vdd.n3174 vdd.n3173 9.3005
R1413 vdd.n2273 vdd.n2272 9.3005
R1414 vdd.n2244 vdd.n2243 9.3005
R1415 vdd.n2229 vdd.n2228 9.3005
R1416 vdd.n2145 vdd.n2144 9.3005
R1417 vdd.n3477 vdd.n3476 9.3005
R1418 vdd.n3433 vdd.n3432 9.3005
R1419 vdd.n3400 vdd.n3399 9.3005
R1420 vdd.n2139 vdd.n2138 9.3005
R1421 vdd.n2110 vdd.n2109 9.3005
R1422 vdd.n2095 vdd.n2094 9.3005
R1423 vdd.n2011 vdd.n2010 9.3005
R1424 vdd.n3708 vdd.n3707 9.3005
R1425 vdd.n3659 vdd.n3658 9.3005
R1426 vdd.n3626 vdd.n3625 9.3005
R1427 vdd.n2005 vdd.n2004 9.3005
R1428 vdd.n1976 vdd.n1975 9.3005
R1429 vdd.n1961 vdd.n1960 9.3005
R1430 vdd.n3597 vdd.n3596 9.3005
R1431 vdd.n3577 vdd.n3576 9.3005
R1432 vdd.n2041 vdd.n2040 9.3005
R1433 vdd.n3536 vdd.n3535 9.3005
R1434 vdd.n3515 vdd.n3514 9.3005
R1435 vdd.n3371 vdd.n3370 9.3005
R1436 vdd.n3351 vdd.n3350 9.3005
R1437 vdd.n2175 vdd.n2174 9.3005
R1438 vdd.n3310 vdd.n3309 9.3005
R1439 vdd.n3289 vdd.n3288 9.3005
R1440 vdd.n3145 vdd.n3144 9.3005
R1441 vdd.n3125 vdd.n3124 9.3005
R1442 vdd.n2309 vdd.n2308 9.3005
R1443 vdd.n3084 vdd.n3083 9.3005
R1444 vdd.n3063 vdd.n3062 9.3005
R1445 vdd.n2919 vdd.n2918 9.3005
R1446 vdd.n2899 vdd.n2898 9.3005
R1447 vdd.n2443 vdd.n2442 9.3005
R1448 vdd.n2837 vdd.n2836 9.3005
R1449 vdd.n2858 vdd.n2857 9.3005
R1450 vdd.n3735 vdd.n3734 9.3005
R1451 vdd.n3754 vdd.n3753 9.3005
R1452 vdd.n3773 vdd.n3772 9.3005
R1453 vdd.n3792 vdd.n3791 9.3005
R1454 vdd.n3811 vdd.n3810 9.3005
R1455 vdd.n3741 vdd.n3740 9.3005
R1456 vdd.n3740 vdd.n3739 9.3005
R1457 vdd.n3760 vdd.n3759 9.3005
R1458 vdd.n3759 vdd.n3758 9.3005
R1459 vdd.n3779 vdd.n3778 9.3005
R1460 vdd.n3778 vdd.n3777 9.3005
R1461 vdd.n3798 vdd.n3797 9.3005
R1462 vdd.n3797 vdd.n3796 9.3005
R1463 vdd.n3817 vdd.n3816 9.3005
R1464 vdd.n3816 vdd.n3815 9.3005
R1465 vdd.n3721 vdd.n3720 9.3005
R1466 vdd.n3720 vdd.n1886 9.3005
R1467 vdd.n3036 vdd.n3035 9.3005
R1468 vdd.n3035 vdd.n3034 9.3005
R1469 vdd.n3004 vdd.n3003 9.3005
R1470 vdd.n3004 vdd.n2358 9.3005
R1471 vdd.n2945 vdd.n2380 9.3005
R1472 vdd.n2945 vdd.n2944 9.3005
R1473 vdd.n2937 vdd.n2936 9.3005
R1474 vdd.n2973 vdd.n2374 9.3005
R1475 vdd.n2974 vdd.n2973 9.3005
R1476 vdd.n3012 vdd.n3011 9.3005
R1477 vdd.n3011 vdd.n3010 9.3005
R1478 vdd.n3262 vdd.n3261 9.3005
R1479 vdd.n3261 vdd.n3260 9.3005
R1480 vdd.n3230 vdd.n3229 9.3005
R1481 vdd.n3230 vdd.n2224 9.3005
R1482 vdd.n3171 vdd.n2246 9.3005
R1483 vdd.n3171 vdd.n3170 9.3005
R1484 vdd.n3163 vdd.n3162 9.3005
R1485 vdd.n3199 vdd.n2240 9.3005
R1486 vdd.n3200 vdd.n3199 9.3005
R1487 vdd.n3238 vdd.n3237 9.3005
R1488 vdd.n3237 vdd.n3236 9.3005
R1489 vdd.n3488 vdd.n3487 9.3005
R1490 vdd.n3487 vdd.n3486 9.3005
R1491 vdd.n3456 vdd.n3455 9.3005
R1492 vdd.n3456 vdd.n2090 9.3005
R1493 vdd.n3397 vdd.n2112 9.3005
R1494 vdd.n3397 vdd.n3396 9.3005
R1495 vdd.n3389 vdd.n3388 9.3005
R1496 vdd.n3425 vdd.n2106 9.3005
R1497 vdd.n3426 vdd.n3425 9.3005
R1498 vdd.n3464 vdd.n3463 9.3005
R1499 vdd.n3463 vdd.n3462 9.3005
R1500 vdd.n3682 vdd.n3681 9.3005
R1501 vdd.n3682 vdd.n1956 9.3005
R1502 vdd.n3623 vdd.n1978 9.3005
R1503 vdd.n3623 vdd.n3622 9.3005
R1504 vdd.n3615 vdd.n3614 9.3005
R1505 vdd.n3651 vdd.n1972 9.3005
R1506 vdd.n3652 vdd.n3651 9.3005
R1507 vdd.n3690 vdd.n3689 9.3005
R1508 vdd.n3689 vdd.n3688 9.3005
R1509 vdd.n3713 vdd.n3712 9.3005
R1510 vdd.n3584 vdd.n3583 9.3005
R1511 vdd.n3583 vdd.n3582 9.3005
R1512 vdd.n3564 vdd.n3563 9.3005
R1513 vdd.n3563 vdd.n2024 9.3005
R1514 vdd.n2024 vdd.n1942 9.3005
R1515 vdd.n3557 vdd.n3556 9.3005
R1516 vdd.n3558 vdd.n3557 9.3005
R1517 vdd.n3558 vdd.n1942 9.3005
R1518 vdd.n3530 vdd.n3529 9.3005
R1519 vdd.n3531 vdd.n3530 9.3005
R1520 vdd.n3531 vdd.n1942 9.3005
R1521 vdd.n3603 vdd.n3602 9.3005
R1522 vdd.n3509 vdd.n3508 9.3005
R1523 vdd.n3510 vdd.n3509 9.3005
R1524 vdd.n3510 vdd.n1942 9.3005
R1525 vdd.n3358 vdd.n3357 9.3005
R1526 vdd.n3357 vdd.n3356 9.3005
R1527 vdd.n3338 vdd.n3337 9.3005
R1528 vdd.n3337 vdd.n2158 9.3005
R1529 vdd.n2158 vdd.n1942 9.3005
R1530 vdd.n3331 vdd.n3330 9.3005
R1531 vdd.n3332 vdd.n3331 9.3005
R1532 vdd.n3332 vdd.n1942 9.3005
R1533 vdd.n3304 vdd.n3303 9.3005
R1534 vdd.n3305 vdd.n3304 9.3005
R1535 vdd.n3305 vdd.n1942 9.3005
R1536 vdd.n3377 vdd.n3376 9.3005
R1537 vdd.n3283 vdd.n3282 9.3005
R1538 vdd.n3284 vdd.n3283 9.3005
R1539 vdd.n3284 vdd.n1942 9.3005
R1540 vdd.n3132 vdd.n3131 9.3005
R1541 vdd.n3131 vdd.n3130 9.3005
R1542 vdd.n3112 vdd.n3111 9.3005
R1543 vdd.n3111 vdd.n2292 9.3005
R1544 vdd.n2292 vdd.n1942 9.3005
R1545 vdd.n3105 vdd.n3104 9.3005
R1546 vdd.n3106 vdd.n3105 9.3005
R1547 vdd.n3106 vdd.n1942 9.3005
R1548 vdd.n3078 vdd.n3077 9.3005
R1549 vdd.n3079 vdd.n3078 9.3005
R1550 vdd.n3079 vdd.n1942 9.3005
R1551 vdd.n3151 vdd.n3150 9.3005
R1552 vdd.n3057 vdd.n3056 9.3005
R1553 vdd.n3058 vdd.n3057 9.3005
R1554 vdd.n3058 vdd.n1942 9.3005
R1555 vdd.n2906 vdd.n2905 9.3005
R1556 vdd.n2905 vdd.n2904 9.3005
R1557 vdd.n2886 vdd.n2885 9.3005
R1558 vdd.n2885 vdd.n2426 9.3005
R1559 vdd.n2426 vdd.n1942 9.3005
R1560 vdd.n2879 vdd.n2878 9.3005
R1561 vdd.n2880 vdd.n2879 9.3005
R1562 vdd.n2880 vdd.n1942 9.3005
R1563 vdd.n2925 vdd.n2924 9.3005
R1564 vdd.n2831 vdd.n2830 9.3005
R1565 vdd.n2852 vdd.n2851 9.3005
R1566 vdd.n2853 vdd.n2852 9.3005
R1567 vdd.n2776 vdd.n2775 9.3005
R1568 vdd.n2806 vdd.n2805 9.3005
R1569 vdd.n2807 vdd.n2806 9.3005
R1570 vdd.n2808 vdd.n2807 9.3005
R1571 vdd.n2700 vdd.n2532 8.98981
R1572 vdd.n2723 vdd.n2517 8.98981
R1573 vdd.t82 vdd.n2622 8.92668
R1574 vdd.n721 vdd.n720 8.92171
R1575 vdd.n729 vdd.n583 8.92171
R1576 vdd.n753 vdd.n752 8.92171
R1577 vdd.n570 vdd.n562 8.92171
R1578 vdd.n800 vdd.n799 8.92171
R1579 vdd.n838 vdd.n837 8.92171
R1580 vdd.n862 vdd.n861 8.92171
R1581 vdd.n870 vdd.n869 8.92171
R1582 vdd.n892 vdd.n890 8.92171
R1583 vdd.n935 vdd.n934 8.92171
R1584 vdd.n972 vdd.n971 8.92171
R1585 vdd.n980 vdd.n449 8.92171
R1586 vdd.n1004 vdd.n1003 8.92171
R1587 vdd.n436 vdd.n428 8.92171
R1588 vdd.n1051 vdd.n1050 8.92171
R1589 vdd.n1089 vdd.n1088 8.92171
R1590 vdd.n1113 vdd.n1112 8.92171
R1591 vdd.n1121 vdd.n1120 8.92171
R1592 vdd.n1143 vdd.n1141 8.92171
R1593 vdd.n1186 vdd.n1185 8.92171
R1594 vdd.n1223 vdd.n1222 8.92171
R1595 vdd.n1231 vdd.n315 8.92171
R1596 vdd.n1255 vdd.n1254 8.92171
R1597 vdd.n302 vdd.n294 8.92171
R1598 vdd.n1302 vdd.n1301 8.92171
R1599 vdd.n1340 vdd.n1339 8.92171
R1600 vdd.n1364 vdd.n1363 8.92171
R1601 vdd.n1372 vdd.n1371 8.92171
R1602 vdd.n1394 vdd.n1392 8.92171
R1603 vdd.n1437 vdd.n1436 8.92171
R1604 vdd.n1474 vdd.n1473 8.92171
R1605 vdd.n1482 vdd.n181 8.92171
R1606 vdd.n1506 vdd.n1505 8.92171
R1607 vdd.n168 vdd.n160 8.92171
R1608 vdd.n1553 vdd.n1552 8.92171
R1609 vdd.n1586 vdd.n1585 8.92171
R1610 vdd.n1610 vdd.n1609 8.92171
R1611 vdd.n1618 vdd.n1617 8.92171
R1612 vdd.n1649 vdd.n1648 8.92171
R1613 vdd.n1671 vdd.n1670 8.92171
R1614 vdd.n1701 vdd.n1700 8.92171
R1615 vdd.n1725 vdd.n1724 8.92171
R1616 vdd.n1733 vdd.n1732 8.92171
R1617 vdd.n1764 vdd.n1763 8.92171
R1618 vdd.n1781 vdd.n1780 8.92171
R1619 vdd.n2836 vdd.n2835 8.92171
R1620 vdd.n2857 vdd.n2856 8.92171
R1621 vdd.n2442 vdd.n2436 8.92171
R1622 vdd.n2900 vdd.n2899 8.92171
R1623 vdd.n2920 vdd.n2919 8.92171
R1624 vdd.n2947 vdd.n2390 8.92171
R1625 vdd.n2391 vdd.n2377 8.92171
R1626 vdd.n2980 vdd.n2979 8.92171
R1627 vdd.n2362 vdd.n2357 8.92171
R1628 vdd.n3026 vdd.n3025 8.92171
R1629 vdd.n3062 vdd.n3061 8.92171
R1630 vdd.n3083 vdd.n3082 8.92171
R1631 vdd.n2308 vdd.n2302 8.92171
R1632 vdd.n3126 vdd.n3125 8.92171
R1633 vdd.n3146 vdd.n3145 8.92171
R1634 vdd.n3173 vdd.n2256 8.92171
R1635 vdd.n2257 vdd.n2243 8.92171
R1636 vdd.n3206 vdd.n3205 8.92171
R1637 vdd.n2228 vdd.n2223 8.92171
R1638 vdd.n3252 vdd.n3251 8.92171
R1639 vdd.n3288 vdd.n3287 8.92171
R1640 vdd.n3309 vdd.n3308 8.92171
R1641 vdd.n2174 vdd.n2168 8.92171
R1642 vdd.n3352 vdd.n3351 8.92171
R1643 vdd.n3372 vdd.n3371 8.92171
R1644 vdd.n3399 vdd.n2122 8.92171
R1645 vdd.n2123 vdd.n2109 8.92171
R1646 vdd.n3432 vdd.n3431 8.92171
R1647 vdd.n2094 vdd.n2089 8.92171
R1648 vdd.n3478 vdd.n3477 8.92171
R1649 vdd.n3514 vdd.n3513 8.92171
R1650 vdd.n3535 vdd.n3534 8.92171
R1651 vdd.n2040 vdd.n2034 8.92171
R1652 vdd.n3578 vdd.n3577 8.92171
R1653 vdd.n3598 vdd.n3597 8.92171
R1654 vdd.n3625 vdd.n1988 8.92171
R1655 vdd.n1989 vdd.n1975 8.92171
R1656 vdd.n3658 vdd.n3657 8.92171
R1657 vdd.n1960 vdd.n1955 8.92171
R1658 vdd.n3709 vdd.n3708 8.92171
R1659 vdd.n3736 vdd.n3735 8.92171
R1660 vdd.n3755 vdd.n3754 8.92171
R1661 vdd.n3774 vdd.n3773 8.92171
R1662 vdd.n3793 vdd.n3792 8.92171
R1663 vdd.n3812 vdd.n3811 8.92171
R1664 vdd.n2518 vdd.n2516 8.85203
R1665 vdd.n3738 vdd.n1886 8.77616
R1666 vdd.n3757 vdd.n1886 8.77616
R1667 vdd.n3776 vdd.n1886 8.77616
R1668 vdd.n3795 vdd.n1886 8.77616
R1669 vdd.n2938 vdd.n1942 8.77616
R1670 vdd.n2975 vdd.n1942 8.77616
R1671 vdd.n3009 vdd.n1942 8.77616
R1672 vdd.n3164 vdd.n1942 8.77616
R1673 vdd.n3201 vdd.n1942 8.77616
R1674 vdd.n3235 vdd.n1942 8.77616
R1675 vdd.n3390 vdd.n1942 8.77616
R1676 vdd.n3427 vdd.n1942 8.77616
R1677 vdd.n3461 vdd.n1942 8.77616
R1678 vdd.n3616 vdd.n1942 8.77616
R1679 vdd.n3653 vdd.n1942 8.77616
R1680 vdd.n3687 vdd.n1942 8.77616
R1681 vdd.n3601 vdd.n1942 8.77616
R1682 vdd.n3375 vdd.n1942 8.77616
R1683 vdd.n3149 vdd.n1942 8.77616
R1684 vdd.n2923 vdd.n1942 8.77616
R1685 vdd.n2452 vdd.n1942 8.77616
R1686 vdd.n2677 vdd.n2520 8.66641
R1687 vdd.n2590 vdd 8.58587
R1688 vdd.t2 vdd.n2605 7.65151
R1689 vdd.t27 vdd.t76 7.65151
R1690 vdd.n2624 vdd.t21 7.65151
R1691 vdd.n2531 vdd.n2529 7.48074
R1692 vdd.n2709 vdd.n2708 7.13332
R1693 vdd.n2683 vdd.n2682 6.84721
R1694 vdd.n673 vdd.n666 6.67284
R1695 vdd.n2704 vdd.n2703 5.8631
R1696 vdd.n668 vdd.n666 5.85582
R1697 vdd.n2703 vdd.n2539 5.66768
R1698 vdd.n2603 vdd.n2577 5.63495
R1699 vdd.n2597 vdd.n2571 5.63495
R1700 vdd.n3814 vdd.n1886 5.63319
R1701 vdd.n2415 vdd.n1942 5.63319
R1702 vdd.n3028 vdd.n1942 5.63319
R1703 vdd.n2977 vdd.n1942 5.63319
R1704 vdd.n2941 vdd.n1942 5.63319
R1705 vdd.n2281 vdd.n1942 5.63319
R1706 vdd.n3254 vdd.n1942 5.63319
R1707 vdd.n3203 vdd.n1942 5.63319
R1708 vdd.n3167 vdd.n1942 5.63319
R1709 vdd.n2147 vdd.n1942 5.63319
R1710 vdd.n3480 vdd.n1942 5.63319
R1711 vdd.n3429 vdd.n1942 5.63319
R1712 vdd.n3393 vdd.n1942 5.63319
R1713 vdd.n2013 vdd.n1942 5.63319
R1714 vdd.n3655 vdd.n1942 5.63319
R1715 vdd.n3619 vdd.n1942 5.63319
R1716 vdd.n2662 vdd.n2661 5.57371
R1717 vdd.n2611 vdd.n2610 5.51246
R1718 vdd.n2642 vdd.n2626 5.51246
R1719 vdd.n2680 vdd.n2550 5.51246
R1720 vdd.n2618 vdd.n2562 5.38997
R1721 vdd.n2673 vdd.n2553 5.38997
R1722 vdd.n2717 vdd.n2525 5.38021
R1723 vdd.n2714 vdd.n2713 5.38021
R1724 vdd.n2599 vdd.n2598 5.32873
R1725 vdd.n2628 vdd.n2627 5.26749
R1726 vdd.n2649 vdd.n2648 5.20624
R1727 vdd.n2832 vdd.n1942 5.1329
R1728 vdd.n3711 vdd.n1942 5.1329
R1729 vdd.n2621 vdd.t85 5.10117
R1730 vdd.n2810 vdd.t55 5.05206
R1731 vdd.t47 vdd.n696 4.95579
R1732 vdd.n2586 vdd.n2578 4.77029
R1733 vdd.n2588 vdd.n2578 4.77029
R1734 vdd.n2507 vdd.t87 4.74591
R1735 vdd.n2667 vdd.n2554 4.71629
R1736 vdd.n675 vdd.n664 4.7039
R1737 vdd.n2681 vdd.n2524 4.67925
R1738 vdd.n674 vdd.n673 4.6505
R1739 vdd.n668 vdd.n665 4.6505
R1740 vdd.n1837 vdd.n1836 4.6505
R1741 vdd.n1805 vdd.n1804 4.6505
R1742 vdd.n2724 vdd.n2723 4.6505
R1743 vdd.n2517 vdd.n2515 4.6505
R1744 vdd.n2703 vdd.n2702 4.6505
R1745 vdd.n2701 vdd.n2700 4.6505
R1746 vdd.n2532 vdd.n2530 4.6505
R1747 vdd.n2710 vdd.n2709 4.6505
R1748 vdd.n2712 vdd.n2711 4.6505
R1749 vdd.n2715 vdd.n2714 4.6505
R1750 vdd.n2717 vdd.n2716 4.6505
R1751 vdd.n2684 vdd.n2683 4.6505
R1752 vdd.n2588 vdd.n2587 4.6505
R1753 vdd.n2601 vdd.n2577 4.6505
R1754 vdd.n2587 vdd.n2586 4.6505
R1755 vdd.n2603 vdd.n2576 4.6505
R1756 vdd.n2593 vdd.n2577 4.6505
R1757 vdd.n2599 vdd.n2594 4.6505
R1758 vdd.n2597 vdd.n2596 4.6505
R1759 vdd.n2595 vdd.n2571 4.6505
R1760 vdd.n2614 vdd.n2569 4.6505
R1761 vdd.n2651 vdd.n2650 4.6505
R1762 vdd.n2629 vdd.n2563 4.6505
R1763 vdd.n2638 vdd.n2637 4.6505
R1764 vdd.n2641 vdd.n2640 4.6505
R1765 vdd.n2659 vdd.n2556 4.6505
R1766 vdd.n2662 vdd.n2555 4.6505
R1767 vdd.n2673 vdd.n2672 4.6505
R1768 vdd.n2670 vdd.n2669 4.6505
R1769 vdd.n2680 vdd.n2548 4.6505
R1770 vdd.n2668 vdd.n2665 4.6505
R1771 vdd.n2671 vdd.n2554 4.6505
R1772 vdd.n2664 vdd.n2663 4.6505
R1773 vdd.n2661 vdd.n2660 4.6505
R1774 vdd.n2628 vdd.n2557 4.6505
R1775 vdd.n2639 vdd.n2626 4.6505
R1776 vdd.n2633 vdd.n2630 4.6505
R1777 vdd.n2649 vdd.n2561 4.6505
R1778 vdd.n2615 vdd.n2614 4.6505
R1779 vdd.n2571 vdd.n2570 4.6505
R1780 vdd.n2597 vdd.n2589 4.6505
R1781 vdd.n2600 vdd.n2599 4.6505
R1782 vdd.n2603 vdd.n2602 4.6505
R1783 vdd.n2681 vdd.n2526 4.6505
R1784 vdd.n2788 vdd.n2787 4.6505
R1785 vdd.n2774 vdd.n2765 4.6505
R1786 vdd.n701 vdd.n607 4.54027
R1787 vdd.n1682 vdd.n1681 4.54027
R1788 vdd.n2830 vdd.n2463 4.54027
R1789 vdd.n3714 vdd.n3713 4.54027
R1790 vdd.n658 vdd.n657 4.52882
R1791 vdd.n2737 vdd.n2736 4.52882
R1792 vdd.n601 vdd.n599 4.5005
R1793 vdd.n591 vdd.n590 4.5005
R1794 vdd.n728 vdd.n591 4.5005
R1795 vdd.n732 vdd.n731 4.5005
R1796 vdd.n718 vdd.n717 4.5005
R1797 vdd.n813 vdd.n812 4.5005
R1798 vdd.n811 vdd.n544 4.5005
R1799 vdd.n534 vdd.n533 4.5005
R1800 vdd.n915 vdd.n914 4.5005
R1801 vdd.n917 vdd.n473 4.5005
R1802 vdd.n969 vdd.n968 4.5005
R1803 vdd.n1064 vdd.n1063 4.5005
R1804 vdd.n1062 vdd.n410 4.5005
R1805 vdd.n400 vdd.n399 4.5005
R1806 vdd.n1166 vdd.n1165 4.5005
R1807 vdd.n1168 vdd.n339 4.5005
R1808 vdd.n1220 vdd.n1219 4.5005
R1809 vdd.n1315 vdd.n1314 4.5005
R1810 vdd.n1313 vdd.n276 4.5005
R1811 vdd.n266 vdd.n265 4.5005
R1812 vdd.n1417 vdd.n1416 4.5005
R1813 vdd.n1419 vdd.n205 4.5005
R1814 vdd.n1471 vdd.n1470 4.5005
R1815 vdd.n1566 vdd.n1565 4.5005
R1816 vdd.n1564 vdd.n142 4.5005
R1817 vdd.n133 vdd.n132 4.5005
R1818 vdd.n84 vdd.n83 4.5005
R1819 vdd.n101 vdd.n99 4.5005
R1820 vdd.n1651 vdd.n89 4.5005
R1821 vdd.n1651 vdd.n1650 4.5005
R1822 vdd.n1640 vdd.n1639 4.5005
R1823 vdd.n1622 vdd.n1621 4.5005
R1824 vdd.n1620 vdd.n97 4.5005
R1825 vdd.n97 vdd.n96 4.5005
R1826 vdd.n1624 vdd.n1623 4.5005
R1827 vdd.n1605 vdd.n116 4.5005
R1828 vdd.n1607 vdd.n1606 4.5005
R1829 vdd.n1607 vdd.n115 4.5005
R1830 vdd.n126 vdd.n117 4.5005
R1831 vdd.n1583 vdd.n1582 4.5005
R1832 vdd.n125 vdd.n123 4.5005
R1833 vdd.n127 vdd.n125 4.5005
R1834 vdd.n1668 vdd.n1667 4.5005
R1835 vdd.n1666 vdd.n74 4.5005
R1836 vdd.n76 vdd.n74 4.5005
R1837 vdd.n1571 vdd.n137 4.5005
R1838 vdd.n1571 vdd.n1570 4.5005
R1839 vdd.n1550 vdd.n1549 4.5005
R1840 vdd.n170 vdd.n159 4.5005
R1841 vdd.n152 vdd.n151 4.5005
R1842 vdd.n151 vdd.n150 4.5005
R1843 vdd.n1524 vdd.n1523 4.5005
R1844 vdd.n1511 vdd.n166 4.5005
R1845 vdd.n1526 vdd.n1525 4.5005
R1846 vdd.n1526 vdd.n165 4.5005
R1847 vdd.n1509 vdd.n1508 4.5005
R1848 vdd.n1486 vdd.n182 4.5005
R1849 vdd.n176 vdd.n175 4.5005
R1850 vdd.n177 vdd.n176 4.5005
R1851 vdd.n1485 vdd.n1484 4.5005
R1852 vdd.n199 vdd.n197 4.5005
R1853 vdd.n189 vdd.n188 4.5005
R1854 vdd.n1481 vdd.n189 4.5005
R1855 vdd.n153 vdd.n145 4.5005
R1856 vdd.n1563 vdd.n141 4.5005
R1857 vdd.n141 vdd.n140 4.5005
R1858 vdd.n198 vdd.n196 4.5005
R1859 vdd.n196 vdd.n195 4.5005
R1860 vdd.n1409 vdd.n1408 4.5005
R1861 vdd.n1397 vdd.n1396 4.5005
R1862 vdd.n225 vdd.n224 4.5005
R1863 vdd.n1393 vdd.n224 4.5005
R1864 vdd.n230 vdd.n229 4.5005
R1865 vdd.n1375 vdd.n1374 4.5005
R1866 vdd.n237 vdd.n236 4.5005
R1867 vdd.n236 vdd.n235 4.5005
R1868 vdd.n243 vdd.n242 4.5005
R1869 vdd.n252 vdd.n250 4.5005
R1870 vdd.n1361 vdd.n1360 4.5005
R1871 vdd.n1361 vdd.n249 4.5005
R1872 vdd.n1350 vdd.n1349 4.5005
R1873 vdd.n1337 vdd.n1336 4.5005
R1874 vdd.n1335 vdd.n258 4.5005
R1875 vdd.n260 vdd.n258 4.5005
R1876 vdd.n217 vdd.n216 4.5005
R1877 vdd.n1434 vdd.n1433 4.5005
R1878 vdd.n1434 vdd.n210 4.5005
R1879 vdd.n1320 vdd.n271 4.5005
R1880 vdd.n1320 vdd.n1319 4.5005
R1881 vdd.n1299 vdd.n1298 4.5005
R1882 vdd.n304 vdd.n293 4.5005
R1883 vdd.n286 vdd.n285 4.5005
R1884 vdd.n285 vdd.n284 4.5005
R1885 vdd.n1273 vdd.n1272 4.5005
R1886 vdd.n1260 vdd.n300 4.5005
R1887 vdd.n1275 vdd.n1274 4.5005
R1888 vdd.n1275 vdd.n299 4.5005
R1889 vdd.n1258 vdd.n1257 4.5005
R1890 vdd.n1235 vdd.n316 4.5005
R1891 vdd.n310 vdd.n309 4.5005
R1892 vdd.n311 vdd.n310 4.5005
R1893 vdd.n1234 vdd.n1233 4.5005
R1894 vdd.n333 vdd.n331 4.5005
R1895 vdd.n323 vdd.n322 4.5005
R1896 vdd.n1230 vdd.n323 4.5005
R1897 vdd.n287 vdd.n279 4.5005
R1898 vdd.n1312 vdd.n275 4.5005
R1899 vdd.n275 vdd.n274 4.5005
R1900 vdd.n332 vdd.n330 4.5005
R1901 vdd.n330 vdd.n329 4.5005
R1902 vdd.n1158 vdd.n1157 4.5005
R1903 vdd.n1146 vdd.n1145 4.5005
R1904 vdd.n359 vdd.n358 4.5005
R1905 vdd.n1142 vdd.n358 4.5005
R1906 vdd.n364 vdd.n363 4.5005
R1907 vdd.n1124 vdd.n1123 4.5005
R1908 vdd.n371 vdd.n370 4.5005
R1909 vdd.n370 vdd.n369 4.5005
R1910 vdd.n377 vdd.n376 4.5005
R1911 vdd.n386 vdd.n384 4.5005
R1912 vdd.n1110 vdd.n1109 4.5005
R1913 vdd.n1110 vdd.n383 4.5005
R1914 vdd.n1099 vdd.n1098 4.5005
R1915 vdd.n1086 vdd.n1085 4.5005
R1916 vdd.n1084 vdd.n392 4.5005
R1917 vdd.n394 vdd.n392 4.5005
R1918 vdd.n351 vdd.n350 4.5005
R1919 vdd.n1183 vdd.n1182 4.5005
R1920 vdd.n1183 vdd.n344 4.5005
R1921 vdd.n1069 vdd.n405 4.5005
R1922 vdd.n1069 vdd.n1068 4.5005
R1923 vdd.n1048 vdd.n1047 4.5005
R1924 vdd.n438 vdd.n427 4.5005
R1925 vdd.n420 vdd.n419 4.5005
R1926 vdd.n419 vdd.n418 4.5005
R1927 vdd.n1022 vdd.n1021 4.5005
R1928 vdd.n1009 vdd.n434 4.5005
R1929 vdd.n1024 vdd.n1023 4.5005
R1930 vdd.n1024 vdd.n433 4.5005
R1931 vdd.n1007 vdd.n1006 4.5005
R1932 vdd.n984 vdd.n450 4.5005
R1933 vdd.n444 vdd.n443 4.5005
R1934 vdd.n445 vdd.n444 4.5005
R1935 vdd.n983 vdd.n982 4.5005
R1936 vdd.n467 vdd.n465 4.5005
R1937 vdd.n457 vdd.n456 4.5005
R1938 vdd.n979 vdd.n457 4.5005
R1939 vdd.n421 vdd.n413 4.5005
R1940 vdd.n1061 vdd.n409 4.5005
R1941 vdd.n409 vdd.n408 4.5005
R1942 vdd.n466 vdd.n464 4.5005
R1943 vdd.n464 vdd.n463 4.5005
R1944 vdd.n907 vdd.n906 4.5005
R1945 vdd.n895 vdd.n894 4.5005
R1946 vdd.n493 vdd.n492 4.5005
R1947 vdd.n891 vdd.n492 4.5005
R1948 vdd.n498 vdd.n497 4.5005
R1949 vdd.n873 vdd.n872 4.5005
R1950 vdd.n505 vdd.n504 4.5005
R1951 vdd.n504 vdd.n503 4.5005
R1952 vdd.n511 vdd.n510 4.5005
R1953 vdd.n520 vdd.n518 4.5005
R1954 vdd.n859 vdd.n858 4.5005
R1955 vdd.n859 vdd.n517 4.5005
R1956 vdd.n848 vdd.n847 4.5005
R1957 vdd.n835 vdd.n834 4.5005
R1958 vdd.n833 vdd.n526 4.5005
R1959 vdd.n528 vdd.n526 4.5005
R1960 vdd.n485 vdd.n484 4.5005
R1961 vdd.n932 vdd.n931 4.5005
R1962 vdd.n932 vdd.n478 4.5005
R1963 vdd.n818 vdd.n539 4.5005
R1964 vdd.n818 vdd.n817 4.5005
R1965 vdd.n797 vdd.n796 4.5005
R1966 vdd.n572 vdd.n561 4.5005
R1967 vdd.n554 vdd.n553 4.5005
R1968 vdd.n553 vdd.n552 4.5005
R1969 vdd.n771 vdd.n770 4.5005
R1970 vdd.n758 vdd.n568 4.5005
R1971 vdd.n773 vdd.n772 4.5005
R1972 vdd.n773 vdd.n567 4.5005
R1973 vdd.n756 vdd.n755 4.5005
R1974 vdd.n733 vdd.n584 4.5005
R1975 vdd.n578 vdd.n577 4.5005
R1976 vdd.n579 vdd.n578 4.5005
R1977 vdd.n555 vdd.n547 4.5005
R1978 vdd.n810 vdd.n543 4.5005
R1979 vdd.n543 vdd.n542 4.5005
R1980 vdd.n600 vdd.n598 4.5005
R1981 vdd.n598 vdd.n597 4.5005
R1982 vdd.n1698 vdd.n1697 4.5005
R1983 vdd.n61 vdd.n59 4.5005
R1984 vdd.n63 vdd.n61 4.5005
R1985 vdd.n62 vdd.n53 4.5005
R1986 vdd.n69 vdd.n68 4.5005
R1987 vdd.n12 vdd.n5 4.5005
R1988 vdd.n21 vdd.n20 4.5005
R1989 vdd.n37 vdd.n35 4.5005
R1990 vdd.n1766 vdd.n25 4.5005
R1991 vdd.n1766 vdd.n1765 4.5005
R1992 vdd.n1755 vdd.n1754 4.5005
R1993 vdd.n1737 vdd.n1736 4.5005
R1994 vdd.n1735 vdd.n33 4.5005
R1995 vdd.n33 vdd.n32 4.5005
R1996 vdd.n1739 vdd.n1738 4.5005
R1997 vdd.n1720 vdd.n52 4.5005
R1998 vdd.n1722 vdd.n1721 4.5005
R1999 vdd.n1722 vdd.n51 4.5005
R2000 vdd.n1778 vdd.n1777 4.5005
R2001 vdd.n11 vdd.n9 4.5005
R2002 vdd.n13 vdd.n11 4.5005
R2003 vdd.n2461 vdd.n2460 4.5005
R2004 vdd.n2462 vdd.n2461 4.5005
R2005 vdd.n2839 vdd.n2838 4.5005
R2006 vdd.n2860 vdd.n2859 4.5005
R2007 vdd.n2411 vdd.n2410 4.5005
R2008 vdd.n2419 vdd.n2403 4.5005
R2009 vdd.n3046 vdd.n2331 4.5005
R2010 vdd.n2343 vdd.n2336 4.5005
R2011 vdd.n3023 vdd.n3022 4.5005
R2012 vdd.n2342 vdd.n2340 4.5005
R2013 vdd.n2344 vdd.n2342 4.5005
R2014 vdd.n3002 vdd.n3001 4.5005
R2015 vdd.n2984 vdd.n2983 4.5005
R2016 vdd.n2982 vdd.n2360 4.5005
R2017 vdd.n2360 vdd.n2359 4.5005
R2018 vdd.n2967 vdd.n2966 4.5005
R2019 vdd.n2950 vdd.n2949 4.5005
R2020 vdd.n2389 vdd.n2387 4.5005
R2021 vdd.n2946 vdd.n2389 4.5005
R2022 vdd.n2388 vdd.n2386 4.5005
R2023 vdd.n2409 vdd.n2408 4.5005
R2024 vdd.n2396 vdd.n2395 4.5005
R2025 vdd.n2395 vdd.n2394 4.5005
R2026 vdd.n2986 vdd.n2985 4.5005
R2027 vdd.n2969 vdd.n2968 4.5005
R2028 vdd.n2971 vdd.n2970 4.5005
R2029 vdd.n2972 vdd.n2971 4.5005
R2030 vdd.n2349 vdd.n2348 4.5005
R2031 vdd.n2366 vdd.n2364 4.5005
R2032 vdd.n2355 vdd.n2353 4.5005
R2033 vdd.n2356 vdd.n2355 4.5005
R2034 vdd.n2277 vdd.n2276 4.5005
R2035 vdd.n2285 vdd.n2269 4.5005
R2036 vdd.n3272 vdd.n2197 4.5005
R2037 vdd.n2209 vdd.n2202 4.5005
R2038 vdd.n3249 vdd.n3248 4.5005
R2039 vdd.n2208 vdd.n2206 4.5005
R2040 vdd.n2210 vdd.n2208 4.5005
R2041 vdd.n3228 vdd.n3227 4.5005
R2042 vdd.n3210 vdd.n3209 4.5005
R2043 vdd.n3208 vdd.n2226 4.5005
R2044 vdd.n2226 vdd.n2225 4.5005
R2045 vdd.n3193 vdd.n3192 4.5005
R2046 vdd.n3176 vdd.n3175 4.5005
R2047 vdd.n2255 vdd.n2253 4.5005
R2048 vdd.n3172 vdd.n2255 4.5005
R2049 vdd.n2254 vdd.n2252 4.5005
R2050 vdd.n2275 vdd.n2274 4.5005
R2051 vdd.n2262 vdd.n2261 4.5005
R2052 vdd.n2261 vdd.n2260 4.5005
R2053 vdd.n3212 vdd.n3211 4.5005
R2054 vdd.n3195 vdd.n3194 4.5005
R2055 vdd.n3197 vdd.n3196 4.5005
R2056 vdd.n3198 vdd.n3197 4.5005
R2057 vdd.n2215 vdd.n2214 4.5005
R2058 vdd.n2232 vdd.n2230 4.5005
R2059 vdd.n2221 vdd.n2219 4.5005
R2060 vdd.n2222 vdd.n2221 4.5005
R2061 vdd.n2143 vdd.n2142 4.5005
R2062 vdd.n2151 vdd.n2135 4.5005
R2063 vdd.n3498 vdd.n2063 4.5005
R2064 vdd.n2075 vdd.n2068 4.5005
R2065 vdd.n3475 vdd.n3474 4.5005
R2066 vdd.n2074 vdd.n2072 4.5005
R2067 vdd.n2076 vdd.n2074 4.5005
R2068 vdd.n3454 vdd.n3453 4.5005
R2069 vdd.n3436 vdd.n3435 4.5005
R2070 vdd.n3434 vdd.n2092 4.5005
R2071 vdd.n2092 vdd.n2091 4.5005
R2072 vdd.n3419 vdd.n3418 4.5005
R2073 vdd.n3402 vdd.n3401 4.5005
R2074 vdd.n2121 vdd.n2119 4.5005
R2075 vdd.n3398 vdd.n2121 4.5005
R2076 vdd.n2120 vdd.n2118 4.5005
R2077 vdd.n2141 vdd.n2140 4.5005
R2078 vdd.n2128 vdd.n2127 4.5005
R2079 vdd.n2127 vdd.n2126 4.5005
R2080 vdd.n3438 vdd.n3437 4.5005
R2081 vdd.n3421 vdd.n3420 4.5005
R2082 vdd.n3423 vdd.n3422 4.5005
R2083 vdd.n3424 vdd.n3423 4.5005
R2084 vdd.n2081 vdd.n2080 4.5005
R2085 vdd.n2098 vdd.n2096 4.5005
R2086 vdd.n2087 vdd.n2085 4.5005
R2087 vdd.n2088 vdd.n2087 4.5005
R2088 vdd.n2009 vdd.n2008 4.5005
R2089 vdd.n2017 vdd.n2001 4.5005
R2090 vdd.n3706 vdd.n3705 4.5005
R2091 vdd.n3680 vdd.n3679 4.5005
R2092 vdd.n3662 vdd.n3661 4.5005
R2093 vdd.n3660 vdd.n1958 4.5005
R2094 vdd.n1958 vdd.n1957 4.5005
R2095 vdd.n3645 vdd.n3644 4.5005
R2096 vdd.n3628 vdd.n3627 4.5005
R2097 vdd.n1987 vdd.n1985 4.5005
R2098 vdd.n3624 vdd.n1987 4.5005
R2099 vdd.n1986 vdd.n1984 4.5005
R2100 vdd.n2007 vdd.n2006 4.5005
R2101 vdd.n1994 vdd.n1993 4.5005
R2102 vdd.n1993 vdd.n1992 4.5005
R2103 vdd.n3664 vdd.n3663 4.5005
R2104 vdd.n3647 vdd.n3646 4.5005
R2105 vdd.n3649 vdd.n3648 4.5005
R2106 vdd.n3650 vdd.n3649 4.5005
R2107 vdd.n1946 vdd.n1945 4.5005
R2108 vdd.n1964 vdd.n1962 4.5005
R2109 vdd.n1953 vdd.n1951 4.5005
R2110 vdd.n1954 vdd.n1953 4.5005
R2111 vdd.n3704 vdd.n1939 4.5005
R2112 vdd.n1941 vdd.n1939 4.5005
R2113 vdd.n3518 vdd.n2052 4.5005
R2114 vdd.n3595 vdd.n3594 4.5005
R2115 vdd.n2028 vdd.n2022 4.5005
R2116 vdd.n2016 vdd.n2015 4.5005
R2117 vdd.n2015 vdd.n2014 4.5005
R2118 vdd.n3575 vdd.n3574 4.5005
R2119 vdd.n2042 vdd.n2033 4.5005
R2120 vdd.n2027 vdd.n2026 4.5005
R2121 vdd.n2026 vdd.n2025 4.5005
R2122 vdd.n3553 vdd.n3552 4.5005
R2123 vdd.n3540 vdd.n2038 4.5005
R2124 vdd.n3555 vdd.n3554 4.5005
R2125 vdd.n3555 vdd.n2037 4.5005
R2126 vdd.n2048 vdd.n2047 4.5005
R2127 vdd.n2049 vdd.n2048 4.5005
R2128 vdd.n3538 vdd.n3537 4.5005
R2129 vdd.n2002 vdd.n2000 4.5005
R2130 vdd.n2012 vdd.n2002 4.5005
R2131 vdd.n2059 vdd.n2058 4.5005
R2132 vdd.n2060 vdd.n2059 4.5005
R2133 vdd.n3517 vdd.n3516 4.5005
R2134 vdd.n3292 vdd.n2186 4.5005
R2135 vdd.n3369 vdd.n3368 4.5005
R2136 vdd.n2162 vdd.n2156 4.5005
R2137 vdd.n2150 vdd.n2149 4.5005
R2138 vdd.n2149 vdd.n2148 4.5005
R2139 vdd.n3349 vdd.n3348 4.5005
R2140 vdd.n2176 vdd.n2167 4.5005
R2141 vdd.n2161 vdd.n2160 4.5005
R2142 vdd.n2160 vdd.n2159 4.5005
R2143 vdd.n3327 vdd.n3326 4.5005
R2144 vdd.n3314 vdd.n2172 4.5005
R2145 vdd.n3329 vdd.n3328 4.5005
R2146 vdd.n3329 vdd.n2171 4.5005
R2147 vdd.n2182 vdd.n2181 4.5005
R2148 vdd.n2183 vdd.n2182 4.5005
R2149 vdd.n3312 vdd.n3311 4.5005
R2150 vdd.n2136 vdd.n2134 4.5005
R2151 vdd.n2146 vdd.n2136 4.5005
R2152 vdd.n2193 vdd.n2192 4.5005
R2153 vdd.n2194 vdd.n2193 4.5005
R2154 vdd.n3291 vdd.n3290 4.5005
R2155 vdd.n3066 vdd.n2320 4.5005
R2156 vdd.n3143 vdd.n3142 4.5005
R2157 vdd.n2296 vdd.n2290 4.5005
R2158 vdd.n2284 vdd.n2283 4.5005
R2159 vdd.n2283 vdd.n2282 4.5005
R2160 vdd.n3123 vdd.n3122 4.5005
R2161 vdd.n2310 vdd.n2301 4.5005
R2162 vdd.n2295 vdd.n2294 4.5005
R2163 vdd.n2294 vdd.n2293 4.5005
R2164 vdd.n3101 vdd.n3100 4.5005
R2165 vdd.n3088 vdd.n2306 4.5005
R2166 vdd.n3103 vdd.n3102 4.5005
R2167 vdd.n3103 vdd.n2305 4.5005
R2168 vdd.n2316 vdd.n2315 4.5005
R2169 vdd.n2317 vdd.n2316 4.5005
R2170 vdd.n3086 vdd.n3085 4.5005
R2171 vdd.n2270 vdd.n2268 4.5005
R2172 vdd.n2280 vdd.n2270 4.5005
R2173 vdd.n2327 vdd.n2326 4.5005
R2174 vdd.n2328 vdd.n2327 4.5005
R2175 vdd.n3065 vdd.n3064 4.5005
R2176 vdd.n2862 vdd.n2440 4.5005
R2177 vdd.n2917 vdd.n2916 4.5005
R2178 vdd.n2430 vdd.n2424 4.5005
R2179 vdd.n2418 vdd.n2417 4.5005
R2180 vdd.n2417 vdd.n2416 4.5005
R2181 vdd.n2897 vdd.n2896 4.5005
R2182 vdd.n2444 vdd.n2435 4.5005
R2183 vdd.n2429 vdd.n2428 4.5005
R2184 vdd.n2428 vdd.n2427 4.5005
R2185 vdd.n2877 vdd.n2876 4.5005
R2186 vdd.n2877 vdd.n2439 4.5005
R2187 vdd.n2875 vdd.n2874 4.5005
R2188 vdd.n2404 vdd.n2402 4.5005
R2189 vdd.n2414 vdd.n2404 4.5005
R2190 vdd.n2450 vdd.n2449 4.5005
R2191 vdd.n2451 vdd.n2450 4.5005
R2192 vdd.n2840 vdd.n2454 4.5005
R2193 vdd.n3809 vdd.n3808 4.5005
R2194 vdd.n1881 vdd.n1879 4.5005
R2195 vdd.n1883 vdd.n1881 4.5005
R2196 vdd.n1882 vdd.n1875 4.5005
R2197 vdd.n1934 vdd.n1933 4.5005
R2198 vdd.n1923 vdd.n1922 4.5005
R2199 vdd.n3733 vdd.n3732 4.5005
R2200 vdd.n1929 vdd.n1927 4.5005
R2201 vdd.n1930 vdd.n1929 4.5005
R2202 vdd.n1912 vdd.n1911 4.5005
R2203 vdd.n3752 vdd.n3751 4.5005
R2204 vdd.n1918 vdd.n1916 4.5005
R2205 vdd.n1919 vdd.n1918 4.5005
R2206 vdd.n1901 vdd.n1900 4.5005
R2207 vdd.n3771 vdd.n3770 4.5005
R2208 vdd.n1907 vdd.n1905 4.5005
R2209 vdd.n1908 vdd.n1907 4.5005
R2210 vdd.n1890 vdd.n1889 4.5005
R2211 vdd.n3790 vdd.n3789 4.5005
R2212 vdd.n1896 vdd.n1894 4.5005
R2213 vdd.n1897 vdd.n1896 4.5005
R2214 vdd.n2778 vdd.n2777 4.5005
R2215 vdd.n2762 vdd.n2760 4.5005
R2216 vdd.n2763 vdd.n2761 4.5005
R2217 vdd.n2801 vdd.n2800 4.43667
R2218 vdd.t14 vdd.t29 4.33345
R2219 vdd vdd.n1870 4.29567
R2220 vdd vdd.n1886 4.28667
R2221 vdd.n2584 vdd 4.16509
R2222 vdd.n695 vdd.n609 3.67129
R2223 vdd.n2811 vdd.n2810 3.52129
R2224 vdd.n2770 vdd.n2766 3.46788
R2225 vdd.n2799 vdd.n2798 3.46651
R2226 vdd.n650 vdd.n649 3.46323
R2227 vdd.n2691 vdd.n2690 3.46323
R2228 vdd.n2657 vdd.n2558 3.46323
R2229 vdd.n2686 vdd.n2547 3.46323
R2230 vdd.n2698 vdd.n2540 3.46323
R2231 vdd.n2726 vdd.n2514 3.46323
R2232 vdd.n2744 vdd.n2743 3.46323
R2233 vdd.n659 vdd.n653 3.46321
R2234 vdd.n2738 vdd.n2732 3.46321
R2235 vdd.n693 vdd.n611 3.45407
R2236 vdd.n646 vdd.n645 3.45407
R2237 vdd.n639 vdd.n638 3.45407
R2238 vdd.n633 vdd.n628 3.45407
R2239 vdd.n624 vdd.n623 3.45407
R2240 vdd.n2752 vdd.n2510 3.45407
R2241 vdd.n2817 vdd.n2816 3.45407
R2242 vdd.n2505 vdd.n2472 3.45407
R2243 vdd.n2487 vdd.n2477 3.45407
R2244 vdd.n2495 vdd.n2494 3.45407
R2245 vdd.n612 vdd.n610 3.45149
R2246 vdd.n643 vdd.n641 3.45149
R2247 vdd.n636 vdd.n630 3.45149
R2248 vdd.n632 vdd.n626 3.45149
R2249 vdd.n621 vdd.n619 3.45149
R2250 vdd.n2511 vdd.n2509 3.45149
R2251 vdd.n2814 vdd.n2468 3.45149
R2252 vdd.n2473 vdd.n2471 3.45149
R2253 vdd.n2486 vdd.n2475 3.45149
R2254 vdd.n2492 vdd.n2479 3.45149
R2255 vdd.n1689 vdd.n1685 3.42985
R2256 vdd.n3724 vdd.n3717 3.42985
R2257 vdd.n2781 vdd.n2763 3.4257
R2258 vdd.n2656 vdd.n2560 3.42509
R2259 vdd.n2688 vdd.n2687 3.42509
R2260 vdd.n2697 vdd.n2542 3.42509
R2261 vdd.n2693 vdd.n2692 3.42509
R2262 vdd.n2728 vdd.n2727 3.42476
R2263 vdd.n1868 vdd.n1867 3.42443
R2264 vdd.n3833 vdd.n3832 3.42443
R2265 vdd.n615 vdd.n607 3.42376
R2266 vdd.n1683 vdd.n1682 3.42376
R2267 vdd.n2822 vdd.n2463 3.42376
R2268 vdd.n3715 vdd.n3714 3.42376
R2269 vdd.n655 vdd.n652 3.41853
R2270 vdd.n2734 vdd.n2731 3.41853
R2271 vdd.n2779 vdd.n2778 3.41388
R2272 vdd.n1684 vdd.n1683 3.41326
R2273 vdd.n3716 vdd.n3715 3.41326
R2274 vdd.n616 vdd.n615 3.41257
R2275 vdd.n2822 vdd.n2821 3.41257
R2276 vdd.n2653 vdd.n2558 3.41222
R2277 vdd.n2559 vdd.n2547 3.41222
R2278 vdd.n2694 vdd.n2540 3.41222
R2279 vdd.n2690 vdd.n2689 3.41222
R2280 vdd.n689 vdd.n611 3.41218
R2281 vdd.n650 vdd.n647 3.41218
R2282 vdd.n646 vdd.n640 3.41218
R2283 vdd.n639 vdd.n629 3.41218
R2284 vdd.n628 vdd.n625 3.41218
R2285 vdd.n624 vdd.n618 3.41218
R2286 vdd.n2541 vdd.n2514 3.41218
R2287 vdd.n2744 vdd.n2742 3.41218
R2288 vdd.n2748 vdd.n2510 3.41218
R2289 vdd.n2817 vdd.n2467 3.41218
R2290 vdd.n2501 vdd.n2472 3.41218
R2291 vdd.n2477 vdd.n2474 3.41218
R2292 vdd.n2495 vdd.n2478 3.41218
R2293 vdd.n654 vdd.n651 3.41162
R2294 vdd.n2733 vdd.n2730 3.41162
R2295 vdd.n703 vdd.n702 3.4105
R2296 vdd.n1604 vdd.n1603 3.4105
R2297 vdd.n1596 vdd.n1595 3.4105
R2298 vdd.n108 vdd.n104 3.4105
R2299 vdd.n119 vdd.n107 3.4105
R2300 vdd.n1638 vdd.n1637 3.4105
R2301 vdd.n1631 vdd.n98 3.4105
R2302 vdd.n1665 vdd.n1664 3.4105
R2303 vdd.n1654 vdd.n1653 3.4105
R2304 vdd.n1658 vdd.n75 3.4105
R2305 vdd.n1581 vdd.n1580 3.4105
R2306 vdd.n1574 vdd.n1573 3.4105
R2307 vdd.n1469 vdd.n1468 3.4105
R2308 vdd.n1465 vdd.n1464 3.4105
R2309 vdd.n1488 vdd.n1487 3.4105
R2310 vdd.n1496 vdd.n1495 3.4105
R2311 vdd.n1510 vdd.n173 3.4105
R2312 vdd.n1515 vdd.n167 3.4105
R2313 vdd.n1522 vdd.n1521 3.4105
R2314 vdd.n1538 vdd.n1537 3.4105
R2315 vdd.n1548 vdd.n1547 3.4105
R2316 vdd.n1562 vdd.n144 3.4105
R2317 vdd.n1421 vdd.n1420 3.4105
R2318 vdd.n1456 vdd.n1455 3.4105
R2319 vdd.n1352 vdd.n1351 3.4105
R2320 vdd.n1327 vdd.n259 3.4105
R2321 vdd.n1377 vdd.n1376 3.4105
R2322 vdd.n1359 vdd.n1358 3.4105
R2323 vdd.n1399 vdd.n1398 3.4105
R2324 vdd.n1384 vdd.n1383 3.4105
R2325 vdd.n1411 vdd.n1410 3.4105
R2326 vdd.n1406 vdd.n1405 3.4105
R2327 vdd.n1418 vdd.n1415 3.4105
R2328 vdd.n1432 vdd.n1431 3.4105
R2329 vdd.n1334 vdd.n1333 3.4105
R2330 vdd.n1323 vdd.n1322 3.4105
R2331 vdd.n1218 vdd.n1217 3.4105
R2332 vdd.n1214 vdd.n1213 3.4105
R2333 vdd.n1237 vdd.n1236 3.4105
R2334 vdd.n1245 vdd.n1244 3.4105
R2335 vdd.n1259 vdd.n307 3.4105
R2336 vdd.n1264 vdd.n301 3.4105
R2337 vdd.n1271 vdd.n1270 3.4105
R2338 vdd.n1287 vdd.n1286 3.4105
R2339 vdd.n1297 vdd.n1296 3.4105
R2340 vdd.n1311 vdd.n278 3.4105
R2341 vdd.n1170 vdd.n1169 3.4105
R2342 vdd.n1205 vdd.n1204 3.4105
R2343 vdd.n1101 vdd.n1100 3.4105
R2344 vdd.n1076 vdd.n393 3.4105
R2345 vdd.n1126 vdd.n1125 3.4105
R2346 vdd.n1108 vdd.n1107 3.4105
R2347 vdd.n1148 vdd.n1147 3.4105
R2348 vdd.n1133 vdd.n1132 3.4105
R2349 vdd.n1160 vdd.n1159 3.4105
R2350 vdd.n1155 vdd.n1154 3.4105
R2351 vdd.n1167 vdd.n1164 3.4105
R2352 vdd.n1181 vdd.n1180 3.4105
R2353 vdd.n1083 vdd.n1082 3.4105
R2354 vdd.n1072 vdd.n1071 3.4105
R2355 vdd.n967 vdd.n966 3.4105
R2356 vdd.n963 vdd.n962 3.4105
R2357 vdd.n986 vdd.n985 3.4105
R2358 vdd.n994 vdd.n993 3.4105
R2359 vdd.n1008 vdd.n441 3.4105
R2360 vdd.n1013 vdd.n435 3.4105
R2361 vdd.n1020 vdd.n1019 3.4105
R2362 vdd.n1036 vdd.n1035 3.4105
R2363 vdd.n1046 vdd.n1045 3.4105
R2364 vdd.n1060 vdd.n412 3.4105
R2365 vdd.n919 vdd.n918 3.4105
R2366 vdd.n954 vdd.n953 3.4105
R2367 vdd.n850 vdd.n849 3.4105
R2368 vdd.n825 vdd.n527 3.4105
R2369 vdd.n875 vdd.n874 3.4105
R2370 vdd.n857 vdd.n856 3.4105
R2371 vdd.n897 vdd.n896 3.4105
R2372 vdd.n882 vdd.n881 3.4105
R2373 vdd.n909 vdd.n908 3.4105
R2374 vdd.n904 vdd.n903 3.4105
R2375 vdd.n916 vdd.n913 3.4105
R2376 vdd.n930 vdd.n929 3.4105
R2377 vdd.n832 vdd.n831 3.4105
R2378 vdd.n821 vdd.n820 3.4105
R2379 vdd.n735 vdd.n734 3.4105
R2380 vdd.n743 vdd.n742 3.4105
R2381 vdd.n757 vdd.n575 3.4105
R2382 vdd.n762 vdd.n569 3.4105
R2383 vdd.n769 vdd.n768 3.4105
R2384 vdd.n785 vdd.n784 3.4105
R2385 vdd.n795 vdd.n794 3.4105
R2386 vdd.n809 vdd.n546 3.4105
R2387 vdd.n712 vdd.n711 3.4105
R2388 vdd.n716 vdd.n715 3.4105
R2389 vdd.n1689 vdd.n1688 3.4105
R2390 vdd.n1696 vdd.n1695 3.4105
R2391 vdd.n1719 vdd.n1718 3.4105
R2392 vdd.n44 vdd.n40 3.4105
R2393 vdd.n55 vdd.n43 3.4105
R2394 vdd.n1753 vdd.n1752 3.4105
R2395 vdd.n1746 vdd.n34 3.4105
R2396 vdd.n1776 vdd.n1775 3.4105
R2397 vdd.n1769 vdd.n1768 3.4105
R2398 vdd.n1863 vdd.n1862 3.4105
R2399 vdd.n1854 vdd.n1853 3.4105
R2400 vdd.n1711 vdd.n1710 3.4105
R2401 vdd.n1865 vdd.n1864 3.4105
R2402 vdd.n1858 vdd.n4 3.4105
R2403 vdd.n8 vdd.n7 3.4105
R2404 vdd.n1857 vdd.n6 3.4105
R2405 vdd.n1861 vdd.n1860 3.4105
R2406 vdd.n1774 vdd.n1773 3.4105
R2407 vdd.n24 vdd.n23 3.4105
R2408 vdd.n1772 vdd.n22 3.4105
R2409 vdd.n1745 vdd.n39 3.4105
R2410 vdd.n1749 vdd.n38 3.4105
R2411 vdd.n1751 vdd.n1750 3.4105
R2412 vdd.n1744 vdd.n1743 3.4105
R2413 vdd.n1715 vdd.n56 3.4105
R2414 vdd.n1742 vdd.n1741 3.4105
R2415 vdd.n58 vdd.n57 3.4105
R2416 vdd.n1714 vdd.n54 3.4105
R2417 vdd.n1717 vdd.n1716 3.4105
R2418 vdd.n1694 vdd.n1693 3.4105
R2419 vdd.n1692 vdd.n70 3.4105
R2420 vdd.n1661 vdd.n86 3.4105
R2421 vdd.n72 vdd.n71 3.4105
R2422 vdd.n1663 vdd.n1662 3.4105
R2423 vdd.n88 vdd.n87 3.4105
R2424 vdd.n1657 vdd.n85 3.4105
R2425 vdd.n1630 vdd.n103 3.4105
R2426 vdd.n1634 vdd.n102 3.4105
R2427 vdd.n1636 vdd.n1635 3.4105
R2428 vdd.n1629 vdd.n1628 3.4105
R2429 vdd.n1600 vdd.n120 3.4105
R2430 vdd.n1627 vdd.n1626 3.4105
R2431 vdd.n122 vdd.n121 3.4105
R2432 vdd.n1599 vdd.n118 3.4105
R2433 vdd.n1602 vdd.n1601 3.4105
R2434 vdd.n1579 vdd.n1578 3.4105
R2435 vdd.n136 vdd.n135 3.4105
R2436 vdd.n1577 vdd.n134 3.4105
R2437 vdd.n1541 vdd.n154 3.4105
R2438 vdd.n1546 vdd.n1545 3.4105
R2439 vdd.n1543 vdd.n1542 3.4105
R2440 vdd.n1540 vdd.n1539 3.4105
R2441 vdd.n1518 vdd.n171 3.4105
R2442 vdd.n1520 vdd.n1519 3.4105
R2443 vdd.n1492 vdd.n185 3.4105
R2444 vdd.n1513 vdd.n174 3.4105
R2445 vdd.n1517 vdd.n1516 3.4105
R2446 vdd.n1494 vdd.n1493 3.4105
R2447 vdd.n187 vdd.n186 3.4105
R2448 vdd.n1490 vdd.n1489 3.4105
R2449 vdd.n1459 vdd.n200 3.4105
R2450 vdd.n1467 vdd.n1460 3.4105
R2451 vdd.n1463 vdd.n1462 3.4105
R2452 vdd.n1458 vdd.n1457 3.4105
R2453 vdd.n1425 vdd.n1424 3.4105
R2454 vdd.n1423 vdd.n1422 3.4105
R2455 vdd.n1414 vdd.n219 3.4105
R2456 vdd.n1428 vdd.n220 3.4105
R2457 vdd.n1427 vdd.n1426 3.4105
R2458 vdd.n1413 vdd.n1412 3.4105
R2459 vdd.n1402 vdd.n226 3.4105
R2460 vdd.n222 vdd.n221 3.4105
R2461 vdd.n1380 vdd.n239 3.4105
R2462 vdd.n228 vdd.n227 3.4105
R2463 vdd.n1401 vdd.n1400 3.4105
R2464 vdd.n1379 vdd.n1378 3.4105
R2465 vdd.n1355 vdd.n254 3.4105
R2466 vdd.n241 vdd.n240 3.4105
R2467 vdd.n1330 vdd.n268 3.4105
R2468 vdd.n256 vdd.n255 3.4105
R2469 vdd.n1354 vdd.n1353 3.4105
R2470 vdd.n1332 vdd.n1331 3.4105
R2471 vdd.n270 vdd.n269 3.4105
R2472 vdd.n1326 vdd.n267 3.4105
R2473 vdd.n1290 vdd.n288 3.4105
R2474 vdd.n1295 vdd.n1294 3.4105
R2475 vdd.n1292 vdd.n1291 3.4105
R2476 vdd.n1289 vdd.n1288 3.4105
R2477 vdd.n1267 vdd.n305 3.4105
R2478 vdd.n1269 vdd.n1268 3.4105
R2479 vdd.n1241 vdd.n319 3.4105
R2480 vdd.n1262 vdd.n308 3.4105
R2481 vdd.n1266 vdd.n1265 3.4105
R2482 vdd.n1243 vdd.n1242 3.4105
R2483 vdd.n321 vdd.n320 3.4105
R2484 vdd.n1239 vdd.n1238 3.4105
R2485 vdd.n1208 vdd.n334 3.4105
R2486 vdd.n1216 vdd.n1209 3.4105
R2487 vdd.n1212 vdd.n1211 3.4105
R2488 vdd.n1207 vdd.n1206 3.4105
R2489 vdd.n1174 vdd.n1173 3.4105
R2490 vdd.n1172 vdd.n1171 3.4105
R2491 vdd.n1163 vdd.n353 3.4105
R2492 vdd.n1177 vdd.n354 3.4105
R2493 vdd.n1176 vdd.n1175 3.4105
R2494 vdd.n1162 vdd.n1161 3.4105
R2495 vdd.n1151 vdd.n360 3.4105
R2496 vdd.n356 vdd.n355 3.4105
R2497 vdd.n1129 vdd.n373 3.4105
R2498 vdd.n362 vdd.n361 3.4105
R2499 vdd.n1150 vdd.n1149 3.4105
R2500 vdd.n1128 vdd.n1127 3.4105
R2501 vdd.n1104 vdd.n388 3.4105
R2502 vdd.n375 vdd.n374 3.4105
R2503 vdd.n1079 vdd.n402 3.4105
R2504 vdd.n390 vdd.n389 3.4105
R2505 vdd.n1103 vdd.n1102 3.4105
R2506 vdd.n1081 vdd.n1080 3.4105
R2507 vdd.n404 vdd.n403 3.4105
R2508 vdd.n1075 vdd.n401 3.4105
R2509 vdd.n1039 vdd.n422 3.4105
R2510 vdd.n1044 vdd.n1043 3.4105
R2511 vdd.n1041 vdd.n1040 3.4105
R2512 vdd.n1038 vdd.n1037 3.4105
R2513 vdd.n1016 vdd.n439 3.4105
R2514 vdd.n1018 vdd.n1017 3.4105
R2515 vdd.n990 vdd.n453 3.4105
R2516 vdd.n1011 vdd.n442 3.4105
R2517 vdd.n1015 vdd.n1014 3.4105
R2518 vdd.n992 vdd.n991 3.4105
R2519 vdd.n455 vdd.n454 3.4105
R2520 vdd.n988 vdd.n987 3.4105
R2521 vdd.n957 vdd.n468 3.4105
R2522 vdd.n965 vdd.n958 3.4105
R2523 vdd.n961 vdd.n960 3.4105
R2524 vdd.n956 vdd.n955 3.4105
R2525 vdd.n923 vdd.n922 3.4105
R2526 vdd.n921 vdd.n920 3.4105
R2527 vdd.n912 vdd.n487 3.4105
R2528 vdd.n926 vdd.n488 3.4105
R2529 vdd.n925 vdd.n924 3.4105
R2530 vdd.n911 vdd.n910 3.4105
R2531 vdd.n900 vdd.n494 3.4105
R2532 vdd.n490 vdd.n489 3.4105
R2533 vdd.n878 vdd.n507 3.4105
R2534 vdd.n496 vdd.n495 3.4105
R2535 vdd.n899 vdd.n898 3.4105
R2536 vdd.n877 vdd.n876 3.4105
R2537 vdd.n853 vdd.n522 3.4105
R2538 vdd.n509 vdd.n508 3.4105
R2539 vdd.n828 vdd.n536 3.4105
R2540 vdd.n524 vdd.n523 3.4105
R2541 vdd.n852 vdd.n851 3.4105
R2542 vdd.n830 vdd.n829 3.4105
R2543 vdd.n538 vdd.n537 3.4105
R2544 vdd.n824 vdd.n535 3.4105
R2545 vdd.n788 vdd.n556 3.4105
R2546 vdd.n793 vdd.n792 3.4105
R2547 vdd.n790 vdd.n789 3.4105
R2548 vdd.n787 vdd.n786 3.4105
R2549 vdd.n765 vdd.n573 3.4105
R2550 vdd.n767 vdd.n766 3.4105
R2551 vdd.n739 vdd.n587 3.4105
R2552 vdd.n760 vdd.n576 3.4105
R2553 vdd.n764 vdd.n763 3.4105
R2554 vdd.n741 vdd.n740 3.4105
R2555 vdd.n589 vdd.n588 3.4105
R2556 vdd.n737 vdd.n736 3.4105
R2557 vdd.n706 vdd.n602 3.4105
R2558 vdd.n714 vdd.n707 3.4105
R2559 vdd.n710 vdd.n709 3.4105
R2560 vdd.n705 vdd.n704 3.4105
R2561 vdd.n614 vdd.n613 3.4105
R2562 vdd.n655 vdd.n654 3.4105
R2563 vdd.n660 vdd.n659 3.4105
R2564 vdd.n687 vdd.n686 3.4105
R2565 vdd.n688 vdd.n687 3.4105
R2566 vdd.n684 vdd.n683 3.4105
R2567 vdd.n685 vdd.n684 3.4105
R2568 vdd.n681 vdd.n680 3.4105
R2569 vdd.n682 vdd.n681 3.4105
R2570 vdd.n678 vdd.n677 3.4105
R2571 vdd.n679 vdd.n678 3.4105
R2572 vdd.n662 vdd.n661 3.4105
R2573 vdd.n663 vdd.n662 3.4105
R2574 vdd.n691 vdd.n690 3.4105
R2575 vdd.n691 vdd.n617 3.4105
R2576 vdd.n2842 vdd.n2841 3.4105
R2577 vdd.n2850 vdd.n2849 3.4105
R2578 vdd.n2935 vdd.n2934 3.4105
R2579 vdd.n2954 vdd.n2381 3.4105
R2580 vdd.n2959 vdd.n2372 3.4105
R2581 vdd.n2993 vdd.n2361 3.4105
R2582 vdd.n3014 vdd.n3013 3.4105
R2583 vdd.n3038 vdd.n3037 3.4105
R2584 vdd.n3048 vdd.n3047 3.4105
R2585 vdd.n3161 vdd.n3160 3.4105
R2586 vdd.n3180 vdd.n2247 3.4105
R2587 vdd.n3185 vdd.n2238 3.4105
R2588 vdd.n3219 vdd.n2227 3.4105
R2589 vdd.n3240 vdd.n3239 3.4105
R2590 vdd.n3264 vdd.n3263 3.4105
R2591 vdd.n3274 vdd.n3273 3.4105
R2592 vdd.n3387 vdd.n3386 3.4105
R2593 vdd.n3406 vdd.n2113 3.4105
R2594 vdd.n3411 vdd.n2104 3.4105
R2595 vdd.n3445 vdd.n2093 3.4105
R2596 vdd.n3466 vdd.n3465 3.4105
R2597 vdd.n3490 vdd.n3489 3.4105
R2598 vdd.n3500 vdd.n3499 3.4105
R2599 vdd.n3613 vdd.n3612 3.4105
R2600 vdd.n3632 vdd.n1979 3.4105
R2601 vdd.n3637 vdd.n1970 3.4105
R2602 vdd.n3671 vdd.n1959 3.4105
R2603 vdd.n3692 vdd.n3691 3.4105
R2604 vdd.n3696 vdd.n1940 3.4105
R2605 vdd.n3703 vdd.n3702 3.4105
R2606 vdd.n3678 vdd.n3677 3.4105
R2607 vdd.n1971 vdd.n1967 3.4105
R2608 vdd.n1981 vdd.n1977 3.4105
R2609 vdd.n3630 vdd.n3629 3.4105
R2610 vdd.n3586 vdd.n3585 3.4105
R2611 vdd.n3573 vdd.n3572 3.4105
R2612 vdd.n3566 vdd.n3565 3.4105
R2613 vdd.n3551 vdd.n3550 3.4105
R2614 vdd.n3544 vdd.n2039 3.4105
R2615 vdd.n3539 vdd.n2045 3.4105
R2616 vdd.n3528 vdd.n3527 3.4105
R2617 vdd.n3520 vdd.n3519 3.4105
R2618 vdd.n3593 vdd.n3592 3.4105
R2619 vdd.n3605 vdd.n3604 3.4105
R2620 vdd.n3507 vdd.n3506 3.4105
R2621 vdd.n3497 vdd.n3496 3.4105
R2622 vdd.n3473 vdd.n3472 3.4105
R2623 vdd.n3452 vdd.n3451 3.4105
R2624 vdd.n2105 vdd.n2101 3.4105
R2625 vdd.n2115 vdd.n2111 3.4105
R2626 vdd.n3404 vdd.n3403 3.4105
R2627 vdd.n3360 vdd.n3359 3.4105
R2628 vdd.n3347 vdd.n3346 3.4105
R2629 vdd.n3340 vdd.n3339 3.4105
R2630 vdd.n3325 vdd.n3324 3.4105
R2631 vdd.n3318 vdd.n2173 3.4105
R2632 vdd.n3313 vdd.n2179 3.4105
R2633 vdd.n3302 vdd.n3301 3.4105
R2634 vdd.n3294 vdd.n3293 3.4105
R2635 vdd.n3367 vdd.n3366 3.4105
R2636 vdd.n3379 vdd.n3378 3.4105
R2637 vdd.n3281 vdd.n3280 3.4105
R2638 vdd.n3271 vdd.n3270 3.4105
R2639 vdd.n3247 vdd.n3246 3.4105
R2640 vdd.n3226 vdd.n3225 3.4105
R2641 vdd.n2239 vdd.n2235 3.4105
R2642 vdd.n2249 vdd.n2245 3.4105
R2643 vdd.n3178 vdd.n3177 3.4105
R2644 vdd.n3134 vdd.n3133 3.4105
R2645 vdd.n3121 vdd.n3120 3.4105
R2646 vdd.n3114 vdd.n3113 3.4105
R2647 vdd.n3099 vdd.n3098 3.4105
R2648 vdd.n3092 vdd.n2307 3.4105
R2649 vdd.n3087 vdd.n2313 3.4105
R2650 vdd.n3076 vdd.n3075 3.4105
R2651 vdd.n3068 vdd.n3067 3.4105
R2652 vdd.n3141 vdd.n3140 3.4105
R2653 vdd.n3153 vdd.n3152 3.4105
R2654 vdd.n3055 vdd.n3054 3.4105
R2655 vdd.n3045 vdd.n3044 3.4105
R2656 vdd.n3021 vdd.n3020 3.4105
R2657 vdd.n3000 vdd.n2999 3.4105
R2658 vdd.n2373 vdd.n2369 3.4105
R2659 vdd.n2383 vdd.n2379 3.4105
R2660 vdd.n2952 vdd.n2951 3.4105
R2661 vdd.n2908 vdd.n2907 3.4105
R2662 vdd.n2895 vdd.n2894 3.4105
R2663 vdd.n2888 vdd.n2887 3.4105
R2664 vdd.n2873 vdd.n2872 3.4105
R2665 vdd.n2866 vdd.n2441 3.4105
R2666 vdd.n2861 vdd.n2447 3.4105
R2667 vdd.n2915 vdd.n2914 3.4105
R2668 vdd.n2927 vdd.n2926 3.4105
R2669 vdd.n2829 vdd.n2828 3.4105
R2670 vdd.n3828 vdd.n3827 3.4105
R2671 vdd.n3724 vdd.n3723 3.4105
R2672 vdd.n3731 vdd.n3730 3.4105
R2673 vdd.n3807 vdd.n3806 3.4105
R2674 vdd.n3800 vdd.n3799 3.4105
R2675 vdd.n3788 vdd.n3787 3.4105
R2676 vdd.n3781 vdd.n3780 3.4105
R2677 vdd.n3769 vdd.n3768 3.4105
R2678 vdd.n3762 vdd.n3761 3.4105
R2679 vdd.n3750 vdd.n3749 3.4105
R2680 vdd.n3743 vdd.n3742 3.4105
R2681 vdd.n3819 vdd.n3818 3.4105
R2682 vdd.n3830 vdd.n3829 3.4105
R2683 vdd.n3823 vdd.n1874 3.4105
R2684 vdd.n3826 vdd.n3825 3.4105
R2685 vdd.n1878 vdd.n1877 3.4105
R2686 vdd.n1893 vdd.n1892 3.4105
R2687 vdd.n3803 vdd.n1891 3.4105
R2688 vdd.n3805 vdd.n3804 3.4105
R2689 vdd.n3786 vdd.n3785 3.4105
R2690 vdd.n1904 vdd.n1903 3.4105
R2691 vdd.n3784 vdd.n1902 3.4105
R2692 vdd.n1915 vdd.n1914 3.4105
R2693 vdd.n3765 vdd.n1913 3.4105
R2694 vdd.n3767 vdd.n3766 3.4105
R2695 vdd.n3748 vdd.n3747 3.4105
R2696 vdd.n1926 vdd.n1925 3.4105
R2697 vdd.n3746 vdd.n1924 3.4105
R2698 vdd.n3727 vdd.n1935 3.4105
R2699 vdd.n3729 vdd.n3728 3.4105
R2700 vdd.n3822 vdd.n1876 3.4105
R2701 vdd.n2824 vdd.n2823 3.4105
R2702 vdd.n2827 vdd.n2826 3.4105
R2703 vdd.n2848 vdd.n2847 3.4105
R2704 vdd.n3699 vdd.n1948 3.4105
R2705 vdd.n1937 vdd.n1936 3.4105
R2706 vdd.n3701 vdd.n3700 3.4105
R2707 vdd.n1950 vdd.n1949 3.4105
R2708 vdd.n3695 vdd.n1947 3.4105
R2709 vdd.n3676 vdd.n3675 3.4105
R2710 vdd.n3670 vdd.n1966 3.4105
R2711 vdd.n3674 vdd.n1965 3.4105
R2712 vdd.n3669 vdd.n3668 3.4105
R2713 vdd.n3638 vdd.n3636 3.4105
R2714 vdd.n3667 vdd.n3666 3.4105
R2715 vdd.n3640 vdd.n3639 3.4105
R2716 vdd.n3634 vdd.n3633 3.4105
R2717 vdd.n3642 vdd.n3641 3.4105
R2718 vdd.n3631 vdd.n1982 3.4105
R2719 vdd.n3608 vdd.n1996 3.4105
R2720 vdd.n3609 vdd.n1983 3.4105
R2721 vdd.n3526 vdd.n3525 3.4105
R2722 vdd.n2057 vdd.n2056 3.4105
R2723 vdd.n3522 vdd.n3521 3.4105
R2724 vdd.n3546 vdd.n3545 3.4105
R2725 vdd.n3524 vdd.n2055 3.4105
R2726 vdd.n3542 vdd.n2046 3.4105
R2727 vdd.n3568 vdd.n3567 3.4105
R2728 vdd.n3547 vdd.n2043 3.4105
R2729 vdd.n3549 vdd.n3548 3.4105
R2730 vdd.n3588 vdd.n3587 3.4105
R2731 vdd.n3569 vdd.n2029 3.4105
R2732 vdd.n3571 vdd.n3570 3.4105
R2733 vdd.n3607 vdd.n3606 3.4105
R2734 vdd.n3589 vdd.n2018 3.4105
R2735 vdd.n3591 vdd.n3590 3.4105
R2736 vdd.n3505 vdd.n3504 3.4105
R2737 vdd.n2067 vdd.n2066 3.4105
R2738 vdd.n3502 vdd.n3501 3.4105
R2739 vdd.n3495 vdd.n3494 3.4105
R2740 vdd.n2071 vdd.n2070 3.4105
R2741 vdd.n3493 vdd.n2069 3.4105
R2742 vdd.n3471 vdd.n3470 3.4105
R2743 vdd.n2084 vdd.n2083 3.4105
R2744 vdd.n3469 vdd.n2082 3.4105
R2745 vdd.n3450 vdd.n3449 3.4105
R2746 vdd.n3444 vdd.n2100 3.4105
R2747 vdd.n3448 vdd.n2099 3.4105
R2748 vdd.n3443 vdd.n3442 3.4105
R2749 vdd.n3412 vdd.n3410 3.4105
R2750 vdd.n3441 vdd.n3440 3.4105
R2751 vdd.n3414 vdd.n3413 3.4105
R2752 vdd.n3408 vdd.n3407 3.4105
R2753 vdd.n3416 vdd.n3415 3.4105
R2754 vdd.n3405 vdd.n2116 3.4105
R2755 vdd.n3382 vdd.n2130 3.4105
R2756 vdd.n3383 vdd.n2117 3.4105
R2757 vdd.n3300 vdd.n3299 3.4105
R2758 vdd.n2191 vdd.n2190 3.4105
R2759 vdd.n3296 vdd.n3295 3.4105
R2760 vdd.n3320 vdd.n3319 3.4105
R2761 vdd.n3298 vdd.n2189 3.4105
R2762 vdd.n3316 vdd.n2180 3.4105
R2763 vdd.n3342 vdd.n3341 3.4105
R2764 vdd.n3321 vdd.n2177 3.4105
R2765 vdd.n3323 vdd.n3322 3.4105
R2766 vdd.n3362 vdd.n3361 3.4105
R2767 vdd.n3343 vdd.n2163 3.4105
R2768 vdd.n3345 vdd.n3344 3.4105
R2769 vdd.n3381 vdd.n3380 3.4105
R2770 vdd.n3363 vdd.n2152 3.4105
R2771 vdd.n3365 vdd.n3364 3.4105
R2772 vdd.n3279 vdd.n3278 3.4105
R2773 vdd.n2201 vdd.n2200 3.4105
R2774 vdd.n3276 vdd.n3275 3.4105
R2775 vdd.n3269 vdd.n3268 3.4105
R2776 vdd.n2205 vdd.n2204 3.4105
R2777 vdd.n3267 vdd.n2203 3.4105
R2778 vdd.n3245 vdd.n3244 3.4105
R2779 vdd.n2218 vdd.n2217 3.4105
R2780 vdd.n3243 vdd.n2216 3.4105
R2781 vdd.n3224 vdd.n3223 3.4105
R2782 vdd.n3218 vdd.n2234 3.4105
R2783 vdd.n3222 vdd.n2233 3.4105
R2784 vdd.n3217 vdd.n3216 3.4105
R2785 vdd.n3186 vdd.n3184 3.4105
R2786 vdd.n3215 vdd.n3214 3.4105
R2787 vdd.n3188 vdd.n3187 3.4105
R2788 vdd.n3182 vdd.n3181 3.4105
R2789 vdd.n3190 vdd.n3189 3.4105
R2790 vdd.n3179 vdd.n2250 3.4105
R2791 vdd.n3156 vdd.n2264 3.4105
R2792 vdd.n3157 vdd.n2251 3.4105
R2793 vdd.n3074 vdd.n3073 3.4105
R2794 vdd.n2325 vdd.n2324 3.4105
R2795 vdd.n3070 vdd.n3069 3.4105
R2796 vdd.n3094 vdd.n3093 3.4105
R2797 vdd.n3072 vdd.n2323 3.4105
R2798 vdd.n3090 vdd.n2314 3.4105
R2799 vdd.n3116 vdd.n3115 3.4105
R2800 vdd.n3095 vdd.n2311 3.4105
R2801 vdd.n3097 vdd.n3096 3.4105
R2802 vdd.n3136 vdd.n3135 3.4105
R2803 vdd.n3117 vdd.n2297 3.4105
R2804 vdd.n3119 vdd.n3118 3.4105
R2805 vdd.n3155 vdd.n3154 3.4105
R2806 vdd.n3137 vdd.n2286 3.4105
R2807 vdd.n3139 vdd.n3138 3.4105
R2808 vdd.n3053 vdd.n3052 3.4105
R2809 vdd.n2335 vdd.n2334 3.4105
R2810 vdd.n3050 vdd.n3049 3.4105
R2811 vdd.n3043 vdd.n3042 3.4105
R2812 vdd.n2339 vdd.n2338 3.4105
R2813 vdd.n3041 vdd.n2337 3.4105
R2814 vdd.n3019 vdd.n3018 3.4105
R2815 vdd.n2352 vdd.n2351 3.4105
R2816 vdd.n3017 vdd.n2350 3.4105
R2817 vdd.n2998 vdd.n2997 3.4105
R2818 vdd.n2992 vdd.n2368 3.4105
R2819 vdd.n2996 vdd.n2367 3.4105
R2820 vdd.n2991 vdd.n2990 3.4105
R2821 vdd.n2960 vdd.n2958 3.4105
R2822 vdd.n2989 vdd.n2988 3.4105
R2823 vdd.n2962 vdd.n2961 3.4105
R2824 vdd.n2956 vdd.n2955 3.4105
R2825 vdd.n2964 vdd.n2963 3.4105
R2826 vdd.n2953 vdd.n2384 3.4105
R2827 vdd.n2930 vdd.n2398 3.4105
R2828 vdd.n2931 vdd.n2385 3.4105
R2829 vdd.n2868 vdd.n2867 3.4105
R2830 vdd.n2846 vdd.n2457 3.4105
R2831 vdd.n2864 vdd.n2448 3.4105
R2832 vdd.n2890 vdd.n2889 3.4105
R2833 vdd.n2869 vdd.n2445 3.4105
R2834 vdd.n2871 vdd.n2870 3.4105
R2835 vdd.n2910 vdd.n2909 3.4105
R2836 vdd.n2891 vdd.n2431 3.4105
R2837 vdd.n2893 vdd.n2892 3.4105
R2838 vdd.n2929 vdd.n2928 3.4105
R2839 vdd.n2911 vdd.n2420 3.4105
R2840 vdd.n2913 vdd.n2912 3.4105
R2841 vdd.n2844 vdd.n2843 3.4105
R2842 vdd.n2459 vdd.n2458 3.4105
R2843 vdd.n2734 vdd.n2733 3.4105
R2844 vdd.n2739 vdd.n2738 3.4105
R2845 vdd.n2499 vdd.n2498 3.4105
R2846 vdd.n2500 vdd.n2499 3.4105
R2847 vdd.n2503 vdd.n2502 3.4105
R2848 vdd.n2503 vdd.n2466 3.4105
R2849 vdd.n2819 vdd.n2818 3.4105
R2850 vdd.n2818 vdd.n2469 3.4105
R2851 vdd.n2750 vdd.n2749 3.4105
R2852 vdd.n2750 vdd.n2747 3.4105
R2853 vdd.n2746 vdd.n2745 3.4105
R2854 vdd.n2745 vdd.n2740 3.4105
R2855 vdd.n2764 vdd.n1871 3.4105
R2856 vdd.n2784 vdd.n2783 3.4105
R2857 vdd.n2786 vdd.n2785 3.4105
R2858 vdd.n2768 vdd.n2767 3.4105
R2859 vdd.n2802 vdd.n2801 3.4105
R2860 vdd.n3622 vdd.n3619 3.38568
R2861 vdd.n3655 vdd.n1956 3.38568
R2862 vdd.n3396 vdd.n3393 3.38568
R2863 vdd.n3429 vdd.n2090 3.38568
R2864 vdd.n3486 vdd.n3480 3.38568
R2865 vdd.n3170 vdd.n3167 3.38568
R2866 vdd.n3203 vdd.n2224 3.38568
R2867 vdd.n3260 vdd.n3254 3.38568
R2868 vdd.n2944 vdd.n2941 3.38568
R2869 vdd.n2977 vdd.n2358 3.38568
R2870 vdd.n3034 vdd.n3028 3.38568
R2871 vdd.n3815 vdd.n3814 3.38568
R2872 vdd.n3582 vdd.n2013 3.38568
R2873 vdd.n3356 vdd.n2147 3.38568
R2874 vdd.n3130 vdd.n2281 3.38568
R2875 vdd.n2904 vdd.n2415 3.38568
R2876 vdd.n2599 vdd.n2592 3.30768
R2877 vdd.n2720 vdd.n2521 3.25021
R2878 vdd.n2619 vdd.n2568 3.24643
R2879 vdd.n2653 vdd.n2652 3.14007
R2880 vdd.n676 vdd.n675 3.11175
R2881 vdd.n720 vdd.n597 3.10353
R2882 vdd.n721 vdd.n592 3.10353
R2883 vdd.n729 vdd.n728 3.10353
R2884 vdd.n746 vdd.n583 3.10353
R2885 vdd.n753 vdd.n579 3.10353
R2886 vdd.n752 vdd.n566 3.10353
R2887 vdd.n570 vdd.n567 3.10353
R2888 vdd.n781 vdd.n562 3.10353
R2889 vdd.n799 vdd.n552 3.10353
R2890 vdd.n800 vdd.n548 3.10353
R2891 vdd.n815 vdd.n542 3.10353
R2892 vdd.n817 vdd.n816 3.10353
R2893 vdd.n839 vdd.n838 3.10353
R2894 vdd.n837 vdd.n528 3.10353
R2895 vdd.n862 vdd.n516 3.10353
R2896 vdd.n861 vdd.n517 3.10353
R2897 vdd.n869 vdd.n868 3.10353
R2898 vdd.n870 vdd.n503 3.10353
R2899 vdd.n890 vdd.n499 3.10353
R2900 vdd.n892 vdd.n891 3.10353
R2901 vdd.n936 vdd.n935 3.10353
R2902 vdd.n934 vdd.n478 3.10353
R2903 vdd.n944 vdd.n943 3.10353
R2904 vdd.n950 vdd.n474 3.10353
R2905 vdd.n971 vdd.n463 3.10353
R2906 vdd.n972 vdd.n458 3.10353
R2907 vdd.n980 vdd.n979 3.10353
R2908 vdd.n997 vdd.n449 3.10353
R2909 vdd.n1004 vdd.n445 3.10353
R2910 vdd.n1003 vdd.n432 3.10353
R2911 vdd.n436 vdd.n433 3.10353
R2912 vdd.n1032 vdd.n428 3.10353
R2913 vdd.n1050 vdd.n418 3.10353
R2914 vdd.n1051 vdd.n414 3.10353
R2915 vdd.n1066 vdd.n408 3.10353
R2916 vdd.n1068 vdd.n1067 3.10353
R2917 vdd.n1090 vdd.n1089 3.10353
R2918 vdd.n1088 vdd.n394 3.10353
R2919 vdd.n1113 vdd.n382 3.10353
R2920 vdd.n1112 vdd.n383 3.10353
R2921 vdd.n1120 vdd.n1119 3.10353
R2922 vdd.n1121 vdd.n369 3.10353
R2923 vdd.n1141 vdd.n365 3.10353
R2924 vdd.n1143 vdd.n1142 3.10353
R2925 vdd.n1187 vdd.n1186 3.10353
R2926 vdd.n1185 vdd.n344 3.10353
R2927 vdd.n1195 vdd.n1194 3.10353
R2928 vdd.n1201 vdd.n340 3.10353
R2929 vdd.n1222 vdd.n329 3.10353
R2930 vdd.n1223 vdd.n324 3.10353
R2931 vdd.n1231 vdd.n1230 3.10353
R2932 vdd.n1248 vdd.n315 3.10353
R2933 vdd.n1255 vdd.n311 3.10353
R2934 vdd.n1254 vdd.n298 3.10353
R2935 vdd.n302 vdd.n299 3.10353
R2936 vdd.n1283 vdd.n294 3.10353
R2937 vdd.n1301 vdd.n284 3.10353
R2938 vdd.n1302 vdd.n280 3.10353
R2939 vdd.n1317 vdd.n274 3.10353
R2940 vdd.n1319 vdd.n1318 3.10353
R2941 vdd.n1341 vdd.n1340 3.10353
R2942 vdd.n1339 vdd.n260 3.10353
R2943 vdd.n1364 vdd.n248 3.10353
R2944 vdd.n1363 vdd.n249 3.10353
R2945 vdd.n1371 vdd.n1370 3.10353
R2946 vdd.n1372 vdd.n235 3.10353
R2947 vdd.n1392 vdd.n231 3.10353
R2948 vdd.n1394 vdd.n1393 3.10353
R2949 vdd.n1438 vdd.n1437 3.10353
R2950 vdd.n1436 vdd.n210 3.10353
R2951 vdd.n1446 vdd.n1445 3.10353
R2952 vdd.n1452 vdd.n206 3.10353
R2953 vdd.n1473 vdd.n195 3.10353
R2954 vdd.n1474 vdd.n190 3.10353
R2955 vdd.n1482 vdd.n1481 3.10353
R2956 vdd.n1499 vdd.n181 3.10353
R2957 vdd.n1506 vdd.n177 3.10353
R2958 vdd.n1505 vdd.n164 3.10353
R2959 vdd.n168 vdd.n165 3.10353
R2960 vdd.n1534 vdd.n160 3.10353
R2961 vdd.n1552 vdd.n150 3.10353
R2962 vdd.n1553 vdd.n146 3.10353
R2963 vdd.n1568 vdd.n140 3.10353
R2964 vdd.n1570 vdd.n1569 3.10353
R2965 vdd.n1587 vdd.n1586 3.10353
R2966 vdd.n1585 vdd.n127 3.10353
R2967 vdd.n1610 vdd.n114 3.10353
R2968 vdd.n1609 vdd.n115 3.10353
R2969 vdd.n1617 vdd.n1616 3.10353
R2970 vdd.n1618 vdd.n96 3.10353
R2971 vdd.n1648 vdd.n92 3.10353
R2972 vdd.n1650 vdd.n1649 3.10353
R2973 vdd.n1672 vdd.n1671 3.10353
R2974 vdd.n1670 vdd.n76 3.10353
R2975 vdd.n1702 vdd.n1701 3.10353
R2976 vdd.n1700 vdd.n63 3.10353
R2977 vdd.n1725 vdd.n50 3.10353
R2978 vdd.n1724 vdd.n51 3.10353
R2979 vdd.n1732 vdd.n1731 3.10353
R2980 vdd.n1733 vdd.n32 3.10353
R2981 vdd.n1763 vdd.n28 3.10353
R2982 vdd.n1765 vdd.n1764 3.10353
R2983 vdd.n1782 vdd.n1781 3.10353
R2984 vdd.n1780 vdd.n13 3.10353
R2985 vdd.n2836 vdd.n2462 3.10353
R2986 vdd.n2835 vdd.n2453 3.10353
R2987 vdd.n2857 vdd.n2451 3.10353
R2988 vdd.n2856 vdd.n2438 3.10353
R2989 vdd.n2442 vdd.n2439 3.10353
R2990 vdd.n2884 vdd.n2436 3.10353
R2991 vdd.n2899 vdd.n2427 3.10353
R2992 vdd.n2900 vdd.n2425 3.10353
R2993 vdd.n2919 vdd.n2416 3.10353
R2994 vdd.n2920 vdd.n2405 3.10353
R2995 vdd.n2414 vdd.n2413 3.10353
R2996 vdd.n2406 vdd.n2394 3.10353
R2997 vdd.n2393 vdd.n2390 3.10353
R2998 vdd.n2947 vdd.n2946 3.10353
R2999 vdd.n2392 vdd.n2391 3.10353
R3000 vdd.n2972 vdd.n2377 3.10353
R3001 vdd.n2979 vdd.n2375 3.10353
R3002 vdd.n2980 vdd.n2359 3.10353
R3003 vdd.n3005 vdd.n2357 3.10353
R3004 vdd.n2362 vdd.n2356 3.10353
R3005 vdd.n3026 vdd.n2347 3.10353
R3006 vdd.n3025 vdd.n2344 3.10353
R3007 vdd.n3031 vdd.n2345 3.10353
R3008 vdd.n3030 vdd.n2330 3.10353
R3009 vdd.n3062 vdd.n2328 3.10353
R3010 vdd.n3061 vdd.n2319 3.10353
R3011 vdd.n3083 vdd.n2317 3.10353
R3012 vdd.n3082 vdd.n2304 3.10353
R3013 vdd.n2308 vdd.n2305 3.10353
R3014 vdd.n3110 vdd.n2302 3.10353
R3015 vdd.n3125 vdd.n2293 3.10353
R3016 vdd.n3126 vdd.n2291 3.10353
R3017 vdd.n3145 vdd.n2282 3.10353
R3018 vdd.n3146 vdd.n2271 3.10353
R3019 vdd.n2280 vdd.n2279 3.10353
R3020 vdd.n2272 vdd.n2260 3.10353
R3021 vdd.n2259 vdd.n2256 3.10353
R3022 vdd.n3173 vdd.n3172 3.10353
R3023 vdd.n2258 vdd.n2257 3.10353
R3024 vdd.n3198 vdd.n2243 3.10353
R3025 vdd.n3205 vdd.n2241 3.10353
R3026 vdd.n3206 vdd.n2225 3.10353
R3027 vdd.n3231 vdd.n2223 3.10353
R3028 vdd.n2228 vdd.n2222 3.10353
R3029 vdd.n3252 vdd.n2213 3.10353
R3030 vdd.n3251 vdd.n2210 3.10353
R3031 vdd.n3257 vdd.n2211 3.10353
R3032 vdd.n3256 vdd.n2196 3.10353
R3033 vdd.n3288 vdd.n2194 3.10353
R3034 vdd.n3287 vdd.n2185 3.10353
R3035 vdd.n3309 vdd.n2183 3.10353
R3036 vdd.n3308 vdd.n2170 3.10353
R3037 vdd.n2174 vdd.n2171 3.10353
R3038 vdd.n3336 vdd.n2168 3.10353
R3039 vdd.n3351 vdd.n2159 3.10353
R3040 vdd.n3352 vdd.n2157 3.10353
R3041 vdd.n3371 vdd.n2148 3.10353
R3042 vdd.n3372 vdd.n2137 3.10353
R3043 vdd.n2146 vdd.n2145 3.10353
R3044 vdd.n2138 vdd.n2126 3.10353
R3045 vdd.n2125 vdd.n2122 3.10353
R3046 vdd.n3399 vdd.n3398 3.10353
R3047 vdd.n2124 vdd.n2123 3.10353
R3048 vdd.n3424 vdd.n2109 3.10353
R3049 vdd.n3431 vdd.n2107 3.10353
R3050 vdd.n3432 vdd.n2091 3.10353
R3051 vdd.n3457 vdd.n2089 3.10353
R3052 vdd.n2094 vdd.n2088 3.10353
R3053 vdd.n3478 vdd.n2079 3.10353
R3054 vdd.n3477 vdd.n2076 3.10353
R3055 vdd.n3483 vdd.n2077 3.10353
R3056 vdd.n3482 vdd.n2062 3.10353
R3057 vdd.n3514 vdd.n2060 3.10353
R3058 vdd.n3513 vdd.n2051 3.10353
R3059 vdd.n3535 vdd.n2049 3.10353
R3060 vdd.n3534 vdd.n2036 3.10353
R3061 vdd.n2040 vdd.n2037 3.10353
R3062 vdd.n3562 vdd.n2034 3.10353
R3063 vdd.n3577 vdd.n2025 3.10353
R3064 vdd.n3578 vdd.n2023 3.10353
R3065 vdd.n3597 vdd.n2014 3.10353
R3066 vdd.n3598 vdd.n2003 3.10353
R3067 vdd.n2012 vdd.n2011 3.10353
R3068 vdd.n2004 vdd.n1992 3.10353
R3069 vdd.n1991 vdd.n1988 3.10353
R3070 vdd.n3625 vdd.n3624 3.10353
R3071 vdd.n1990 vdd.n1989 3.10353
R3072 vdd.n3650 vdd.n1975 3.10353
R3073 vdd.n3657 vdd.n1973 3.10353
R3074 vdd.n3658 vdd.n1957 3.10353
R3075 vdd.n3683 vdd.n1955 3.10353
R3076 vdd.n1960 vdd.n1954 3.10353
R3077 vdd.n3709 vdd.n1944 3.10353
R3078 vdd.n3708 vdd.n1941 3.10353
R3079 vdd.n3736 vdd.n1932 3.10353
R3080 vdd.n3735 vdd.n1930 3.10353
R3081 vdd.n3755 vdd.n1921 3.10353
R3082 vdd.n3754 vdd.n1919 3.10353
R3083 vdd.n3774 vdd.n1910 3.10353
R3084 vdd.n3773 vdd.n1908 3.10353
R3085 vdd.n3793 vdd.n1899 3.10353
R3086 vdd.n3792 vdd.n1897 3.10353
R3087 vdd.n3812 vdd.n1888 3.10353
R3088 vdd.n3811 vdd.n1883 3.10353
R3089 vdd.n1833 vdd.n1832 3.03311
R3090 vdd.n2760 vdd.n2758 3.03311
R3091 vdd.n2723 vdd.n2722 2.9318
R3092 vdd.n2491 vdd 2.90898
R3093 vdd.n2587 vdd.n2575 2.81772
R3094 vdd.n2603 vdd.n2575 2.81772
R3095 vdd.n2636 vdd.n2635 2.69524
R3096 vdd.n1824 vdd.n1823 2.64177
R3097 vdd.n2789 vdd.n2759 2.64177
R3098 vdd.n2634 vdd.n2633 2.63399
R3099 vdd.n2581 vdd 2.55084
R3100 vdd.n2646 vdd.t27 2.55084
R3101 vdd.n1686 vdd.n67 2.54483
R3102 vdd.n3722 vdd.n3721 2.54394
R3103 vdd.n2704 vdd.n2538 2.54096
R3104 vdd.n1832 vdd.n1822 2.4386
R3105 vdd.n2775 vdd.n2758 2.4386
R3106 vdd.n2592 vdd.n2577 2.32777
R3107 vdd.n2618 vdd.n2617 2.3255
R3108 vdd.n1845 vdd.n14 2.28608
R3109 vdd.n2482 vdd.n1884 2.28608
R3110 vdd vdd.n2820 2.28482
R3111 vdd.n694 vdd.n610 2.24869
R3112 vdd.n644 vdd.n643 2.24869
R3113 vdd.n637 vdd.n636 2.24869
R3114 vdd.n634 vdd.n632 2.24869
R3115 vdd.n622 vdd.n621 2.24869
R3116 vdd.n2753 vdd.n2509 2.24869
R3117 vdd.n2815 vdd.n2814 2.24869
R3118 vdd.n2506 vdd.n2471 2.24869
R3119 vdd.n2488 vdd.n2486 2.24869
R3120 vdd.n2493 vdd.n2492 2.24869
R3121 vdd.n2720 vdd.n2520 2.16698
R3122 vdd.n1845 vdd.n1844 2.15377
R3123 vdd.n2485 vdd.n2482 2.15377
R3124 vdd.n2616 vdd 2.13331
R3125 vdd.n2590 vdd 2.02977
R3126 vdd.n2490 vdd.n2489 1.99051
R3127 vdd.n1842 vdd.n3 1.94045
R3128 vdd.n1803 vdd.n1802 1.94045
R3129 vdd.n2483 vdd.n1873 1.94045
R3130 vdd.n2691 vdd.n2527 1.94045
R3131 vdd.n2699 vdd.n2698 1.94045
R3132 vdd.n2726 vdd.n2725 1.94045
R3133 vdd.n2658 vdd.n2657 1.94045
R3134 vdd.n2686 vdd.n2685 1.94045
R3135 vdd.n2798 vdd.n2797 1.94045
R3136 vdd.n2771 vdd.n2770 1.94045
R3137 vdd.n2708 vdd.n2532 1.85699
R3138 vdd.n2722 vdd.n2518 1.85699
R3139 vdd.n2718 vdd.n2524 1.85557
R3140 vdd.n1588 vdd.n130 1.76521
R3141 vdd.n1592 vdd.n113 1.76521
R3142 vdd.n1615 vdd.n111 1.76521
R3143 vdd.n1643 vdd.n93 1.76521
R3144 vdd.n1673 vdd.n81 1.76521
R3145 vdd.n1679 vdd.n79 1.76521
R3146 vdd.n1451 vdd.n194 1.76521
R3147 vdd.n1479 vdd.n192 1.76521
R3148 vdd.n1500 vdd.n178 1.76521
R3149 vdd.n1529 vdd.n163 1.76521
R3150 vdd.n1533 vdd.n149 1.76521
R3151 vdd.n1559 vdd.n147 1.76521
R3152 vdd.n1342 vdd.n263 1.76521
R3153 vdd.n1346 vdd.n247 1.76521
R3154 vdd.n1369 vdd.n245 1.76521
R3155 vdd.n1387 vdd.n232 1.76521
R3156 vdd.n1439 vdd.n214 1.76521
R3157 vdd.n1443 vdd.n209 1.76521
R3158 vdd.n1200 vdd.n328 1.76521
R3159 vdd.n1228 vdd.n326 1.76521
R3160 vdd.n1249 vdd.n312 1.76521
R3161 vdd.n1278 vdd.n297 1.76521
R3162 vdd.n1282 vdd.n283 1.76521
R3163 vdd.n1308 vdd.n281 1.76521
R3164 vdd.n1091 vdd.n397 1.76521
R3165 vdd.n1095 vdd.n381 1.76521
R3166 vdd.n1118 vdd.n379 1.76521
R3167 vdd.n1136 vdd.n366 1.76521
R3168 vdd.n1188 vdd.n348 1.76521
R3169 vdd.n1192 vdd.n343 1.76521
R3170 vdd.n949 vdd.n462 1.76521
R3171 vdd.n977 vdd.n460 1.76521
R3172 vdd.n998 vdd.n446 1.76521
R3173 vdd.n1027 vdd.n431 1.76521
R3174 vdd.n1031 vdd.n417 1.76521
R3175 vdd.n1057 vdd.n415 1.76521
R3176 vdd.n840 vdd.n531 1.76521
R3177 vdd.n844 vdd.n515 1.76521
R3178 vdd.n867 vdd.n513 1.76521
R3179 vdd.n885 vdd.n500 1.76521
R3180 vdd.n937 vdd.n482 1.76521
R3181 vdd.n941 vdd.n477 1.76521
R3182 vdd.n608 vdd.n596 1.76521
R3183 vdd.n726 vdd.n594 1.76521
R3184 vdd.n747 vdd.n580 1.76521
R3185 vdd.n776 vdd.n565 1.76521
R3186 vdd.n780 vdd.n551 1.76521
R3187 vdd.n806 vdd.n549 1.76521
R3188 vdd.n1703 vdd.n66 1.76521
R3189 vdd.n1707 vdd.n49 1.76521
R3190 vdd.n1730 vdd.n47 1.76521
R3191 vdd.n1758 vdd.n29 1.76521
R3192 vdd.n1783 vdd.n18 1.76521
R3193 vdd.n1850 vdd.n16 1.76521
R3194 vdd.n3622 vdd.n3621 1.76521
R3195 vdd.n3684 vdd.n1956 1.76521
R3196 vdd.n3510 vdd.n2061 1.76521
R3197 vdd.n3531 vdd.n2050 1.76521
R3198 vdd.n3558 vdd.n2035 1.76521
R3199 vdd.n3561 vdd.n2024 1.76521
R3200 vdd.n3582 vdd.n3581 1.76521
R3201 vdd.n3396 vdd.n3395 1.76521
R3202 vdd.n3458 vdd.n2090 1.76521
R3203 vdd.n3486 vdd.n3485 1.76521
R3204 vdd.n3284 vdd.n2195 1.76521
R3205 vdd.n3305 vdd.n2184 1.76521
R3206 vdd.n3332 vdd.n2169 1.76521
R3207 vdd.n3335 vdd.n2158 1.76521
R3208 vdd.n3356 vdd.n3355 1.76521
R3209 vdd.n3170 vdd.n3169 1.76521
R3210 vdd.n3232 vdd.n2224 1.76521
R3211 vdd.n3260 vdd.n3259 1.76521
R3212 vdd.n3058 vdd.n2329 1.76521
R3213 vdd.n3079 vdd.n2318 1.76521
R3214 vdd.n3106 vdd.n2303 1.76521
R3215 vdd.n3109 vdd.n2292 1.76521
R3216 vdd.n3130 vdd.n3129 1.76521
R3217 vdd.n2944 vdd.n2943 1.76521
R3218 vdd.n3006 vdd.n2358 1.76521
R3219 vdd.n3034 vdd.n3033 1.76521
R3220 vdd.n2880 vdd.n2437 1.76521
R3221 vdd.n2883 vdd.n2426 1.76521
R3222 vdd.n2904 vdd.n2903 1.76521
R3223 vdd.n3720 vdd.n3719 1.76521
R3224 vdd.n3815 vdd.n1885 1.76521
R3225 vdd.n2613 vdd.n2568 1.71533
R3226 vdd.n2497 vdd.n2496 1.706
R3227 vdd.n2491 vdd.t0 1.68435
R3228 vdd.n3738 vdd.n1920 1.66612
R3229 vdd.n3757 vdd.n1909 1.66612
R3230 vdd.n3776 vdd.n1898 1.66612
R3231 vdd.n3795 vdd.n1887 1.66612
R3232 vdd.n2939 vdd.n2938 1.66612
R3233 vdd.n2976 vdd.n2975 1.66612
R3234 vdd.n3009 vdd.n2346 1.66612
R3235 vdd.n3165 vdd.n3164 1.66612
R3236 vdd.n3202 vdd.n3201 1.66612
R3237 vdd.n3235 vdd.n2212 1.66612
R3238 vdd.n3391 vdd.n3390 1.66612
R3239 vdd.n3428 vdd.n3427 1.66612
R3240 vdd.n3461 vdd.n2078 1.66612
R3241 vdd.n3617 vdd.n3616 1.66612
R3242 vdd.n3654 vdd.n3653 1.66612
R3243 vdd.n3687 vdd.n1943 1.66612
R3244 vdd.n3601 vdd.n3600 1.66612
R3245 vdd.n3375 vdd.n3374 1.66612
R3246 vdd.n3149 vdd.n3148 1.66612
R3247 vdd.n2923 vdd.n2922 1.66612
R3248 vdd.n2833 vdd.n2452 1.66612
R3249 vdd.n2539 vdd.n2517 1.36844
R3250 vdd.n1820 vdd.n1819 1.35607
R3251 vdd.n702 vdd.n701 1.35607
R3252 vdd.n1595 vdd.n1594 1.35607
R3253 vdd.n109 vdd.n107 1.35607
R3254 vdd.n1641 vdd.n98 1.35607
R3255 vdd.n1653 vdd.n1652 1.35607
R3256 vdd.n1681 vdd.n75 1.35607
R3257 vdd.n1573 vdd.n1572 1.35607
R3258 vdd.n1465 vdd.n191 1.35607
R3259 vdd.n1497 vdd.n1496 1.35607
R3260 vdd.n1527 vdd.n167 1.35607
R3261 vdd.n1537 vdd.n1536 1.35607
R3262 vdd.n1562 vdd.n1561 1.35607
R3263 vdd.n1455 vdd.n1454 1.35607
R3264 vdd.n1348 vdd.n259 1.35607
R3265 vdd.n1359 vdd.n251 1.35607
R3266 vdd.n1385 vdd.n1384 1.35607
R3267 vdd.n1407 vdd.n1406 1.35607
R3268 vdd.n1432 vdd.n211 1.35607
R3269 vdd.n1322 vdd.n1321 1.35607
R3270 vdd.n1214 vdd.n325 1.35607
R3271 vdd.n1246 vdd.n1245 1.35607
R3272 vdd.n1276 vdd.n301 1.35607
R3273 vdd.n1286 vdd.n1285 1.35607
R3274 vdd.n1311 vdd.n1310 1.35607
R3275 vdd.n1204 vdd.n1203 1.35607
R3276 vdd.n1097 vdd.n393 1.35607
R3277 vdd.n1108 vdd.n385 1.35607
R3278 vdd.n1134 vdd.n1133 1.35607
R3279 vdd.n1156 vdd.n1155 1.35607
R3280 vdd.n1181 vdd.n345 1.35607
R3281 vdd.n1071 vdd.n1070 1.35607
R3282 vdd.n963 vdd.n459 1.35607
R3283 vdd.n995 vdd.n994 1.35607
R3284 vdd.n1025 vdd.n435 1.35607
R3285 vdd.n1035 vdd.n1034 1.35607
R3286 vdd.n1060 vdd.n1059 1.35607
R3287 vdd.n953 vdd.n952 1.35607
R3288 vdd.n846 vdd.n527 1.35607
R3289 vdd.n857 vdd.n519 1.35607
R3290 vdd.n883 vdd.n882 1.35607
R3291 vdd.n905 vdd.n904 1.35607
R3292 vdd.n930 vdd.n479 1.35607
R3293 vdd.n820 vdd.n819 1.35607
R3294 vdd.n744 vdd.n743 1.35607
R3295 vdd.n774 vdd.n569 1.35607
R3296 vdd.n784 vdd.n783 1.35607
R3297 vdd.n809 vdd.n808 1.35607
R3298 vdd.n712 vdd.n593 1.35607
R3299 vdd.n45 vdd.n43 1.35607
R3300 vdd.n1756 vdd.n34 1.35607
R3301 vdd.n1768 vdd.n1767 1.35607
R3302 vdd.n1853 vdd.n1852 1.35607
R3303 vdd.n1710 vdd.n1709 1.35607
R3304 vdd.n2851 vdd.n2850 1.35607
R3305 vdd.n2936 vdd.n2935 1.35607
R3306 vdd.n2381 vdd.n2380 1.35607
R3307 vdd.n2374 vdd.n2372 1.35607
R3308 vdd.n3003 vdd.n2361 1.35607
R3309 vdd.n3013 vdd.n3012 1.35607
R3310 vdd.n3037 vdd.n3036 1.35607
R3311 vdd.n3162 vdd.n3161 1.35607
R3312 vdd.n2247 vdd.n2246 1.35607
R3313 vdd.n2240 vdd.n2238 1.35607
R3314 vdd.n3229 vdd.n2227 1.35607
R3315 vdd.n3239 vdd.n3238 1.35607
R3316 vdd.n3263 vdd.n3262 1.35607
R3317 vdd.n3388 vdd.n3387 1.35607
R3318 vdd.n2113 vdd.n2112 1.35607
R3319 vdd.n2106 vdd.n2104 1.35607
R3320 vdd.n3455 vdd.n2093 1.35607
R3321 vdd.n3465 vdd.n3464 1.35607
R3322 vdd.n3489 vdd.n3488 1.35607
R3323 vdd.n3614 vdd.n3613 1.35607
R3324 vdd.n1979 vdd.n1978 1.35607
R3325 vdd.n1972 vdd.n1970 1.35607
R3326 vdd.n3681 vdd.n1959 1.35607
R3327 vdd.n3691 vdd.n3690 1.35607
R3328 vdd.n3713 vdd.n1940 1.35607
R3329 vdd.n3585 vdd.n3584 1.35607
R3330 vdd.n3565 vdd.n3564 1.35607
R3331 vdd.n3556 vdd.n2039 1.35607
R3332 vdd.n3529 vdd.n3528 1.35607
R3333 vdd.n3604 vdd.n3603 1.35607
R3334 vdd.n3508 vdd.n3507 1.35607
R3335 vdd.n3359 vdd.n3358 1.35607
R3336 vdd.n3339 vdd.n3338 1.35607
R3337 vdd.n3330 vdd.n2173 1.35607
R3338 vdd.n3303 vdd.n3302 1.35607
R3339 vdd.n3378 vdd.n3377 1.35607
R3340 vdd.n3282 vdd.n3281 1.35607
R3341 vdd.n3133 vdd.n3132 1.35607
R3342 vdd.n3113 vdd.n3112 1.35607
R3343 vdd.n3104 vdd.n2307 1.35607
R3344 vdd.n3077 vdd.n3076 1.35607
R3345 vdd.n3152 vdd.n3151 1.35607
R3346 vdd.n3056 vdd.n3055 1.35607
R3347 vdd.n2907 vdd.n2906 1.35607
R3348 vdd.n2887 vdd.n2886 1.35607
R3349 vdd.n2878 vdd.n2441 1.35607
R3350 vdd.n2926 vdd.n2925 1.35607
R3351 vdd.n2830 vdd.n2829 1.35607
R3352 vdd.n3799 vdd.n3798 1.35607
R3353 vdd.n3780 vdd.n3779 1.35607
R3354 vdd.n3761 vdd.n3760 1.35607
R3355 vdd.n3742 vdd.n3741 1.35607
R3356 vdd.n3818 vdd.n3817 1.35607
R3357 vdd.n2804 vdd.n2803 1.35607
R3358 vdd.n648 vdd.n647 1.13981
R3359 vdd.n2742 vdd.n2741 1.13981
R3360 vdd.n10 vdd.n6 1.13717
R3361 vdd.n26 vdd.n22 1.13717
R3362 vdd.n38 vdd.n36 1.13717
R3363 vdd.n1741 vdd.n1740 1.13717
R3364 vdd.n60 vdd.n54 1.13717
R3365 vdd.n1687 vdd.n70 1.13717
R3366 vdd.n1691 vdd.n1690 1.13717
R3367 vdd.n1713 vdd.n1712 1.13717
R3368 vdd.n42 vdd.n41 1.13717
R3369 vdd.n1748 vdd.n1747 1.13717
R3370 vdd.n1771 vdd.n1770 1.13717
R3371 vdd.n1856 vdd.n1855 1.13717
R3372 vdd.n73 vdd.n72 1.13717
R3373 vdd.n90 vdd.n85 1.13717
R3374 vdd.n102 vdd.n100 1.13717
R3375 vdd.n1626 vdd.n1625 1.13717
R3376 vdd.n124 vdd.n118 1.13717
R3377 vdd.n138 vdd.n134 1.13717
R3378 vdd.n1546 vdd.n143 1.13717
R3379 vdd.n1520 vdd.n158 1.13717
R3380 vdd.n1513 vdd.n1512 1.13717
R3381 vdd.n1489 vdd.n183 1.13717
R3382 vdd.n1467 vdd.n1466 1.13717
R3383 vdd.n1422 vdd.n204 1.13717
R3384 vdd.n220 vdd.n218 1.13717
R3385 vdd.n223 vdd.n222 1.13717
R3386 vdd.n238 vdd.n228 1.13717
R3387 vdd.n253 vdd.n241 1.13717
R3388 vdd.n257 vdd.n256 1.13717
R3389 vdd.n272 vdd.n267 1.13717
R3390 vdd.n1295 vdd.n277 1.13717
R3391 vdd.n1269 vdd.n292 1.13717
R3392 vdd.n1262 vdd.n1261 1.13717
R3393 vdd.n1238 vdd.n317 1.13717
R3394 vdd.n1216 vdd.n1215 1.13717
R3395 vdd.n1171 vdd.n338 1.13717
R3396 vdd.n354 vdd.n352 1.13717
R3397 vdd.n357 vdd.n356 1.13717
R3398 vdd.n372 vdd.n362 1.13717
R3399 vdd.n387 vdd.n375 1.13717
R3400 vdd.n391 vdd.n390 1.13717
R3401 vdd.n406 vdd.n401 1.13717
R3402 vdd.n1044 vdd.n411 1.13717
R3403 vdd.n1018 vdd.n426 1.13717
R3404 vdd.n1011 vdd.n1010 1.13717
R3405 vdd.n987 vdd.n451 1.13717
R3406 vdd.n965 vdd.n964 1.13717
R3407 vdd.n920 vdd.n472 1.13717
R3408 vdd.n488 vdd.n486 1.13717
R3409 vdd.n491 vdd.n490 1.13717
R3410 vdd.n506 vdd.n496 1.13717
R3411 vdd.n521 vdd.n509 1.13717
R3412 vdd.n525 vdd.n524 1.13717
R3413 vdd.n540 vdd.n535 1.13717
R3414 vdd.n793 vdd.n545 1.13717
R3415 vdd.n767 vdd.n560 1.13717
R3416 vdd.n760 vdd.n759 1.13717
R3417 vdd.n736 vdd.n585 1.13717
R3418 vdd.n714 vdd.n713 1.13717
R3419 vdd.n614 vdd.n606 1.13717
R3420 vdd.n605 vdd.n604 1.13717
R3421 vdd.n708 vdd.n603 1.13717
R3422 vdd.n738 vdd.n586 1.13717
R3423 vdd.n761 vdd.n574 1.13717
R3424 vdd.n559 vdd.n558 1.13717
R3425 vdd.n791 vdd.n557 1.13717
R3426 vdd.n823 vdd.n822 1.13717
R3427 vdd.n827 vdd.n826 1.13717
R3428 vdd.n855 vdd.n854 1.13717
R3429 vdd.n880 vdd.n879 1.13717
R3430 vdd.n902 vdd.n901 1.13717
R3431 vdd.n928 vdd.n927 1.13717
R3432 vdd.n471 vdd.n470 1.13717
R3433 vdd.n959 vdd.n469 1.13717
R3434 vdd.n989 vdd.n452 1.13717
R3435 vdd.n1012 vdd.n440 1.13717
R3436 vdd.n425 vdd.n424 1.13717
R3437 vdd.n1042 vdd.n423 1.13717
R3438 vdd.n1074 vdd.n1073 1.13717
R3439 vdd.n1078 vdd.n1077 1.13717
R3440 vdd.n1106 vdd.n1105 1.13717
R3441 vdd.n1131 vdd.n1130 1.13717
R3442 vdd.n1153 vdd.n1152 1.13717
R3443 vdd.n1179 vdd.n1178 1.13717
R3444 vdd.n337 vdd.n336 1.13717
R3445 vdd.n1210 vdd.n335 1.13717
R3446 vdd.n1240 vdd.n318 1.13717
R3447 vdd.n1263 vdd.n306 1.13717
R3448 vdd.n291 vdd.n290 1.13717
R3449 vdd.n1293 vdd.n289 1.13717
R3450 vdd.n1325 vdd.n1324 1.13717
R3451 vdd.n1329 vdd.n1328 1.13717
R3452 vdd.n1357 vdd.n1356 1.13717
R3453 vdd.n1382 vdd.n1381 1.13717
R3454 vdd.n1404 vdd.n1403 1.13717
R3455 vdd.n1430 vdd.n1429 1.13717
R3456 vdd.n203 vdd.n202 1.13717
R3457 vdd.n1461 vdd.n201 1.13717
R3458 vdd.n1491 vdd.n184 1.13717
R3459 vdd.n1514 vdd.n172 1.13717
R3460 vdd.n157 vdd.n156 1.13717
R3461 vdd.n1544 vdd.n155 1.13717
R3462 vdd.n1576 vdd.n1575 1.13717
R3463 vdd.n1598 vdd.n1597 1.13717
R3464 vdd.n106 vdd.n105 1.13717
R3465 vdd.n1633 vdd.n1632 1.13717
R3466 vdd.n1656 vdd.n1655 1.13717
R3467 vdd.n1660 vdd.n1659 1.13717
R3468 vdd.n1880 vdd.n1876 1.13717
R3469 vdd.n1895 vdd.n1891 1.13717
R3470 vdd.n1906 vdd.n1902 1.13717
R3471 vdd.n1917 vdd.n1913 1.13717
R3472 vdd.n1928 vdd.n1924 1.13717
R3473 vdd.n3718 vdd.n1935 1.13717
R3474 vdd.n3726 vdd.n3725 1.13717
R3475 vdd.n3745 vdd.n3744 1.13717
R3476 vdd.n3764 vdd.n3763 1.13717
R3477 vdd.n3783 vdd.n3782 1.13717
R3478 vdd.n3802 vdd.n3801 1.13717
R3479 vdd.n3821 vdd.n3820 1.13717
R3480 vdd.n3698 vdd.n3697 1.13717
R3481 vdd.n2823 vdd.n2464 1.13717
R3482 vdd.n1938 vdd.n1937 1.13717
R3483 vdd.n3694 vdd.n3693 1.13717
R3484 vdd.n1952 vdd.n1947 1.13717
R3485 vdd.n3673 vdd.n3672 1.13717
R3486 vdd.n1965 vdd.n1963 1.13717
R3487 vdd.n1969 vdd.n1968 1.13717
R3488 vdd.n3666 vdd.n3665 1.13717
R3489 vdd.n3635 vdd.n1980 1.13717
R3490 vdd.n3643 vdd.n3642 1.13717
R3491 vdd.n3611 vdd.n3610 1.13717
R3492 vdd.n1995 vdd.n1983 1.13717
R3493 vdd.n3523 vdd.n2054 1.13717
R3494 vdd.n3521 vdd.n2053 1.13717
R3495 vdd.n3543 vdd.n2044 1.13717
R3496 vdd.n3542 vdd.n3541 1.13717
R3497 vdd.n2031 vdd.n2030 1.13717
R3498 vdd.n3549 vdd.n2032 1.13717
R3499 vdd.n2020 vdd.n2019 1.13717
R3500 vdd.n3571 vdd.n2021 1.13717
R3501 vdd.n1998 vdd.n1997 1.13717
R3502 vdd.n3591 vdd.n1999 1.13717
R3503 vdd.n3503 vdd.n2065 1.13717
R3504 vdd.n3501 vdd.n2064 1.13717
R3505 vdd.n3492 vdd.n3491 1.13717
R3506 vdd.n2073 vdd.n2069 1.13717
R3507 vdd.n3468 vdd.n3467 1.13717
R3508 vdd.n2086 vdd.n2082 1.13717
R3509 vdd.n3447 vdd.n3446 1.13717
R3510 vdd.n2099 vdd.n2097 1.13717
R3511 vdd.n2103 vdd.n2102 1.13717
R3512 vdd.n3440 vdd.n3439 1.13717
R3513 vdd.n3409 vdd.n2114 1.13717
R3514 vdd.n3417 vdd.n3416 1.13717
R3515 vdd.n3385 vdd.n3384 1.13717
R3516 vdd.n2129 vdd.n2117 1.13717
R3517 vdd.n3297 vdd.n2188 1.13717
R3518 vdd.n3295 vdd.n2187 1.13717
R3519 vdd.n3317 vdd.n2178 1.13717
R3520 vdd.n3316 vdd.n3315 1.13717
R3521 vdd.n2165 vdd.n2164 1.13717
R3522 vdd.n3323 vdd.n2166 1.13717
R3523 vdd.n2154 vdd.n2153 1.13717
R3524 vdd.n3345 vdd.n2155 1.13717
R3525 vdd.n2132 vdd.n2131 1.13717
R3526 vdd.n3365 vdd.n2133 1.13717
R3527 vdd.n3277 vdd.n2199 1.13717
R3528 vdd.n3275 vdd.n2198 1.13717
R3529 vdd.n3266 vdd.n3265 1.13717
R3530 vdd.n2207 vdd.n2203 1.13717
R3531 vdd.n3242 vdd.n3241 1.13717
R3532 vdd.n2220 vdd.n2216 1.13717
R3533 vdd.n3221 vdd.n3220 1.13717
R3534 vdd.n2233 vdd.n2231 1.13717
R3535 vdd.n2237 vdd.n2236 1.13717
R3536 vdd.n3214 vdd.n3213 1.13717
R3537 vdd.n3183 vdd.n2248 1.13717
R3538 vdd.n3191 vdd.n3190 1.13717
R3539 vdd.n3159 vdd.n3158 1.13717
R3540 vdd.n2263 vdd.n2251 1.13717
R3541 vdd.n3071 vdd.n2322 1.13717
R3542 vdd.n3069 vdd.n2321 1.13717
R3543 vdd.n3091 vdd.n2312 1.13717
R3544 vdd.n3090 vdd.n3089 1.13717
R3545 vdd.n2299 vdd.n2298 1.13717
R3546 vdd.n3097 vdd.n2300 1.13717
R3547 vdd.n2288 vdd.n2287 1.13717
R3548 vdd.n3119 vdd.n2289 1.13717
R3549 vdd.n2266 vdd.n2265 1.13717
R3550 vdd.n3139 vdd.n2267 1.13717
R3551 vdd.n3051 vdd.n2333 1.13717
R3552 vdd.n3049 vdd.n2332 1.13717
R3553 vdd.n3040 vdd.n3039 1.13717
R3554 vdd.n2341 vdd.n2337 1.13717
R3555 vdd.n3016 vdd.n3015 1.13717
R3556 vdd.n2354 vdd.n2350 1.13717
R3557 vdd.n2995 vdd.n2994 1.13717
R3558 vdd.n2367 vdd.n2365 1.13717
R3559 vdd.n2371 vdd.n2370 1.13717
R3560 vdd.n2988 vdd.n2987 1.13717
R3561 vdd.n2957 vdd.n2382 1.13717
R3562 vdd.n2965 vdd.n2964 1.13717
R3563 vdd.n2933 vdd.n2932 1.13717
R3564 vdd.n2397 vdd.n2385 1.13717
R3565 vdd.n2865 vdd.n2446 1.13717
R3566 vdd.n2864 vdd.n2863 1.13717
R3567 vdd.n2433 vdd.n2432 1.13717
R3568 vdd.n2871 vdd.n2434 1.13717
R3569 vdd.n2422 vdd.n2421 1.13717
R3570 vdd.n2893 vdd.n2423 1.13717
R3571 vdd.n2400 vdd.n2399 1.13717
R3572 vdd.n2913 vdd.n2401 1.13717
R3573 vdd.n2843 vdd.n2455 1.13717
R3574 vdd.n2845 vdd.n2456 1.13717
R3575 vdd.n2825 vdd.n2465 1.13717
R3576 vdd.n2802 vdd.n2780 1.13717
R3577 vdd.n619 vdd.n618 1.13462
R3578 vdd.n626 vdd.n625 1.13462
R3579 vdd.n630 vdd.n629 1.13462
R3580 vdd.n641 vdd.n640 1.13462
R3581 vdd.n689 vdd.n612 1.13462
R3582 vdd.n2479 vdd.n2478 1.13462
R3583 vdd.n2475 vdd.n2474 1.13462
R3584 vdd.n2501 vdd.n2473 1.13462
R3585 vdd.n2468 vdd.n2467 1.13462
R3586 vdd.n2748 vdd.n2511 1.13462
R3587 vdd.n659 vdd.n658 1.13005
R3588 vdd.n2738 vdd.n2737 1.13005
R3589 vdd.n2535 vdd.n2521 1.08374
R3590 vdd.n2535 vdd.n2534 1.08374
R3591 vdd.n694 vdd.n693 1.04017
R3592 vdd.n645 vdd.n644 1.04017
R3593 vdd.n638 vdd.n637 1.04017
R3594 vdd.n634 vdd.n633 1.04017
R3595 vdd.n623 vdd.n622 1.04017
R3596 vdd.n2753 vdd.n2752 1.04017
R3597 vdd.n2816 vdd.n2815 1.04017
R3598 vdd.n2506 vdd.n2505 1.04017
R3599 vdd.n2488 vdd.n2487 1.04017
R3600 vdd.n2494 vdd.n2493 1.04017
R3601 vdd.n1832 vdd.n1831 1.01637
R3602 vdd.n2806 vdd.n2758 1.01637
R3603 vdd vdd.n2583 0.91916
R3604 vdd.t0 vdd 0.918966
R3605 vdd.n2767 vdd.n2766 0.870766
R3606 vdd.n1810 vdd.n1809 0.870578
R3607 vdd.n1799 vdd.n1798 0.870578
R3608 vdd.n2799 vdd.n2786 0.870578
R3609 vdd.n2669 vdd.n2667 0.857916
R3610 vdd.n652 vdd.n651 0.853291
R3611 vdd.n2731 vdd.n2730 0.853291
R3612 vdd.n1866 vdd.n2 0.853
R3613 vdd.n687 vdd.n620 0.853
R3614 vdd.n684 vdd.n627 0.853
R3615 vdd.n681 vdd.n631 0.853
R3616 vdd.n678 vdd.n642 0.853
R3617 vdd.n692 vdd.n691 0.853
R3618 vdd.n1819 vdd.n1817 0.853
R3619 vdd.n3831 vdd.n1872 0.853
R3620 vdd.n2496 vdd.n2480 0.853
R3621 vdd.n2499 vdd.n2476 0.853
R3622 vdd.n2504 vdd.n2503 0.853
R3623 vdd.n2818 vdd.n2470 0.853
R3624 vdd.n2751 vdd.n2750 0.853
R3625 vdd.n2513 vdd.n2512 0.853
R3626 vdd.n2696 vdd.n2695 0.853
R3627 vdd.n2546 vdd.n2545 0.853
R3628 vdd.n2655 vdd.n2654 0.853
R3629 vdd.n2544 vdd.n2543 0.853
R3630 vdd.n2803 vdd.n2802 0.853
R3631 vdd.n3723 vdd.n3722 0.849634
R3632 vdd.n1688 vdd.n1686 0.849012
R3633 vdd.n1838 vdd.n1786 0.813198
R3634 vdd.n1831 vdd.n1824 0.813198
R3635 vdd.n2773 vdd.n2772 0.813198
R3636 vdd.n2806 vdd.n2759 0.813198
R3637 vdd.n635 vdd.n609 0.734658
R3638 vdd.n697 vdd.n595 0.734658
R3639 vdd.n725 vdd.n724 0.734658
R3640 vdd.n749 vdd.n748 0.734658
R3641 vdd.n777 vdd.n564 0.734658
R3642 vdd.n779 vdd.n550 0.734658
R3643 vdd.n805 vdd.n803 0.734658
R3644 vdd.n841 vdd.n530 0.734658
R3645 vdd.n843 vdd.n514 0.734658
R3646 vdd.n866 vdd.n865 0.734658
R3647 vdd.n887 vdd.n886 0.734658
R3648 vdd.n938 vdd.n481 0.734658
R3649 vdd.n940 vdd.n476 0.734658
R3650 vdd.n948 vdd.n461 0.734658
R3651 vdd.n976 vdd.n975 0.734658
R3652 vdd.n1000 vdd.n999 0.734658
R3653 vdd.n1028 vdd.n430 0.734658
R3654 vdd.n1030 vdd.n416 0.734658
R3655 vdd.n1056 vdd.n1054 0.734658
R3656 vdd.n1092 vdd.n396 0.734658
R3657 vdd.n1094 vdd.n380 0.734658
R3658 vdd.n1117 vdd.n1116 0.734658
R3659 vdd.n1138 vdd.n1137 0.734658
R3660 vdd.n1189 vdd.n347 0.734658
R3661 vdd.n1191 vdd.n342 0.734658
R3662 vdd.n1199 vdd.n327 0.734658
R3663 vdd.n1227 vdd.n1226 0.734658
R3664 vdd.n1251 vdd.n1250 0.734658
R3665 vdd.n1279 vdd.n296 0.734658
R3666 vdd.n1281 vdd.n282 0.734658
R3667 vdd.n1307 vdd.n1305 0.734658
R3668 vdd.n1343 vdd.n262 0.734658
R3669 vdd.n1345 vdd.n246 0.734658
R3670 vdd.n1368 vdd.n1367 0.734658
R3671 vdd.n1389 vdd.n1388 0.734658
R3672 vdd.n1440 vdd.n213 0.734658
R3673 vdd.n1442 vdd.n208 0.734658
R3674 vdd.n1450 vdd.n193 0.734658
R3675 vdd.n1478 vdd.n1477 0.734658
R3676 vdd.n1502 vdd.n1501 0.734658
R3677 vdd.n1530 vdd.n162 0.734658
R3678 vdd.n1532 vdd.n148 0.734658
R3679 vdd.n1558 vdd.n1556 0.734658
R3680 vdd.n1589 vdd.n129 0.734658
R3681 vdd.n1591 vdd.n112 0.734658
R3682 vdd.n1614 vdd.n1613 0.734658
R3683 vdd.n1645 vdd.n1644 0.734658
R3684 vdd.n1674 vdd.n80 0.734658
R3685 vdd.n1678 vdd.n1677 0.734658
R3686 vdd.n1704 vdd.n65 0.734658
R3687 vdd.n1706 vdd.n48 0.734658
R3688 vdd.n1729 vdd.n1728 0.734658
R3689 vdd.n1760 vdd.n1759 0.734658
R3690 vdd.n1784 vdd.n17 0.734658
R3691 vdd.n1849 vdd.n1848 0.734658
R3692 vdd.n3834 vdd 0.685225
R3693 vdd.n649 vdd.n648 0.684595
R3694 vdd.n2743 vdd.n2741 0.684595
R3695 vdd.n2682 vdd.n2681 0.684469
R3696 vdd.n1802 vdd.n1801 0.682713
R3697 vdd.n1813 vdd.n1812 0.682713
R3698 vdd.n2798 vdd.n2782 0.682713
R3699 vdd.n2770 vdd.n2769 0.682713
R3700 vdd.n2727 vdd.n2726 0.682697
R3701 vdd.n2692 vdd.n2691 0.682639
R3702 vdd.n2657 vdd.n2656 0.682639
R3703 vdd.n2687 vdd.n2686 0.682639
R3704 vdd.n2698 vdd.n2697 0.682639
R3705 vdd.n1867 vdd.n3 0.682447
R3706 vdd.n3832 vdd.n1873 0.682447
R3707 vdd.t61 vdd.n2490 0.612811
R3708 vdd.n2700 vdd.n2538 0.58676
R3709 vdd.n2619 vdd.n2618 0.551696
R3710 vdd.n804 vdd 0.534441
R3711 vdd.n1055 vdd 0.534441
R3712 vdd.n1306 vdd 0.534441
R3713 vdd.n1557 vdd 0.534441
R3714 vdd.t32 vdd.n2754 0.459883
R3715 vdd.n1942 vdd.n1886 0.459733
R3716 vdd.n2754 vdd.t11 0.457214
R3717 vdd.n1791 vdd.n1790 0.406849
R3718 vdd.n2795 vdd.n2794 0.406849
R3719 vdd.n2648 vdd.n2563 0.367964
R3720 vdd.n661 vdd.n660 0.357419
R3721 vdd.n914 vdd.n473 0.314894
R3722 vdd.n1165 vdd.n339 0.314894
R3723 vdd.n1416 vdd.n205 0.314894
R3724 vdd.n2343 vdd.n2331 0.314894
R3725 vdd.n2209 vdd.n2197 0.314894
R3726 vdd.n2075 vdd.n2063 0.314894
R3727 vdd.n2740 vdd.n2739 0.312073
R3728 vdd.n2714 vdd.n2525 0.309679
R3729 vdd.n2713 vdd.n2712 0.309679
R3730 vdd.n2712 vdd.n2529 0.309679
R3731 vdd.n2598 vdd.n2597 0.30672
R3732 vdd.n2627 vdd.n2556 0.30672
R3733 vdd.n2812 vdd.n2811 0.306655
R3734 vdd.n813 vdd.n544 0.30353
R3735 vdd.n1064 vdd.n410 0.30353
R3736 vdd.n1315 vdd.n276 0.30353
R3737 vdd.n1566 vdd.n142 0.30353
R3738 vdd.n812 vdd.n811 0.30353
R3739 vdd.n1063 vdd.n1062 0.30353
R3740 vdd.n1314 vdd.n1313 0.30353
R3741 vdd.n1565 vdd.n1564 0.30353
R3742 vdd.n2411 vdd.n2408 0.30353
R3743 vdd.n2277 vdd.n2274 0.30353
R3744 vdd.n2143 vdd.n2140 0.30353
R3745 vdd.n2009 vdd.n2006 0.30353
R3746 vdd.n2410 vdd.n2409 0.30353
R3747 vdd.n2276 vdd.n2275 0.30353
R3748 vdd.n2142 vdd.n2141 0.30353
R3749 vdd.n2008 vdd.n2007 0.30353
R3750 vdd.n918 vdd.n916 0.288379
R3751 vdd.n1169 vdd.n1167 0.288379
R3752 vdd.n1420 vdd.n1418 0.288379
R3753 vdd.n3047 vdd.n3045 0.288379
R3754 vdd.n3273 vdd.n3271 0.288379
R3755 vdd.n3499 vdd.n3497 0.288379
R3756 vdd.n2585 vdd.n2584 0.245476
R3757 vdd.n1 vdd.n0 0.2355
R3758 vdd.n2801 vdd.n1871 0.2355
R3759 vdd.n2709 vdd.n2531 0.19592
R3760 vdd.n700 vdd.n597 0.194439
R3761 vdd.n727 vdd.n592 0.194439
R3762 vdd.n728 vdd.n727 0.194439
R3763 vdd.n746 vdd.n745 0.194439
R3764 vdd.n745 vdd.n579 0.194439
R3765 vdd.n775 vdd.n566 0.194439
R3766 vdd.n775 vdd.n567 0.194439
R3767 vdd.n782 vdd.n781 0.194439
R3768 vdd.n782 vdd.n552 0.194439
R3769 vdd.n807 vdd.n548 0.194439
R3770 vdd.n807 vdd.n542 0.194439
R3771 vdd.n817 vdd.n532 0.194439
R3772 vdd.n839 vdd.n532 0.194439
R3773 vdd.n845 vdd.n528 0.194439
R3774 vdd.n845 vdd.n516 0.194439
R3775 vdd.n517 vdd.n512 0.194439
R3776 vdd.n868 vdd.n512 0.194439
R3777 vdd.n884 vdd.n503 0.194439
R3778 vdd.n884 vdd.n499 0.194439
R3779 vdd.n891 vdd.n483 0.194439
R3780 vdd.n936 vdd.n483 0.194439
R3781 vdd.n942 vdd.n478 0.194439
R3782 vdd.n943 vdd.n942 0.194439
R3783 vdd.n951 vdd.n950 0.194439
R3784 vdd.n951 vdd.n463 0.194439
R3785 vdd.n978 vdd.n458 0.194439
R3786 vdd.n979 vdd.n978 0.194439
R3787 vdd.n997 vdd.n996 0.194439
R3788 vdd.n996 vdd.n445 0.194439
R3789 vdd.n1026 vdd.n432 0.194439
R3790 vdd.n1026 vdd.n433 0.194439
R3791 vdd.n1033 vdd.n1032 0.194439
R3792 vdd.n1033 vdd.n418 0.194439
R3793 vdd.n1058 vdd.n414 0.194439
R3794 vdd.n1058 vdd.n408 0.194439
R3795 vdd.n1068 vdd.n398 0.194439
R3796 vdd.n1090 vdd.n398 0.194439
R3797 vdd.n1096 vdd.n394 0.194439
R3798 vdd.n1096 vdd.n382 0.194439
R3799 vdd.n383 vdd.n378 0.194439
R3800 vdd.n1119 vdd.n378 0.194439
R3801 vdd.n1135 vdd.n369 0.194439
R3802 vdd.n1135 vdd.n365 0.194439
R3803 vdd.n1142 vdd.n349 0.194439
R3804 vdd.n1187 vdd.n349 0.194439
R3805 vdd.n1193 vdd.n344 0.194439
R3806 vdd.n1194 vdd.n1193 0.194439
R3807 vdd.n1202 vdd.n1201 0.194439
R3808 vdd.n1202 vdd.n329 0.194439
R3809 vdd.n1229 vdd.n324 0.194439
R3810 vdd.n1230 vdd.n1229 0.194439
R3811 vdd.n1248 vdd.n1247 0.194439
R3812 vdd.n1247 vdd.n311 0.194439
R3813 vdd.n1277 vdd.n298 0.194439
R3814 vdd.n1277 vdd.n299 0.194439
R3815 vdd.n1284 vdd.n1283 0.194439
R3816 vdd.n1284 vdd.n284 0.194439
R3817 vdd.n1309 vdd.n280 0.194439
R3818 vdd.n1309 vdd.n274 0.194439
R3819 vdd.n1319 vdd.n264 0.194439
R3820 vdd.n1341 vdd.n264 0.194439
R3821 vdd.n1347 vdd.n260 0.194439
R3822 vdd.n1347 vdd.n248 0.194439
R3823 vdd.n249 vdd.n244 0.194439
R3824 vdd.n1370 vdd.n244 0.194439
R3825 vdd.n1386 vdd.n235 0.194439
R3826 vdd.n1386 vdd.n231 0.194439
R3827 vdd.n1393 vdd.n215 0.194439
R3828 vdd.n1438 vdd.n215 0.194439
R3829 vdd.n1444 vdd.n210 0.194439
R3830 vdd.n1445 vdd.n1444 0.194439
R3831 vdd.n1453 vdd.n1452 0.194439
R3832 vdd.n1453 vdd.n195 0.194439
R3833 vdd.n1480 vdd.n190 0.194439
R3834 vdd.n1481 vdd.n1480 0.194439
R3835 vdd.n1499 vdd.n1498 0.194439
R3836 vdd.n1498 vdd.n177 0.194439
R3837 vdd.n1528 vdd.n164 0.194439
R3838 vdd.n1528 vdd.n165 0.194439
R3839 vdd.n1535 vdd.n1534 0.194439
R3840 vdd.n1535 vdd.n150 0.194439
R3841 vdd.n1560 vdd.n146 0.194439
R3842 vdd.n1560 vdd.n140 0.194439
R3843 vdd.n1570 vdd.n131 0.194439
R3844 vdd.n1587 vdd.n131 0.194439
R3845 vdd.n1593 vdd.n127 0.194439
R3846 vdd.n1593 vdd.n114 0.194439
R3847 vdd.n115 vdd.n110 0.194439
R3848 vdd.n1616 vdd.n110 0.194439
R3849 vdd.n1642 vdd.n96 0.194439
R3850 vdd.n1642 vdd.n92 0.194439
R3851 vdd.n1650 vdd.n82 0.194439
R3852 vdd.n1672 vdd.n82 0.194439
R3853 vdd.n1680 vdd.n76 0.194439
R3854 vdd.n1702 vdd.n67 0.194439
R3855 vdd.n1708 vdd.n63 0.194439
R3856 vdd.n1708 vdd.n50 0.194439
R3857 vdd.n51 vdd.n46 0.194439
R3858 vdd.n1731 vdd.n46 0.194439
R3859 vdd.n1757 vdd.n32 0.194439
R3860 vdd.n1757 vdd.n28 0.194439
R3861 vdd.n1765 vdd.n19 0.194439
R3862 vdd.n1782 vdd.n19 0.194439
R3863 vdd.n1851 vdd.n13 0.194439
R3864 vdd.n1851 vdd.n14 0.194439
R3865 vdd.n2831 vdd.n2462 0.194439
R3866 vdd.n2852 vdd.n2453 0.194439
R3867 vdd.n2852 vdd.n2451 0.194439
R3868 vdd.n2879 vdd.n2438 0.194439
R3869 vdd.n2879 vdd.n2439 0.194439
R3870 vdd.n2885 vdd.n2884 0.194439
R3871 vdd.n2885 vdd.n2427 0.194439
R3872 vdd.n2905 vdd.n2425 0.194439
R3873 vdd.n2905 vdd.n2416 0.194439
R3874 vdd.n2924 vdd.n2405 0.194439
R3875 vdd.n2924 vdd.n2414 0.194439
R3876 vdd.n2937 vdd.n2394 0.194439
R3877 vdd.n2937 vdd.n2393 0.194439
R3878 vdd.n2946 vdd.n2945 0.194439
R3879 vdd.n2945 vdd.n2392 0.194439
R3880 vdd.n2973 vdd.n2972 0.194439
R3881 vdd.n2973 vdd.n2375 0.194439
R3882 vdd.n3004 vdd.n2359 0.194439
R3883 vdd.n3005 vdd.n3004 0.194439
R3884 vdd.n3011 vdd.n2356 0.194439
R3885 vdd.n3011 vdd.n2347 0.194439
R3886 vdd.n3035 vdd.n2344 0.194439
R3887 vdd.n3035 vdd.n2345 0.194439
R3888 vdd.n3057 vdd.n2330 0.194439
R3889 vdd.n3057 vdd.n2328 0.194439
R3890 vdd.n3078 vdd.n2319 0.194439
R3891 vdd.n3078 vdd.n2317 0.194439
R3892 vdd.n3105 vdd.n2304 0.194439
R3893 vdd.n3105 vdd.n2305 0.194439
R3894 vdd.n3111 vdd.n3110 0.194439
R3895 vdd.n3111 vdd.n2293 0.194439
R3896 vdd.n3131 vdd.n2291 0.194439
R3897 vdd.n3131 vdd.n2282 0.194439
R3898 vdd.n3150 vdd.n2271 0.194439
R3899 vdd.n3150 vdd.n2280 0.194439
R3900 vdd.n3163 vdd.n2260 0.194439
R3901 vdd.n3163 vdd.n2259 0.194439
R3902 vdd.n3172 vdd.n3171 0.194439
R3903 vdd.n3171 vdd.n2258 0.194439
R3904 vdd.n3199 vdd.n3198 0.194439
R3905 vdd.n3199 vdd.n2241 0.194439
R3906 vdd.n3230 vdd.n2225 0.194439
R3907 vdd.n3231 vdd.n3230 0.194439
R3908 vdd.n3237 vdd.n2222 0.194439
R3909 vdd.n3237 vdd.n2213 0.194439
R3910 vdd.n3261 vdd.n2210 0.194439
R3911 vdd.n3261 vdd.n2211 0.194439
R3912 vdd.n3283 vdd.n2196 0.194439
R3913 vdd.n3283 vdd.n2194 0.194439
R3914 vdd.n3304 vdd.n2185 0.194439
R3915 vdd.n3304 vdd.n2183 0.194439
R3916 vdd.n3331 vdd.n2170 0.194439
R3917 vdd.n3331 vdd.n2171 0.194439
R3918 vdd.n3337 vdd.n3336 0.194439
R3919 vdd.n3337 vdd.n2159 0.194439
R3920 vdd.n3357 vdd.n2157 0.194439
R3921 vdd.n3357 vdd.n2148 0.194439
R3922 vdd.n3376 vdd.n2137 0.194439
R3923 vdd.n3376 vdd.n2146 0.194439
R3924 vdd.n3389 vdd.n2126 0.194439
R3925 vdd.n3389 vdd.n2125 0.194439
R3926 vdd.n3398 vdd.n3397 0.194439
R3927 vdd.n3397 vdd.n2124 0.194439
R3928 vdd.n3425 vdd.n3424 0.194439
R3929 vdd.n3425 vdd.n2107 0.194439
R3930 vdd.n3456 vdd.n2091 0.194439
R3931 vdd.n3457 vdd.n3456 0.194439
R3932 vdd.n3463 vdd.n2088 0.194439
R3933 vdd.n3463 vdd.n2079 0.194439
R3934 vdd.n3487 vdd.n2076 0.194439
R3935 vdd.n3487 vdd.n2077 0.194439
R3936 vdd.n3509 vdd.n2062 0.194439
R3937 vdd.n3509 vdd.n2060 0.194439
R3938 vdd.n3530 vdd.n2051 0.194439
R3939 vdd.n3530 vdd.n2049 0.194439
R3940 vdd.n3557 vdd.n2036 0.194439
R3941 vdd.n3557 vdd.n2037 0.194439
R3942 vdd.n3563 vdd.n3562 0.194439
R3943 vdd.n3563 vdd.n2025 0.194439
R3944 vdd.n3583 vdd.n2023 0.194439
R3945 vdd.n3583 vdd.n2014 0.194439
R3946 vdd.n3602 vdd.n2003 0.194439
R3947 vdd.n3602 vdd.n2012 0.194439
R3948 vdd.n3615 vdd.n1992 0.194439
R3949 vdd.n3615 vdd.n1991 0.194439
R3950 vdd.n3624 vdd.n3623 0.194439
R3951 vdd.n3623 vdd.n1990 0.194439
R3952 vdd.n3651 vdd.n3650 0.194439
R3953 vdd.n3651 vdd.n1973 0.194439
R3954 vdd.n3682 vdd.n1957 0.194439
R3955 vdd.n3683 vdd.n3682 0.194439
R3956 vdd.n3689 vdd.n1954 0.194439
R3957 vdd.n3689 vdd.n1944 0.194439
R3958 vdd.n3712 vdd.n1941 0.194439
R3959 vdd.n3721 vdd.n1932 0.194439
R3960 vdd.n3740 vdd.n1930 0.194439
R3961 vdd.n3740 vdd.n1921 0.194439
R3962 vdd.n3759 vdd.n1919 0.194439
R3963 vdd.n3759 vdd.n1910 0.194439
R3964 vdd.n3778 vdd.n1908 0.194439
R3965 vdd.n3778 vdd.n1899 0.194439
R3966 vdd.n3797 vdd.n1897 0.194439
R3967 vdd.n3797 vdd.n1888 0.194439
R3968 vdd.n3816 vdd.n1883 0.194439
R3969 vdd.n3816 vdd.n1884 0.194439
R3970 vdd.n2583 vdd.n2578 0.184232
R3971 vdd.n2650 vdd.n2562 0.184232
R3972 vdd.n2663 vdd.n2553 0.184232
R3973 vdd.n1869 vdd 0.142102
R3974 vdd.n1843 vdd.n1842 0.132407
R3975 vdd.n2484 vdd.n2483 0.132407
R3976 vdd.n1842 vdd.n12 0.127283
R3977 vdd.n2483 vdd.n1882 0.127283
R3978 vdd.n2718 vdd.n2717 0.124172
R3979 vdd.n2587 vdd.n2585 0.122988
R3980 vdd.n2614 vdd.n2613 0.122988
R3981 vdd.n2635 vdd.n2634 0.122988
R3982 vdd.n2637 vdd.n2636 0.122988
R3983 vdd.n2586 vdd.n2576 0.120292
R3984 vdd.n2593 vdd.n2576 0.120292
R3985 vdd.n2594 vdd.n2593 0.120292
R3986 vdd.n2596 vdd.n2594 0.120292
R3987 vdd.n2596 vdd.n2595 0.120292
R3988 vdd.n2595 vdd.n2569 0.120292
R3989 vdd.n2602 vdd.n2588 0.120292
R3990 vdd.n2602 vdd.n2601 0.120292
R3991 vdd.n2601 vdd.n2600 0.120292
R3992 vdd.n2600 vdd.n2589 0.120292
R3993 vdd.n2589 vdd.n2570 0.120292
R3994 vdd.n2615 vdd.n2570 0.120292
R3995 vdd.n617 vdd 0.103754
R3996 vdd.n789 vdd.n538 0.102103
R3997 vdd.n1040 vdd.n404 0.102103
R3998 vdd.n1291 vdd.n270 0.102103
R3999 vdd.n1542 vdd.n136 0.102103
R4000 vdd.n2928 vdd.n2398 0.102103
R4001 vdd.n3154 vdd.n2264 0.102103
R4002 vdd.n3380 vdd.n2130 0.102103
R4003 vdd.n3606 vdd.n1996 0.102103
R4004 vdd.n924 vdd.n923 0.100721
R4005 vdd.n1175 vdd.n1174 0.100721
R4006 vdd.n1426 vdd.n1425 0.100721
R4007 vdd.n3043 vdd.n2335 0.100721
R4008 vdd.n3269 vdd.n2201 0.100721
R4009 vdd.n3495 vdd.n2067 0.100721
R4010 vdd.n1685 vdd 0.100533
R4011 vdd.n3717 vdd 0.100533
R4012 vdd.n1836 vdd.n1835 0.0981562
R4013 vdd.n2777 vdd.n2765 0.0981562
R4014 vdd.n2616 vdd 0.0968542
R4015 vdd.n790 vdd.n537 0.0890769
R4016 vdd.n1041 vdd.n403 0.0890769
R4017 vdd.n1292 vdd.n269 0.0890769
R4018 vdd.n1543 vdd.n135 0.0890769
R4019 vdd.n2930 vdd.n2929 0.0890769
R4020 vdd.n3156 vdd.n3155 0.0890769
R4021 vdd.n3382 vdd.n3381 0.0890769
R4022 vdd.n3608 vdd.n3607 0.0890769
R4023 vdd.n3653 vdd.n3652 0.0847059
R4024 vdd.n3688 vdd.n3687 0.0847059
R4025 vdd.n3427 vdd.n3426 0.0847059
R4026 vdd.n3462 vdd.n3461 0.0847059
R4027 vdd.n3201 vdd.n3200 0.0847059
R4028 vdd.n3236 vdd.n3235 0.0847059
R4029 vdd.n2975 vdd.n2974 0.0847059
R4030 vdd.n3010 vdd.n3009 0.0847059
R4031 vdd.n2853 vdd.n2452 0.0847059
R4032 vdd.n3739 vdd.n3738 0.0847059
R4033 vdd.n3758 vdd.n3757 0.0847059
R4034 vdd.n3777 vdd.n3776 0.0847059
R4035 vdd.n3796 vdd.n3795 0.0847059
R4036 vdd.n2616 vdd.n2569 0.0838333
R4037 vdd.n2616 vdd.n2615 0.0838333
R4038 vdd.n1864 vdd.n1863 0.0796667
R4039 vdd.n3829 vdd.n3828 0.0796667
R4040 vdd.n3834 vdd 0.0794477
R4041 vdd.n718 vdd.n599 0.0705758
R4042 vdd.n731 vdd.n584 0.0705758
R4043 vdd.n755 vdd.n568 0.0705758
R4044 vdd.n770 vdd.n561 0.0705758
R4045 vdd.n797 vdd.n547 0.0705758
R4046 vdd.n835 vdd.n533 0.0705758
R4047 vdd.n847 vdd.n518 0.0705758
R4048 vdd.n872 vdd.n511 0.0705758
R4049 vdd.n894 vdd.n498 0.0705758
R4050 vdd.n906 vdd.n484 0.0705758
R4051 vdd.n969 vdd.n465 0.0705758
R4052 vdd.n982 vdd.n450 0.0705758
R4053 vdd.n1006 vdd.n434 0.0705758
R4054 vdd.n1021 vdd.n427 0.0705758
R4055 vdd.n1048 vdd.n413 0.0705758
R4056 vdd.n1086 vdd.n399 0.0705758
R4057 vdd.n1098 vdd.n384 0.0705758
R4058 vdd.n1123 vdd.n377 0.0705758
R4059 vdd.n1145 vdd.n364 0.0705758
R4060 vdd.n1157 vdd.n350 0.0705758
R4061 vdd.n1220 vdd.n331 0.0705758
R4062 vdd.n1233 vdd.n316 0.0705758
R4063 vdd.n1257 vdd.n300 0.0705758
R4064 vdd.n1272 vdd.n293 0.0705758
R4065 vdd.n1299 vdd.n279 0.0705758
R4066 vdd.n1337 vdd.n265 0.0705758
R4067 vdd.n1349 vdd.n250 0.0705758
R4068 vdd.n1374 vdd.n243 0.0705758
R4069 vdd.n1396 vdd.n230 0.0705758
R4070 vdd.n1408 vdd.n216 0.0705758
R4071 vdd.n1471 vdd.n197 0.0705758
R4072 vdd.n1484 vdd.n182 0.0705758
R4073 vdd.n1508 vdd.n166 0.0705758
R4074 vdd.n1523 vdd.n159 0.0705758
R4075 vdd.n1550 vdd.n145 0.0705758
R4076 vdd.n1583 vdd.n132 0.0705758
R4077 vdd.n126 vdd.n116 0.0705758
R4078 vdd.n1623 vdd.n1622 0.0705758
R4079 vdd.n1640 vdd.n99 0.0705758
R4080 vdd.n1668 vdd.n83 0.0705758
R4081 vdd.n1698 vdd.n68 0.0705758
R4082 vdd.n62 vdd.n52 0.0705758
R4083 vdd.n1738 vdd.n1737 0.0705758
R4084 vdd.n1755 vdd.n35 0.0705758
R4085 vdd.n1778 vdd.n20 0.0705758
R4086 vdd.n2838 vdd.n2454 0.0705758
R4087 vdd.n2859 vdd.n2440 0.0705758
R4088 vdd.n2874 vdd.n2435 0.0705758
R4089 vdd.n2897 vdd.n2424 0.0705758
R4090 vdd.n2917 vdd.n2403 0.0705758
R4091 vdd.n2949 vdd.n2388 0.0705758
R4092 vdd.n2968 vdd.n2967 0.0705758
R4093 vdd.n2985 vdd.n2984 0.0705758
R4094 vdd.n3002 vdd.n2364 0.0705758
R4095 vdd.n3023 vdd.n2348 0.0705758
R4096 vdd.n3064 vdd.n2320 0.0705758
R4097 vdd.n3085 vdd.n2306 0.0705758
R4098 vdd.n3100 vdd.n2301 0.0705758
R4099 vdd.n3123 vdd.n2290 0.0705758
R4100 vdd.n3143 vdd.n2269 0.0705758
R4101 vdd.n3175 vdd.n2254 0.0705758
R4102 vdd.n3194 vdd.n3193 0.0705758
R4103 vdd.n3211 vdd.n3210 0.0705758
R4104 vdd.n3228 vdd.n2230 0.0705758
R4105 vdd.n3249 vdd.n2214 0.0705758
R4106 vdd.n3290 vdd.n2186 0.0705758
R4107 vdd.n3311 vdd.n2172 0.0705758
R4108 vdd.n3326 vdd.n2167 0.0705758
R4109 vdd.n3349 vdd.n2156 0.0705758
R4110 vdd.n3369 vdd.n2135 0.0705758
R4111 vdd.n3401 vdd.n2120 0.0705758
R4112 vdd.n3420 vdd.n3419 0.0705758
R4113 vdd.n3437 vdd.n3436 0.0705758
R4114 vdd.n3454 vdd.n2096 0.0705758
R4115 vdd.n3475 vdd.n2080 0.0705758
R4116 vdd.n3516 vdd.n2052 0.0705758
R4117 vdd.n3537 vdd.n2038 0.0705758
R4118 vdd.n3552 vdd.n2033 0.0705758
R4119 vdd.n3575 vdd.n2022 0.0705758
R4120 vdd.n3595 vdd.n2001 0.0705758
R4121 vdd.n3627 vdd.n1986 0.0705758
R4122 vdd.n3646 vdd.n3645 0.0705758
R4123 vdd.n3663 vdd.n3662 0.0705758
R4124 vdd.n3680 vdd.n1962 0.0705758
R4125 vdd.n3706 vdd.n1945 0.0705758
R4126 vdd.n3733 vdd.n1933 0.0705758
R4127 vdd.n3752 vdd.n1922 0.0705758
R4128 vdd.n3771 vdd.n1911 0.0705758
R4129 vdd.n3790 vdd.n1900 0.0705758
R4130 vdd.n3809 vdd.n1889 0.0705758
R4131 vdd.n2716 vdd.n2526 0.0651067
R4132 vdd.n2716 vdd.n2715 0.0651067
R4133 vdd.n2711 vdd.n2710 0.0651067
R4134 vdd.n2710 vdd.n2530 0.0651067
R4135 vdd.n2702 vdd.n2701 0.0651067
R4136 vdd.n2724 vdd.n2516 0.0651067
R4137 vdd.n925 vdd 0.0619615
R4138 vdd.n1176 vdd 0.0619615
R4139 vdd.n1427 vdd 0.0619615
R4140 vdd vdd.n1684 0.0619615
R4141 vdd.n3042 vdd 0.0619615
R4142 vdd.n3268 vdd 0.0619615
R4143 vdd.n3494 vdd 0.0619615
R4144 vdd vdd.n3716 0.0619615
R4145 vdd.n2610 vdd.n2571 0.061744
R4146 vdd.n2614 vdd.n2611 0.061744
R4147 vdd.n2650 vdd.n2649 0.061744
R4148 vdd.n2633 vdd.n2563 0.061744
R4149 vdd.n2637 vdd.n2626 0.061744
R4150 vdd.n2642 vdd.n2641 0.061744
R4151 vdd.n2641 vdd.n2628 0.061744
R4152 vdd.n2661 vdd.n2556 0.061744
R4153 vdd.n2663 vdd.n2662 0.061744
R4154 vdd.n2673 vdd.n2554 0.061744
R4155 vdd.n2669 vdd.n2668 0.061744
R4156 vdd.n2668 vdd.n2550 0.061744
R4157 vdd.n2683 vdd.n2680 0.061744
R4158 vdd.n1805 vdd.n1803 0.0616979
R4159 vdd.n2797 vdd.n2787 0.0616979
R4160 vdd vdd.n1805 0.0603958
R4161 vdd.n2787 vdd 0.0603958
R4162 vdd.n1803 vdd.n1792 0.0590938
R4163 vdd.n2797 vdd.n2796 0.0590938
R4164 vdd.n1859 vdd 0.0579444
R4165 vdd.n3824 vdd 0.0579444
R4166 vdd.n1836 vdd.n1787 0.0577917
R4167 vdd.n2771 vdd.n2765 0.0577917
R4168 vdd.n717 vdd.n716 0.0573182
R4169 vdd.n734 vdd.n732 0.0573182
R4170 vdd.n757 vdd.n756 0.0573182
R4171 vdd.n771 vdd.n769 0.0573182
R4172 vdd.n796 vdd.n795 0.0573182
R4173 vdd.n834 vdd.n832 0.0573182
R4174 vdd.n849 vdd.n520 0.0573182
R4175 vdd.n874 vdd.n873 0.0573182
R4176 vdd.n896 vdd.n895 0.0573182
R4177 vdd.n908 vdd.n485 0.0573182
R4178 vdd.n968 vdd.n967 0.0573182
R4179 vdd.n985 vdd.n983 0.0573182
R4180 vdd.n1008 vdd.n1007 0.0573182
R4181 vdd.n1022 vdd.n1020 0.0573182
R4182 vdd.n1047 vdd.n1046 0.0573182
R4183 vdd.n1085 vdd.n1083 0.0573182
R4184 vdd.n1100 vdd.n386 0.0573182
R4185 vdd.n1125 vdd.n1124 0.0573182
R4186 vdd.n1147 vdd.n1146 0.0573182
R4187 vdd.n1159 vdd.n351 0.0573182
R4188 vdd.n1219 vdd.n1218 0.0573182
R4189 vdd.n1236 vdd.n1234 0.0573182
R4190 vdd.n1259 vdd.n1258 0.0573182
R4191 vdd.n1273 vdd.n1271 0.0573182
R4192 vdd.n1298 vdd.n1297 0.0573182
R4193 vdd.n1336 vdd.n1334 0.0573182
R4194 vdd.n1351 vdd.n252 0.0573182
R4195 vdd.n1376 vdd.n1375 0.0573182
R4196 vdd.n1398 vdd.n1397 0.0573182
R4197 vdd.n1410 vdd.n217 0.0573182
R4198 vdd.n1470 vdd.n1469 0.0573182
R4199 vdd.n1487 vdd.n1485 0.0573182
R4200 vdd.n1510 vdd.n1509 0.0573182
R4201 vdd.n1524 vdd.n1522 0.0573182
R4202 vdd.n1549 vdd.n1548 0.0573182
R4203 vdd.n1582 vdd.n1581 0.0573182
R4204 vdd.n1605 vdd.n1604 0.0573182
R4205 vdd.n1621 vdd.n108 0.0573182
R4206 vdd.n1638 vdd.n101 0.0573182
R4207 vdd.n1667 vdd.n1665 0.0573182
R4208 vdd.n1697 vdd.n1696 0.0573182
R4209 vdd.n1720 vdd.n1719 0.0573182
R4210 vdd.n1736 vdd.n44 0.0573182
R4211 vdd.n1753 vdd.n37 0.0573182
R4212 vdd.n1777 vdd.n1776 0.0573182
R4213 vdd.n2841 vdd.n2839 0.0573182
R4214 vdd.n2861 vdd.n2860 0.0573182
R4215 vdd.n2875 vdd.n2873 0.0573182
R4216 vdd.n2896 vdd.n2895 0.0573182
R4217 vdd.n2916 vdd.n2915 0.0573182
R4218 vdd.n2951 vdd.n2950 0.0573182
R4219 vdd.n2969 vdd.n2379 0.0573182
R4220 vdd.n2983 vdd.n2373 0.0573182
R4221 vdd.n3000 vdd.n2366 0.0573182
R4222 vdd.n3022 vdd.n3021 0.0573182
R4223 vdd.n3067 vdd.n3065 0.0573182
R4224 vdd.n3087 vdd.n3086 0.0573182
R4225 vdd.n3101 vdd.n3099 0.0573182
R4226 vdd.n3122 vdd.n3121 0.0573182
R4227 vdd.n3142 vdd.n3141 0.0573182
R4228 vdd.n3177 vdd.n3176 0.0573182
R4229 vdd.n3195 vdd.n2245 0.0573182
R4230 vdd.n3209 vdd.n2239 0.0573182
R4231 vdd.n3226 vdd.n2232 0.0573182
R4232 vdd.n3248 vdd.n3247 0.0573182
R4233 vdd.n3293 vdd.n3291 0.0573182
R4234 vdd.n3313 vdd.n3312 0.0573182
R4235 vdd.n3327 vdd.n3325 0.0573182
R4236 vdd.n3348 vdd.n3347 0.0573182
R4237 vdd.n3368 vdd.n3367 0.0573182
R4238 vdd.n3403 vdd.n3402 0.0573182
R4239 vdd.n3421 vdd.n2111 0.0573182
R4240 vdd.n3435 vdd.n2105 0.0573182
R4241 vdd.n3452 vdd.n2098 0.0573182
R4242 vdd.n3474 vdd.n3473 0.0573182
R4243 vdd.n3519 vdd.n3517 0.0573182
R4244 vdd.n3539 vdd.n3538 0.0573182
R4245 vdd.n3553 vdd.n3551 0.0573182
R4246 vdd.n3574 vdd.n3573 0.0573182
R4247 vdd.n3594 vdd.n3593 0.0573182
R4248 vdd.n3629 vdd.n3628 0.0573182
R4249 vdd.n3647 vdd.n1977 0.0573182
R4250 vdd.n3661 vdd.n1971 0.0573182
R4251 vdd.n3678 vdd.n1964 0.0573182
R4252 vdd.n3705 vdd.n3703 0.0573182
R4253 vdd.n3732 vdd.n3731 0.0573182
R4254 vdd.n3751 vdd.n3750 0.0573182
R4255 vdd.n3770 vdd.n3769 0.0573182
R4256 vdd.n3789 vdd.n3788 0.0573182
R4257 vdd.n3808 vdd.n3807 0.0573182
R4258 vdd.n674 vdd.n665 0.0563252
R4259 vdd.n2560 vdd.n2559 0.0532517
R4260 vdd.n1809 vdd.n1 0.0517727
R4261 vdd.n2767 vdd.n1871 0.0517727
R4262 vdd.n1864 vdd.n3 0.0455
R4263 vdd.n3829 vdd.n1873 0.0455
R4264 vdd.n2689 vdd.n2688 0.0443776
R4265 vdd.n1798 vdd.n1797 0.0438377
R4266 vdd.n2786 vdd.n2783 0.0438377
R4267 vdd.n1686 vdd.n68 0.0434423
R4268 vdd.n3722 vdd.n1933 0.0434103
R4269 vdd.n2629 vdd.n2561 0.0424742
R4270 vdd.n2638 vdd.n2630 0.0424742
R4271 vdd.n2640 vdd.n2639 0.0424742
R4272 vdd.n2660 vdd.n2555 0.0424742
R4273 vdd.n2672 vdd.n2664 0.0424742
R4274 vdd.n2671 vdd.n2670 0.0424742
R4275 vdd.n2665 vdd.n2548 0.0424742
R4276 vdd.n1815 vdd.n1814 0.041625
R4277 vdd.n2768 vdd.n2764 0.041625
R4278 vdd.n1787 vdd 0.0408646
R4279 vdd vdd.n2771 0.0408646
R4280 vdd.n599 vdd.n593 0.0402727
R4281 vdd.n744 vdd.n584 0.0402727
R4282 vdd.n774 vdd.n568 0.0402727
R4283 vdd.n783 vdd.n561 0.0402727
R4284 vdd.n808 vdd.n547 0.0402727
R4285 vdd.n819 vdd.n533 0.0402727
R4286 vdd.n847 vdd.n846 0.0402727
R4287 vdd.n519 vdd.n511 0.0402727
R4288 vdd.n883 vdd.n498 0.0402727
R4289 vdd.n906 vdd.n905 0.0402727
R4290 vdd.n914 vdd.n479 0.0402727
R4291 vdd.n952 vdd.n473 0.0402727
R4292 vdd.n465 vdd.n459 0.0402727
R4293 vdd.n995 vdd.n450 0.0402727
R4294 vdd.n1025 vdd.n434 0.0402727
R4295 vdd.n1034 vdd.n427 0.0402727
R4296 vdd.n1059 vdd.n413 0.0402727
R4297 vdd.n1070 vdd.n399 0.0402727
R4298 vdd.n1098 vdd.n1097 0.0402727
R4299 vdd.n385 vdd.n377 0.0402727
R4300 vdd.n1134 vdd.n364 0.0402727
R4301 vdd.n1157 vdd.n1156 0.0402727
R4302 vdd.n1165 vdd.n345 0.0402727
R4303 vdd.n1203 vdd.n339 0.0402727
R4304 vdd.n331 vdd.n325 0.0402727
R4305 vdd.n1246 vdd.n316 0.0402727
R4306 vdd.n1276 vdd.n300 0.0402727
R4307 vdd.n1285 vdd.n293 0.0402727
R4308 vdd.n1310 vdd.n279 0.0402727
R4309 vdd.n1321 vdd.n265 0.0402727
R4310 vdd.n1349 vdd.n1348 0.0402727
R4311 vdd.n251 vdd.n243 0.0402727
R4312 vdd.n1385 vdd.n230 0.0402727
R4313 vdd.n1408 vdd.n1407 0.0402727
R4314 vdd.n1416 vdd.n211 0.0402727
R4315 vdd.n1454 vdd.n205 0.0402727
R4316 vdd.n197 vdd.n191 0.0402727
R4317 vdd.n1497 vdd.n182 0.0402727
R4318 vdd.n1527 vdd.n166 0.0402727
R4319 vdd.n1536 vdd.n159 0.0402727
R4320 vdd.n1561 vdd.n145 0.0402727
R4321 vdd.n1572 vdd.n132 0.0402727
R4322 vdd.n1594 vdd.n126 0.0402727
R4323 vdd.n1623 vdd.n109 0.0402727
R4324 vdd.n1641 vdd.n1640 0.0402727
R4325 vdd.n1652 vdd.n83 0.0402727
R4326 vdd.n717 vdd.n600 0.0402727
R4327 vdd.n732 vdd.n590 0.0402727
R4328 vdd.n756 vdd.n577 0.0402727
R4329 vdd.n772 vdd.n771 0.0402727
R4330 vdd.n796 vdd.n554 0.0402727
R4331 vdd.n812 vdd.n810 0.0402727
R4332 vdd.n811 vdd.n539 0.0402727
R4333 vdd.n834 vdd.n833 0.0402727
R4334 vdd.n858 vdd.n520 0.0402727
R4335 vdd.n873 vdd.n505 0.0402727
R4336 vdd.n895 vdd.n493 0.0402727
R4337 vdd.n931 vdd.n485 0.0402727
R4338 vdd.n968 vdd.n466 0.0402727
R4339 vdd.n983 vdd.n456 0.0402727
R4340 vdd.n1007 vdd.n443 0.0402727
R4341 vdd.n1023 vdd.n1022 0.0402727
R4342 vdd.n1047 vdd.n420 0.0402727
R4343 vdd.n1063 vdd.n1061 0.0402727
R4344 vdd.n1062 vdd.n405 0.0402727
R4345 vdd.n1085 vdd.n1084 0.0402727
R4346 vdd.n1109 vdd.n386 0.0402727
R4347 vdd.n1124 vdd.n371 0.0402727
R4348 vdd.n1146 vdd.n359 0.0402727
R4349 vdd.n1182 vdd.n351 0.0402727
R4350 vdd.n1219 vdd.n332 0.0402727
R4351 vdd.n1234 vdd.n322 0.0402727
R4352 vdd.n1258 vdd.n309 0.0402727
R4353 vdd.n1274 vdd.n1273 0.0402727
R4354 vdd.n1298 vdd.n286 0.0402727
R4355 vdd.n1314 vdd.n1312 0.0402727
R4356 vdd.n1313 vdd.n271 0.0402727
R4357 vdd.n1336 vdd.n1335 0.0402727
R4358 vdd.n1360 vdd.n252 0.0402727
R4359 vdd.n1375 vdd.n237 0.0402727
R4360 vdd.n1397 vdd.n225 0.0402727
R4361 vdd.n1433 vdd.n217 0.0402727
R4362 vdd.n1470 vdd.n198 0.0402727
R4363 vdd.n1485 vdd.n188 0.0402727
R4364 vdd.n1509 vdd.n175 0.0402727
R4365 vdd.n1525 vdd.n1524 0.0402727
R4366 vdd.n1549 vdd.n152 0.0402727
R4367 vdd.n1565 vdd.n1563 0.0402727
R4368 vdd.n1564 vdd.n137 0.0402727
R4369 vdd.n1582 vdd.n123 0.0402727
R4370 vdd.n1606 vdd.n1605 0.0402727
R4371 vdd.n1621 vdd.n1620 0.0402727
R4372 vdd.n101 vdd.n89 0.0402727
R4373 vdd.n1667 vdd.n1666 0.0402727
R4374 vdd.n1709 vdd.n62 0.0402727
R4375 vdd.n1738 vdd.n45 0.0402727
R4376 vdd.n1756 vdd.n1755 0.0402727
R4377 vdd.n1767 vdd.n20 0.0402727
R4378 vdd.n1852 vdd.n12 0.0402727
R4379 vdd.n1697 vdd.n59 0.0402727
R4380 vdd.n1721 vdd.n1720 0.0402727
R4381 vdd.n1736 vdd.n1735 0.0402727
R4382 vdd.n37 vdd.n25 0.0402727
R4383 vdd.n1777 vdd.n9 0.0402727
R4384 vdd.n2851 vdd.n2454 0.0402727
R4385 vdd.n2878 vdd.n2440 0.0402727
R4386 vdd.n2886 vdd.n2435 0.0402727
R4387 vdd.n2906 vdd.n2424 0.0402727
R4388 vdd.n2925 vdd.n2403 0.0402727
R4389 vdd.n2936 vdd.n2388 0.0402727
R4390 vdd.n2967 vdd.n2380 0.0402727
R4391 vdd.n2985 vdd.n2374 0.0402727
R4392 vdd.n3003 vdd.n3002 0.0402727
R4393 vdd.n3012 vdd.n2348 0.0402727
R4394 vdd.n3036 vdd.n2343 0.0402727
R4395 vdd.n3056 vdd.n2331 0.0402727
R4396 vdd.n3077 vdd.n2320 0.0402727
R4397 vdd.n3104 vdd.n2306 0.0402727
R4398 vdd.n3112 vdd.n2301 0.0402727
R4399 vdd.n3132 vdd.n2290 0.0402727
R4400 vdd.n3151 vdd.n2269 0.0402727
R4401 vdd.n3162 vdd.n2254 0.0402727
R4402 vdd.n3193 vdd.n2246 0.0402727
R4403 vdd.n3211 vdd.n2240 0.0402727
R4404 vdd.n3229 vdd.n3228 0.0402727
R4405 vdd.n3238 vdd.n2214 0.0402727
R4406 vdd.n3262 vdd.n2209 0.0402727
R4407 vdd.n3282 vdd.n2197 0.0402727
R4408 vdd.n3303 vdd.n2186 0.0402727
R4409 vdd.n3330 vdd.n2172 0.0402727
R4410 vdd.n3338 vdd.n2167 0.0402727
R4411 vdd.n3358 vdd.n2156 0.0402727
R4412 vdd.n3377 vdd.n2135 0.0402727
R4413 vdd.n3388 vdd.n2120 0.0402727
R4414 vdd.n3419 vdd.n2112 0.0402727
R4415 vdd.n3437 vdd.n2106 0.0402727
R4416 vdd.n3455 vdd.n3454 0.0402727
R4417 vdd.n3464 vdd.n2080 0.0402727
R4418 vdd.n3488 vdd.n2075 0.0402727
R4419 vdd.n3508 vdd.n2063 0.0402727
R4420 vdd.n3529 vdd.n2052 0.0402727
R4421 vdd.n3556 vdd.n2038 0.0402727
R4422 vdd.n3564 vdd.n2033 0.0402727
R4423 vdd.n3584 vdd.n2022 0.0402727
R4424 vdd.n3603 vdd.n2001 0.0402727
R4425 vdd.n3614 vdd.n1986 0.0402727
R4426 vdd.n3645 vdd.n1978 0.0402727
R4427 vdd.n3663 vdd.n1972 0.0402727
R4428 vdd.n3681 vdd.n3680 0.0402727
R4429 vdd.n3690 vdd.n1945 0.0402727
R4430 vdd.n2839 vdd.n2460 0.0402727
R4431 vdd.n2860 vdd.n2449 0.0402727
R4432 vdd.n2876 vdd.n2875 0.0402727
R4433 vdd.n2896 vdd.n2429 0.0402727
R4434 vdd.n2916 vdd.n2418 0.0402727
R4435 vdd.n2410 vdd.n2402 0.0402727
R4436 vdd.n2409 vdd.n2396 0.0402727
R4437 vdd.n2950 vdd.n2387 0.0402727
R4438 vdd.n2970 vdd.n2969 0.0402727
R4439 vdd.n2983 vdd.n2982 0.0402727
R4440 vdd.n2366 vdd.n2353 0.0402727
R4441 vdd.n3022 vdd.n2340 0.0402727
R4442 vdd.n3065 vdd.n2326 0.0402727
R4443 vdd.n3086 vdd.n2315 0.0402727
R4444 vdd.n3102 vdd.n3101 0.0402727
R4445 vdd.n3122 vdd.n2295 0.0402727
R4446 vdd.n3142 vdd.n2284 0.0402727
R4447 vdd.n2276 vdd.n2268 0.0402727
R4448 vdd.n2275 vdd.n2262 0.0402727
R4449 vdd.n3176 vdd.n2253 0.0402727
R4450 vdd.n3196 vdd.n3195 0.0402727
R4451 vdd.n3209 vdd.n3208 0.0402727
R4452 vdd.n2232 vdd.n2219 0.0402727
R4453 vdd.n3248 vdd.n2206 0.0402727
R4454 vdd.n3291 vdd.n2192 0.0402727
R4455 vdd.n3312 vdd.n2181 0.0402727
R4456 vdd.n3328 vdd.n3327 0.0402727
R4457 vdd.n3348 vdd.n2161 0.0402727
R4458 vdd.n3368 vdd.n2150 0.0402727
R4459 vdd.n2142 vdd.n2134 0.0402727
R4460 vdd.n2141 vdd.n2128 0.0402727
R4461 vdd.n3402 vdd.n2119 0.0402727
R4462 vdd.n3422 vdd.n3421 0.0402727
R4463 vdd.n3435 vdd.n3434 0.0402727
R4464 vdd.n2098 vdd.n2085 0.0402727
R4465 vdd.n3474 vdd.n2072 0.0402727
R4466 vdd.n3517 vdd.n2058 0.0402727
R4467 vdd.n3538 vdd.n2047 0.0402727
R4468 vdd.n3554 vdd.n3553 0.0402727
R4469 vdd.n3574 vdd.n2027 0.0402727
R4470 vdd.n3594 vdd.n2016 0.0402727
R4471 vdd.n2008 vdd.n2000 0.0402727
R4472 vdd.n2007 vdd.n1994 0.0402727
R4473 vdd.n3628 vdd.n1985 0.0402727
R4474 vdd.n3648 vdd.n3647 0.0402727
R4475 vdd.n3661 vdd.n3660 0.0402727
R4476 vdd.n1964 vdd.n1951 0.0402727
R4477 vdd.n3705 vdd.n3704 0.0402727
R4478 vdd.n3741 vdd.n1922 0.0402727
R4479 vdd.n3760 vdd.n1911 0.0402727
R4480 vdd.n3779 vdd.n1900 0.0402727
R4481 vdd.n3798 vdd.n1889 0.0402727
R4482 vdd.n3817 vdd.n1882 0.0402727
R4483 vdd.n3732 vdd.n1927 0.0402727
R4484 vdd.n3751 vdd.n1916 0.0402727
R4485 vdd.n3770 vdd.n1905 0.0402727
R4486 vdd.n3789 vdd.n1894 0.0402727
R4487 vdd.n3808 vdd.n1879 0.0402727
R4488 vdd.n2725 vdd.n2515 0.0391236
R4489 vdd.n2658 vdd.n2557 0.0378616
R4490 vdd.n2715 vdd.n2527 0.0377191
R4491 vdd.n607 vdd.n606 0.0364848
R4492 vdd.n713 vdd.n601 0.0364848
R4493 vdd.n733 vdd.n585 0.0364848
R4494 vdd.n759 vdd.n758 0.0364848
R4495 vdd.n572 vdd.n560 0.0364848
R4496 vdd.n555 vdd.n545 0.0364848
R4497 vdd.n540 vdd.n534 0.0364848
R4498 vdd.n848 vdd.n525 0.0364848
R4499 vdd.n521 vdd.n510 0.0364848
R4500 vdd.n506 vdd.n497 0.0364848
R4501 vdd.n907 vdd.n491 0.0364848
R4502 vdd.n915 vdd.n486 0.0364848
R4503 vdd.n917 vdd.n472 0.0364848
R4504 vdd.n964 vdd.n467 0.0364848
R4505 vdd.n984 vdd.n451 0.0364848
R4506 vdd.n1010 vdd.n1009 0.0364848
R4507 vdd.n438 vdd.n426 0.0364848
R4508 vdd.n421 vdd.n411 0.0364848
R4509 vdd.n406 vdd.n400 0.0364848
R4510 vdd.n1099 vdd.n391 0.0364848
R4511 vdd.n387 vdd.n376 0.0364848
R4512 vdd.n372 vdd.n363 0.0364848
R4513 vdd.n1158 vdd.n357 0.0364848
R4514 vdd.n1166 vdd.n352 0.0364848
R4515 vdd.n1168 vdd.n338 0.0364848
R4516 vdd.n1215 vdd.n333 0.0364848
R4517 vdd.n1235 vdd.n317 0.0364848
R4518 vdd.n1261 vdd.n1260 0.0364848
R4519 vdd.n304 vdd.n292 0.0364848
R4520 vdd.n287 vdd.n277 0.0364848
R4521 vdd.n272 vdd.n266 0.0364848
R4522 vdd.n1350 vdd.n257 0.0364848
R4523 vdd.n253 vdd.n242 0.0364848
R4524 vdd.n238 vdd.n229 0.0364848
R4525 vdd.n1409 vdd.n223 0.0364848
R4526 vdd.n1417 vdd.n218 0.0364848
R4527 vdd.n1419 vdd.n204 0.0364848
R4528 vdd.n1466 vdd.n199 0.0364848
R4529 vdd.n1486 vdd.n183 0.0364848
R4530 vdd.n1512 vdd.n1511 0.0364848
R4531 vdd.n170 vdd.n158 0.0364848
R4532 vdd.n153 vdd.n143 0.0364848
R4533 vdd.n138 vdd.n133 0.0364848
R4534 vdd.n124 vdd.n117 0.0364848
R4535 vdd.n1625 vdd.n1624 0.0364848
R4536 vdd.n1639 vdd.n100 0.0364848
R4537 vdd.n90 vdd.n84 0.0364848
R4538 vdd.n1682 vdd.n73 0.0364848
R4539 vdd.n1687 vdd.n69 0.0364848
R4540 vdd.n60 vdd.n53 0.0364848
R4541 vdd.n1740 vdd.n1739 0.0364848
R4542 vdd.n1754 vdd.n36 0.0364848
R4543 vdd.n26 vdd.n21 0.0364848
R4544 vdd.n10 vdd.n5 0.0364848
R4545 vdd.n2464 vdd.n2463 0.0364848
R4546 vdd.n2840 vdd.n2455 0.0364848
R4547 vdd.n2863 vdd.n2862 0.0364848
R4548 vdd.n2444 vdd.n2434 0.0364848
R4549 vdd.n2430 vdd.n2423 0.0364848
R4550 vdd.n2419 vdd.n2401 0.0364848
R4551 vdd.n2397 vdd.n2386 0.0364848
R4552 vdd.n2966 vdd.n2965 0.0364848
R4553 vdd.n2987 vdd.n2986 0.0364848
R4554 vdd.n3001 vdd.n2365 0.0364848
R4555 vdd.n2354 vdd.n2349 0.0364848
R4556 vdd.n2341 vdd.n2336 0.0364848
R4557 vdd.n3046 vdd.n2332 0.0364848
R4558 vdd.n3066 vdd.n2321 0.0364848
R4559 vdd.n3089 vdd.n3088 0.0364848
R4560 vdd.n2310 vdd.n2300 0.0364848
R4561 vdd.n2296 vdd.n2289 0.0364848
R4562 vdd.n2285 vdd.n2267 0.0364848
R4563 vdd.n2263 vdd.n2252 0.0364848
R4564 vdd.n3192 vdd.n3191 0.0364848
R4565 vdd.n3213 vdd.n3212 0.0364848
R4566 vdd.n3227 vdd.n2231 0.0364848
R4567 vdd.n2220 vdd.n2215 0.0364848
R4568 vdd.n2207 vdd.n2202 0.0364848
R4569 vdd.n3272 vdd.n2198 0.0364848
R4570 vdd.n3292 vdd.n2187 0.0364848
R4571 vdd.n3315 vdd.n3314 0.0364848
R4572 vdd.n2176 vdd.n2166 0.0364848
R4573 vdd.n2162 vdd.n2155 0.0364848
R4574 vdd.n2151 vdd.n2133 0.0364848
R4575 vdd.n2129 vdd.n2118 0.0364848
R4576 vdd.n3418 vdd.n3417 0.0364848
R4577 vdd.n3439 vdd.n3438 0.0364848
R4578 vdd.n3453 vdd.n2097 0.0364848
R4579 vdd.n2086 vdd.n2081 0.0364848
R4580 vdd.n2073 vdd.n2068 0.0364848
R4581 vdd.n3498 vdd.n2064 0.0364848
R4582 vdd.n3518 vdd.n2053 0.0364848
R4583 vdd.n3541 vdd.n3540 0.0364848
R4584 vdd.n2042 vdd.n2032 0.0364848
R4585 vdd.n2028 vdd.n2021 0.0364848
R4586 vdd.n2017 vdd.n1999 0.0364848
R4587 vdd.n1995 vdd.n1984 0.0364848
R4588 vdd.n3644 vdd.n3643 0.0364848
R4589 vdd.n3665 vdd.n3664 0.0364848
R4590 vdd.n3679 vdd.n1963 0.0364848
R4591 vdd.n1952 vdd.n1946 0.0364848
R4592 vdd.n3714 vdd.n1938 0.0364848
R4593 vdd.n3718 vdd.n1934 0.0364848
R4594 vdd.n1928 vdd.n1923 0.0364848
R4595 vdd.n1917 vdd.n1912 0.0364848
R4596 vdd.n1906 vdd.n1901 0.0364848
R4597 vdd.n1895 vdd.n1890 0.0364848
R4598 vdd.n1880 vdd.n1875 0.0364848
R4599 vdd.n2694 vdd.n2693 0.0353392
R4600 vdd.n1795 vdd.n1794 0.0351948
R4601 vdd.n2785 vdd.n2784 0.0351948
R4602 vdd.n2699 vdd.n2530 0.0349101
R4603 vdd.n2542 vdd.n2541 0.0336958
R4604 vdd vdd.n2526 0.0335056
R4605 vdd.n2702 vdd 0.0328034
R4606 vdd.n1819 vdd.n1818 0.0309054
R4607 vdd.n2803 vdd.n2763 0.0309054
R4608 vdd.n719 vdd.n598 0.030803
R4609 vdd.n730 vdd.n591 0.030803
R4610 vdd.n754 vdd.n578 0.030803
R4611 vdd.n773 vdd.n571 0.030803
R4612 vdd.n798 vdd.n553 0.030803
R4613 vdd.n814 vdd.n543 0.030803
R4614 vdd.n818 vdd.n541 0.030803
R4615 vdd.n836 vdd.n526 0.030803
R4616 vdd.n860 vdd.n859 0.030803
R4617 vdd.n871 vdd.n504 0.030803
R4618 vdd.n893 vdd.n492 0.030803
R4619 vdd.n933 vdd.n932 0.030803
R4620 vdd.n970 vdd.n464 0.030803
R4621 vdd.n981 vdd.n457 0.030803
R4622 vdd.n1005 vdd.n444 0.030803
R4623 vdd.n1024 vdd.n437 0.030803
R4624 vdd.n1049 vdd.n419 0.030803
R4625 vdd.n1065 vdd.n409 0.030803
R4626 vdd.n1069 vdd.n407 0.030803
R4627 vdd.n1087 vdd.n392 0.030803
R4628 vdd.n1111 vdd.n1110 0.030803
R4629 vdd.n1122 vdd.n370 0.030803
R4630 vdd.n1144 vdd.n358 0.030803
R4631 vdd.n1184 vdd.n1183 0.030803
R4632 vdd.n1221 vdd.n330 0.030803
R4633 vdd.n1232 vdd.n323 0.030803
R4634 vdd.n1256 vdd.n310 0.030803
R4635 vdd.n1275 vdd.n303 0.030803
R4636 vdd.n1300 vdd.n285 0.030803
R4637 vdd.n1316 vdd.n275 0.030803
R4638 vdd.n1320 vdd.n273 0.030803
R4639 vdd.n1338 vdd.n258 0.030803
R4640 vdd.n1362 vdd.n1361 0.030803
R4641 vdd.n1373 vdd.n236 0.030803
R4642 vdd.n1395 vdd.n224 0.030803
R4643 vdd.n1435 vdd.n1434 0.030803
R4644 vdd.n1472 vdd.n196 0.030803
R4645 vdd.n1483 vdd.n189 0.030803
R4646 vdd.n1507 vdd.n176 0.030803
R4647 vdd.n1526 vdd.n169 0.030803
R4648 vdd.n1551 vdd.n151 0.030803
R4649 vdd.n1567 vdd.n141 0.030803
R4650 vdd.n1571 vdd.n139 0.030803
R4651 vdd.n1584 vdd.n125 0.030803
R4652 vdd.n1608 vdd.n1607 0.030803
R4653 vdd.n1619 vdd.n97 0.030803
R4654 vdd.n1651 vdd.n91 0.030803
R4655 vdd.n1669 vdd.n74 0.030803
R4656 vdd.n1699 vdd.n61 0.030803
R4657 vdd.n1723 vdd.n1722 0.030803
R4658 vdd.n1734 vdd.n33 0.030803
R4659 vdd.n1766 vdd.n27 0.030803
R4660 vdd.n1779 vdd.n11 0.030803
R4661 vdd.n2837 vdd.n2461 0.030803
R4662 vdd.n2858 vdd.n2450 0.030803
R4663 vdd.n2877 vdd.n2443 0.030803
R4664 vdd.n2898 vdd.n2428 0.030803
R4665 vdd.n2918 vdd.n2417 0.030803
R4666 vdd.n2412 vdd.n2404 0.030803
R4667 vdd.n2407 vdd.n2395 0.030803
R4668 vdd.n2948 vdd.n2389 0.030803
R4669 vdd.n2971 vdd.n2378 0.030803
R4670 vdd.n2981 vdd.n2360 0.030803
R4671 vdd.n2363 vdd.n2355 0.030803
R4672 vdd.n3024 vdd.n2342 0.030803
R4673 vdd.n3063 vdd.n2327 0.030803
R4674 vdd.n3084 vdd.n2316 0.030803
R4675 vdd.n3103 vdd.n2309 0.030803
R4676 vdd.n3124 vdd.n2294 0.030803
R4677 vdd.n3144 vdd.n2283 0.030803
R4678 vdd.n2278 vdd.n2270 0.030803
R4679 vdd.n2273 vdd.n2261 0.030803
R4680 vdd.n3174 vdd.n2255 0.030803
R4681 vdd.n3197 vdd.n2244 0.030803
R4682 vdd.n3207 vdd.n2226 0.030803
R4683 vdd.n2229 vdd.n2221 0.030803
R4684 vdd.n3250 vdd.n2208 0.030803
R4685 vdd.n3289 vdd.n2193 0.030803
R4686 vdd.n3310 vdd.n2182 0.030803
R4687 vdd.n3329 vdd.n2175 0.030803
R4688 vdd.n3350 vdd.n2160 0.030803
R4689 vdd.n3370 vdd.n2149 0.030803
R4690 vdd.n2144 vdd.n2136 0.030803
R4691 vdd.n2139 vdd.n2127 0.030803
R4692 vdd.n3400 vdd.n2121 0.030803
R4693 vdd.n3423 vdd.n2110 0.030803
R4694 vdd.n3433 vdd.n2092 0.030803
R4695 vdd.n2095 vdd.n2087 0.030803
R4696 vdd.n3476 vdd.n2074 0.030803
R4697 vdd.n3515 vdd.n2059 0.030803
R4698 vdd.n3536 vdd.n2048 0.030803
R4699 vdd.n3555 vdd.n2041 0.030803
R4700 vdd.n3576 vdd.n2026 0.030803
R4701 vdd.n3596 vdd.n2015 0.030803
R4702 vdd.n2010 vdd.n2002 0.030803
R4703 vdd.n2005 vdd.n1993 0.030803
R4704 vdd.n3626 vdd.n1987 0.030803
R4705 vdd.n3649 vdd.n1976 0.030803
R4706 vdd.n3659 vdd.n1958 0.030803
R4707 vdd.n1961 vdd.n1953 0.030803
R4708 vdd.n3707 vdd.n1939 0.030803
R4709 vdd.n3734 vdd.n1929 0.030803
R4710 vdd.n3753 vdd.n1918 0.030803
R4711 vdd.n3772 vdd.n1907 0.030803
R4712 vdd.n3791 vdd.n1896 0.030803
R4713 vdd.n3810 vdd.n1881 0.030803
R4714 vdd.n2701 vdd.n2699 0.0306966
R4715 vdd.n1808 vdd.n1807 0.0292162
R4716 vdd.n2778 vdd.n2762 0.0292162
R4717 vdd.n2747 vdd.n2746 0.0282727
R4718 vdd.n2711 vdd.n2527 0.0278876
R4719 vdd.n1806 vdd 0.0265417
R4720 vdd vdd.n2761 0.0265417
R4721 vdd.n2725 vdd.n2724 0.0264831
R4722 vdd.n692 vdd.n610 0.0242893
R4723 vdd.n643 vdd.n642 0.0242893
R4724 vdd.n636 vdd.n631 0.0242893
R4725 vdd.n632 vdd.n627 0.0242893
R4726 vdd.n621 vdd.n620 0.0242893
R4727 vdd.n2751 vdd.n2509 0.0242893
R4728 vdd.n2814 vdd.n2470 0.0242893
R4729 vdd.n2504 vdd.n2471 0.0242893
R4730 vdd.n2486 vdd.n2476 0.0242893
R4731 vdd.n2492 vdd.n2480 0.0242893
R4732 vdd.n1820 vdd.n1806 0.0239375
R4733 vdd.n2804 vdd.n2761 0.0239375
R4734 vdd.n657 vdd.n656 0.0234759
R4735 vdd.n2736 vdd.n2735 0.0234759
R4736 vdd.n1792 vdd 0.0226354
R4737 vdd.n2796 vdd 0.0226354
R4738 vdd.n2729 vdd.n2728 0.0213706
R4739 vdd.n1861 vdd.n4 0.0206084
R4740 vdd.n3826 vdd.n1874 0.0206084
R4741 vdd.n704 vdd.n703 0.0205441
R4742 vdd.n711 vdd.n710 0.0205441
R4743 vdd.n742 vdd.n741 0.0205441
R4744 vdd.n763 vdd.n762 0.0205441
R4745 vdd.n786 vdd.n785 0.0205441
R4746 vdd.n789 vdd.n546 0.0205441
R4747 vdd.n955 vdd.n954 0.0205441
R4748 vdd.n962 vdd.n961 0.0205441
R4749 vdd.n993 vdd.n992 0.0205441
R4750 vdd.n1014 vdd.n1013 0.0205441
R4751 vdd.n1037 vdd.n1036 0.0205441
R4752 vdd.n1040 vdd.n412 0.0205441
R4753 vdd.n1206 vdd.n1205 0.0205441
R4754 vdd.n1213 vdd.n1212 0.0205441
R4755 vdd.n1244 vdd.n1243 0.0205441
R4756 vdd.n1265 vdd.n1264 0.0205441
R4757 vdd.n1288 vdd.n1287 0.0205441
R4758 vdd.n1291 vdd.n278 0.0205441
R4759 vdd.n1457 vdd.n1456 0.0205441
R4760 vdd.n1464 vdd.n1463 0.0205441
R4761 vdd.n1495 vdd.n1494 0.0205441
R4762 vdd.n1516 vdd.n1515 0.0205441
R4763 vdd.n1539 vdd.n1538 0.0205441
R4764 vdd.n1542 vdd.n144 0.0205441
R4765 vdd.n2828 vdd.n2827 0.0205441
R4766 vdd.n2849 vdd.n2848 0.0205441
R4767 vdd.n2867 vdd.n2866 0.0205441
R4768 vdd.n2889 vdd.n2888 0.0205441
R4769 vdd.n2909 vdd.n2908 0.0205441
R4770 vdd.n2928 vdd.n2927 0.0205441
R4771 vdd.n3054 vdd.n3053 0.0205441
R4772 vdd.n3075 vdd.n3074 0.0205441
R4773 vdd.n3093 vdd.n3092 0.0205441
R4774 vdd.n3115 vdd.n3114 0.0205441
R4775 vdd.n3135 vdd.n3134 0.0205441
R4776 vdd.n3154 vdd.n3153 0.0205441
R4777 vdd.n3280 vdd.n3279 0.0205441
R4778 vdd.n3301 vdd.n3300 0.0205441
R4779 vdd.n3319 vdd.n3318 0.0205441
R4780 vdd.n3341 vdd.n3340 0.0205441
R4781 vdd.n3361 vdd.n3360 0.0205441
R4782 vdd.n3380 vdd.n3379 0.0205441
R4783 vdd.n3506 vdd.n3505 0.0205441
R4784 vdd.n3527 vdd.n3526 0.0205441
R4785 vdd.n3545 vdd.n3544 0.0205441
R4786 vdd.n3567 vdd.n3566 0.0205441
R4787 vdd.n3587 vdd.n3586 0.0205441
R4788 vdd.n3606 vdd.n3605 0.0205441
R4789 vdd.n821 vdd.n538 0.0198529
R4790 vdd.n825 vdd.n536 0.0198529
R4791 vdd.n856 vdd.n522 0.0198529
R4792 vdd.n881 vdd.n507 0.0198529
R4793 vdd.n903 vdd.n494 0.0198529
R4794 vdd.n929 vdd.n487 0.0198529
R4795 vdd.n1072 vdd.n404 0.0198529
R4796 vdd.n1076 vdd.n402 0.0198529
R4797 vdd.n1107 vdd.n388 0.0198529
R4798 vdd.n1132 vdd.n373 0.0198529
R4799 vdd.n1154 vdd.n360 0.0198529
R4800 vdd.n1180 vdd.n353 0.0198529
R4801 vdd.n1323 vdd.n270 0.0198529
R4802 vdd.n1327 vdd.n268 0.0198529
R4803 vdd.n1358 vdd.n254 0.0198529
R4804 vdd.n1383 vdd.n239 0.0198529
R4805 vdd.n1405 vdd.n226 0.0198529
R4806 vdd.n1431 vdd.n219 0.0198529
R4807 vdd.n1574 vdd.n136 0.0198529
R4808 vdd.n1596 vdd.n122 0.0198529
R4809 vdd.n120 vdd.n119 0.0198529
R4810 vdd.n1631 vdd.n1630 0.0198529
R4811 vdd.n1654 vdd.n88 0.0198529
R4812 vdd.n1658 vdd.n86 0.0198529
R4813 vdd.n1711 vdd.n58 0.0198529
R4814 vdd.n56 vdd.n55 0.0198529
R4815 vdd.n1746 vdd.n1745 0.0198529
R4816 vdd.n1769 vdd.n24 0.0198529
R4817 vdd.n1854 vdd.n8 0.0198529
R4818 vdd.n2934 vdd.n2398 0.0198529
R4819 vdd.n2955 vdd.n2954 0.0198529
R4820 vdd.n2960 vdd.n2959 0.0198529
R4821 vdd.n2993 vdd.n2992 0.0198529
R4822 vdd.n3014 vdd.n2352 0.0198529
R4823 vdd.n3038 vdd.n2339 0.0198529
R4824 vdd.n3160 vdd.n2264 0.0198529
R4825 vdd.n3181 vdd.n3180 0.0198529
R4826 vdd.n3186 vdd.n3185 0.0198529
R4827 vdd.n3219 vdd.n3218 0.0198529
R4828 vdd.n3240 vdd.n2218 0.0198529
R4829 vdd.n3264 vdd.n2205 0.0198529
R4830 vdd.n3386 vdd.n2130 0.0198529
R4831 vdd.n3407 vdd.n3406 0.0198529
R4832 vdd.n3412 vdd.n3411 0.0198529
R4833 vdd.n3445 vdd.n3444 0.0198529
R4834 vdd.n3466 vdd.n2084 0.0198529
R4835 vdd.n3490 vdd.n2071 0.0198529
R4836 vdd.n3612 vdd.n1996 0.0198529
R4837 vdd.n3633 vdd.n3632 0.0198529
R4838 vdd.n3638 vdd.n3637 0.0198529
R4839 vdd.n3671 vdd.n3670 0.0198529
R4840 vdd.n3692 vdd.n1950 0.0198529
R4841 vdd.n3696 vdd.n1948 0.0198529
R4842 vdd.n3743 vdd.n1926 0.0198529
R4843 vdd.n3762 vdd.n1915 0.0198529
R4844 vdd.n3781 vdd.n1904 0.0198529
R4845 vdd.n3800 vdd.n1893 0.0198529
R4846 vdd.n3819 vdd.n1878 0.0198529
R4847 vdd.n677 vdd.n676 0.018827
R4848 vdd.n1796 vdd.n1 0.0188117
R4849 vdd.n1797 vdd.n1796 0.0188117
R4850 vdd.n2780 vdd.n1871 0.0188117
R4851 vdd.n2783 vdd.n2780 0.0188117
R4852 vdd vdd.n2515 0.0187584
R4853 vdd.n705 vdd.n604 0.0185769
R4854 vdd.n709 vdd.n708 0.0185769
R4855 vdd.n740 vdd.n738 0.0185769
R4856 vdd.n764 vdd.n574 0.0185769
R4857 vdd.n787 vdd.n558 0.0185769
R4858 vdd.n791 vdd.n790 0.0185769
R4859 vdd.n829 vdd.n824 0.0185769
R4860 vdd.n852 vdd.n523 0.0185769
R4861 vdd.n877 vdd.n508 0.0185769
R4862 vdd.n899 vdd.n495 0.0185769
R4863 vdd.n911 vdd.n489 0.0185769
R4864 vdd.n926 vdd.n925 0.0185769
R4865 vdd.n956 vdd.n470 0.0185769
R4866 vdd.n960 vdd.n959 0.0185769
R4867 vdd.n991 vdd.n989 0.0185769
R4868 vdd.n1015 vdd.n440 0.0185769
R4869 vdd.n1038 vdd.n424 0.0185769
R4870 vdd.n1042 vdd.n1041 0.0185769
R4871 vdd.n1080 vdd.n1075 0.0185769
R4872 vdd.n1103 vdd.n389 0.0185769
R4873 vdd.n1128 vdd.n374 0.0185769
R4874 vdd.n1150 vdd.n361 0.0185769
R4875 vdd.n1162 vdd.n355 0.0185769
R4876 vdd.n1177 vdd.n1176 0.0185769
R4877 vdd.n1207 vdd.n336 0.0185769
R4878 vdd.n1211 vdd.n1210 0.0185769
R4879 vdd.n1242 vdd.n1240 0.0185769
R4880 vdd.n1266 vdd.n306 0.0185769
R4881 vdd.n1289 vdd.n290 0.0185769
R4882 vdd.n1293 vdd.n1292 0.0185769
R4883 vdd.n1331 vdd.n1326 0.0185769
R4884 vdd.n1354 vdd.n255 0.0185769
R4885 vdd.n1379 vdd.n240 0.0185769
R4886 vdd.n1401 vdd.n227 0.0185769
R4887 vdd.n1413 vdd.n221 0.0185769
R4888 vdd.n1428 vdd.n1427 0.0185769
R4889 vdd.n1458 vdd.n202 0.0185769
R4890 vdd.n1462 vdd.n1461 0.0185769
R4891 vdd.n1493 vdd.n1491 0.0185769
R4892 vdd.n1517 vdd.n172 0.0185769
R4893 vdd.n1540 vdd.n156 0.0185769
R4894 vdd.n1544 vdd.n1543 0.0185769
R4895 vdd.n1578 vdd.n1577 0.0185769
R4896 vdd.n1601 vdd.n1599 0.0185769
R4897 vdd.n1628 vdd.n1627 0.0185769
R4898 vdd.n1635 vdd.n1634 0.0185769
R4899 vdd.n1662 vdd.n1657 0.0185769
R4900 vdd.n1684 vdd.n71 0.0185769
R4901 vdd.n2826 vdd.n2825 0.0185769
R4902 vdd.n2847 vdd.n2845 0.0185769
R4903 vdd.n2868 vdd.n2446 0.0185769
R4904 vdd.n2890 vdd.n2432 0.0185769
R4905 vdd.n2910 vdd.n2421 0.0185769
R4906 vdd.n2929 vdd.n2399 0.0185769
R4907 vdd.n2931 vdd.n2384 0.0185769
R4908 vdd.n2963 vdd.n2962 0.0185769
R4909 vdd.n2990 vdd.n2989 0.0185769
R4910 vdd.n2997 vdd.n2996 0.0185769
R4911 vdd.n3018 vdd.n3017 0.0185769
R4912 vdd.n3042 vdd.n3041 0.0185769
R4913 vdd.n3052 vdd.n3051 0.0185769
R4914 vdd.n3073 vdd.n3071 0.0185769
R4915 vdd.n3094 vdd.n2312 0.0185769
R4916 vdd.n3116 vdd.n2298 0.0185769
R4917 vdd.n3136 vdd.n2287 0.0185769
R4918 vdd.n3155 vdd.n2265 0.0185769
R4919 vdd.n3157 vdd.n2250 0.0185769
R4920 vdd.n3189 vdd.n3188 0.0185769
R4921 vdd.n3216 vdd.n3215 0.0185769
R4922 vdd.n3223 vdd.n3222 0.0185769
R4923 vdd.n3244 vdd.n3243 0.0185769
R4924 vdd.n3268 vdd.n3267 0.0185769
R4925 vdd.n3278 vdd.n3277 0.0185769
R4926 vdd.n3299 vdd.n3297 0.0185769
R4927 vdd.n3320 vdd.n2178 0.0185769
R4928 vdd.n3342 vdd.n2164 0.0185769
R4929 vdd.n3362 vdd.n2153 0.0185769
R4930 vdd.n3381 vdd.n2131 0.0185769
R4931 vdd.n3383 vdd.n2116 0.0185769
R4932 vdd.n3415 vdd.n3414 0.0185769
R4933 vdd.n3442 vdd.n3441 0.0185769
R4934 vdd.n3449 vdd.n3448 0.0185769
R4935 vdd.n3470 vdd.n3469 0.0185769
R4936 vdd.n3494 vdd.n3493 0.0185769
R4937 vdd.n3504 vdd.n3503 0.0185769
R4938 vdd.n3525 vdd.n3523 0.0185769
R4939 vdd.n3546 vdd.n2044 0.0185769
R4940 vdd.n3568 vdd.n2030 0.0185769
R4941 vdd.n3588 vdd.n2019 0.0185769
R4942 vdd.n3607 vdd.n1997 0.0185769
R4943 vdd.n3609 vdd.n1982 0.0185769
R4944 vdd.n3641 vdd.n3640 0.0185769
R4945 vdd.n3668 vdd.n3667 0.0185769
R4946 vdd.n3675 vdd.n3674 0.0185769
R4947 vdd.n3700 vdd.n3695 0.0185769
R4948 vdd.n3716 vdd.n1936 0.0185769
R4949 vdd.n1859 vdd.n1858 0.0185349
R4950 vdd.n3824 vdd.n3823 0.0185349
R4951 vdd.n615 vdd.n614 0.0184706
R4952 vdd.n715 vdd.n714 0.0184706
R4953 vdd.n736 vdd.n735 0.0184706
R4954 vdd.n760 vdd.n575 0.0184706
R4955 vdd.n768 vdd.n767 0.0184706
R4956 vdd.n794 vdd.n793 0.0184706
R4957 vdd.n831 vdd.n535 0.0184706
R4958 vdd.n850 vdd.n524 0.0184706
R4959 vdd.n875 vdd.n509 0.0184706
R4960 vdd.n897 vdd.n496 0.0184706
R4961 vdd.n909 vdd.n490 0.0184706
R4962 vdd.n913 vdd.n488 0.0184706
R4963 vdd.n920 vdd.n919 0.0184706
R4964 vdd.n966 vdd.n965 0.0184706
R4965 vdd.n987 vdd.n986 0.0184706
R4966 vdd.n1011 vdd.n441 0.0184706
R4967 vdd.n1019 vdd.n1018 0.0184706
R4968 vdd.n1045 vdd.n1044 0.0184706
R4969 vdd.n1082 vdd.n401 0.0184706
R4970 vdd.n1101 vdd.n390 0.0184706
R4971 vdd.n1126 vdd.n375 0.0184706
R4972 vdd.n1148 vdd.n362 0.0184706
R4973 vdd.n1160 vdd.n356 0.0184706
R4974 vdd.n1164 vdd.n354 0.0184706
R4975 vdd.n1171 vdd.n1170 0.0184706
R4976 vdd.n1217 vdd.n1216 0.0184706
R4977 vdd.n1238 vdd.n1237 0.0184706
R4978 vdd.n1262 vdd.n307 0.0184706
R4979 vdd.n1270 vdd.n1269 0.0184706
R4980 vdd.n1296 vdd.n1295 0.0184706
R4981 vdd.n1333 vdd.n267 0.0184706
R4982 vdd.n1352 vdd.n256 0.0184706
R4983 vdd.n1377 vdd.n241 0.0184706
R4984 vdd.n1399 vdd.n228 0.0184706
R4985 vdd.n1411 vdd.n222 0.0184706
R4986 vdd.n1415 vdd.n220 0.0184706
R4987 vdd.n1422 vdd.n1421 0.0184706
R4988 vdd.n1468 vdd.n1467 0.0184706
R4989 vdd.n1489 vdd.n1488 0.0184706
R4990 vdd.n1513 vdd.n173 0.0184706
R4991 vdd.n1521 vdd.n1520 0.0184706
R4992 vdd.n1547 vdd.n1546 0.0184706
R4993 vdd.n1580 vdd.n134 0.0184706
R4994 vdd.n1603 vdd.n118 0.0184706
R4995 vdd.n1626 vdd.n104 0.0184706
R4996 vdd.n1637 vdd.n102 0.0184706
R4997 vdd.n1664 vdd.n85 0.0184706
R4998 vdd.n1683 vdd.n72 0.0184706
R4999 vdd.n1695 vdd.n70 0.0184706
R5000 vdd.n1718 vdd.n54 0.0184706
R5001 vdd.n1741 vdd.n40 0.0184706
R5002 vdd.n1752 vdd.n38 0.0184706
R5003 vdd.n1775 vdd.n22 0.0184706
R5004 vdd.n1862 vdd.n6 0.0184706
R5005 vdd.n2823 vdd.n2822 0.0184706
R5006 vdd.n2843 vdd.n2842 0.0184706
R5007 vdd.n2864 vdd.n2447 0.0184706
R5008 vdd.n2872 vdd.n2871 0.0184706
R5009 vdd.n2894 vdd.n2893 0.0184706
R5010 vdd.n2914 vdd.n2913 0.0184706
R5011 vdd.n2952 vdd.n2385 0.0184706
R5012 vdd.n2964 vdd.n2383 0.0184706
R5013 vdd.n2988 vdd.n2369 0.0184706
R5014 vdd.n2999 vdd.n2367 0.0184706
R5015 vdd.n3020 vdd.n2350 0.0184706
R5016 vdd.n3044 vdd.n2337 0.0184706
R5017 vdd.n3049 vdd.n3048 0.0184706
R5018 vdd.n3069 vdd.n3068 0.0184706
R5019 vdd.n3090 vdd.n2313 0.0184706
R5020 vdd.n3098 vdd.n3097 0.0184706
R5021 vdd.n3120 vdd.n3119 0.0184706
R5022 vdd.n3140 vdd.n3139 0.0184706
R5023 vdd.n3178 vdd.n2251 0.0184706
R5024 vdd.n3190 vdd.n2249 0.0184706
R5025 vdd.n3214 vdd.n2235 0.0184706
R5026 vdd.n3225 vdd.n2233 0.0184706
R5027 vdd.n3246 vdd.n2216 0.0184706
R5028 vdd.n3270 vdd.n2203 0.0184706
R5029 vdd.n3275 vdd.n3274 0.0184706
R5030 vdd.n3295 vdd.n3294 0.0184706
R5031 vdd.n3316 vdd.n2179 0.0184706
R5032 vdd.n3324 vdd.n3323 0.0184706
R5033 vdd.n3346 vdd.n3345 0.0184706
R5034 vdd.n3366 vdd.n3365 0.0184706
R5035 vdd.n3404 vdd.n2117 0.0184706
R5036 vdd.n3416 vdd.n2115 0.0184706
R5037 vdd.n3440 vdd.n2101 0.0184706
R5038 vdd.n3451 vdd.n2099 0.0184706
R5039 vdd.n3472 vdd.n2082 0.0184706
R5040 vdd.n3496 vdd.n2069 0.0184706
R5041 vdd.n3501 vdd.n3500 0.0184706
R5042 vdd.n3521 vdd.n3520 0.0184706
R5043 vdd.n3542 vdd.n2045 0.0184706
R5044 vdd.n3550 vdd.n3549 0.0184706
R5045 vdd.n3572 vdd.n3571 0.0184706
R5046 vdd.n3592 vdd.n3591 0.0184706
R5047 vdd.n3630 vdd.n1983 0.0184706
R5048 vdd.n3642 vdd.n1981 0.0184706
R5049 vdd.n3666 vdd.n1967 0.0184706
R5050 vdd.n3677 vdd.n1965 0.0184706
R5051 vdd.n3702 vdd.n1947 0.0184706
R5052 vdd.n3715 vdd.n1937 0.0184706
R5053 vdd.n3730 vdd.n1935 0.0184706
R5054 vdd.n3749 vdd.n1924 0.0184706
R5055 vdd.n3768 vdd.n1913 0.0184706
R5056 vdd.n3787 vdd.n1902 0.0184706
R5057 vdd.n3806 vdd.n1891 0.0184706
R5058 vdd.n3827 vdd.n1876 0.0184706
R5059 vdd.n616 vdd.n613 0.0179744
R5060 vdd.n707 vdd.n706 0.0179744
R5061 vdd.n737 vdd.n588 0.0179744
R5062 vdd.n739 vdd.n576 0.0179744
R5063 vdd.n766 vdd.n765 0.0179744
R5064 vdd.n792 vdd.n788 0.0179744
R5065 vdd.n823 vdd.n537 0.0179744
R5066 vdd.n828 vdd.n827 0.0179744
R5067 vdd.n854 vdd.n853 0.0179744
R5068 vdd.n879 vdd.n878 0.0179744
R5069 vdd.n901 vdd.n900 0.0179744
R5070 vdd.n927 vdd.n912 0.0179744
R5071 vdd.n922 vdd.n921 0.0179744
R5072 vdd.n958 vdd.n957 0.0179744
R5073 vdd.n988 vdd.n454 0.0179744
R5074 vdd.n990 vdd.n442 0.0179744
R5075 vdd.n1017 vdd.n1016 0.0179744
R5076 vdd.n1043 vdd.n1039 0.0179744
R5077 vdd.n1074 vdd.n403 0.0179744
R5078 vdd.n1079 vdd.n1078 0.0179744
R5079 vdd.n1105 vdd.n1104 0.0179744
R5080 vdd.n1130 vdd.n1129 0.0179744
R5081 vdd.n1152 vdd.n1151 0.0179744
R5082 vdd.n1178 vdd.n1163 0.0179744
R5083 vdd.n1173 vdd.n1172 0.0179744
R5084 vdd.n1209 vdd.n1208 0.0179744
R5085 vdd.n1239 vdd.n320 0.0179744
R5086 vdd.n1241 vdd.n308 0.0179744
R5087 vdd.n1268 vdd.n1267 0.0179744
R5088 vdd.n1294 vdd.n1290 0.0179744
R5089 vdd.n1325 vdd.n269 0.0179744
R5090 vdd.n1330 vdd.n1329 0.0179744
R5091 vdd.n1356 vdd.n1355 0.0179744
R5092 vdd.n1381 vdd.n1380 0.0179744
R5093 vdd.n1403 vdd.n1402 0.0179744
R5094 vdd.n1429 vdd.n1414 0.0179744
R5095 vdd.n1424 vdd.n1423 0.0179744
R5096 vdd.n1460 vdd.n1459 0.0179744
R5097 vdd.n1490 vdd.n186 0.0179744
R5098 vdd.n1492 vdd.n174 0.0179744
R5099 vdd.n1519 vdd.n1518 0.0179744
R5100 vdd.n1545 vdd.n1541 0.0179744
R5101 vdd.n1576 vdd.n135 0.0179744
R5102 vdd.n1598 vdd.n121 0.0179744
R5103 vdd.n1600 vdd.n105 0.0179744
R5104 vdd.n1633 vdd.n103 0.0179744
R5105 vdd.n1656 vdd.n87 0.0179744
R5106 vdd.n1661 vdd.n1660 0.0179744
R5107 vdd.n2824 vdd.n2821 0.0179744
R5108 vdd.n2844 vdd.n2458 0.0179744
R5109 vdd.n2846 vdd.n2448 0.0179744
R5110 vdd.n2870 vdd.n2869 0.0179744
R5111 vdd.n2892 vdd.n2891 0.0179744
R5112 vdd.n2912 vdd.n2911 0.0179744
R5113 vdd.n2932 vdd.n2930 0.0179744
R5114 vdd.n2957 vdd.n2956 0.0179744
R5115 vdd.n2958 vdd.n2370 0.0179744
R5116 vdd.n2995 vdd.n2368 0.0179744
R5117 vdd.n3016 vdd.n2351 0.0179744
R5118 vdd.n3040 vdd.n2338 0.0179744
R5119 vdd.n3050 vdd.n2334 0.0179744
R5120 vdd.n3070 vdd.n2324 0.0179744
R5121 vdd.n3072 vdd.n2314 0.0179744
R5122 vdd.n3096 vdd.n3095 0.0179744
R5123 vdd.n3118 vdd.n3117 0.0179744
R5124 vdd.n3138 vdd.n3137 0.0179744
R5125 vdd.n3158 vdd.n3156 0.0179744
R5126 vdd.n3183 vdd.n3182 0.0179744
R5127 vdd.n3184 vdd.n2236 0.0179744
R5128 vdd.n3221 vdd.n2234 0.0179744
R5129 vdd.n3242 vdd.n2217 0.0179744
R5130 vdd.n3266 vdd.n2204 0.0179744
R5131 vdd.n3276 vdd.n2200 0.0179744
R5132 vdd.n3296 vdd.n2190 0.0179744
R5133 vdd.n3298 vdd.n2180 0.0179744
R5134 vdd.n3322 vdd.n3321 0.0179744
R5135 vdd.n3344 vdd.n3343 0.0179744
R5136 vdd.n3364 vdd.n3363 0.0179744
R5137 vdd.n3384 vdd.n3382 0.0179744
R5138 vdd.n3409 vdd.n3408 0.0179744
R5139 vdd.n3410 vdd.n2102 0.0179744
R5140 vdd.n3447 vdd.n2100 0.0179744
R5141 vdd.n3468 vdd.n2083 0.0179744
R5142 vdd.n3492 vdd.n2070 0.0179744
R5143 vdd.n3502 vdd.n2066 0.0179744
R5144 vdd.n3522 vdd.n2056 0.0179744
R5145 vdd.n3524 vdd.n2046 0.0179744
R5146 vdd.n3548 vdd.n3547 0.0179744
R5147 vdd.n3570 vdd.n3569 0.0179744
R5148 vdd.n3590 vdd.n3589 0.0179744
R5149 vdd.n3610 vdd.n3608 0.0179744
R5150 vdd.n3635 vdd.n3634 0.0179744
R5151 vdd.n3636 vdd.n1968 0.0179744
R5152 vdd.n3673 vdd.n1966 0.0179744
R5153 vdd.n3694 vdd.n1949 0.0179744
R5154 vdd.n3699 vdd.n3698 0.0179744
R5155 vdd.n1693 vdd.n1692 0.0179074
R5156 vdd.n1716 vdd.n1714 0.0179074
R5157 vdd.n1743 vdd.n1742 0.0179074
R5158 vdd.n1750 vdd.n1749 0.0179074
R5159 vdd.n1773 vdd.n1772 0.0179074
R5160 vdd.n1860 vdd.n1857 0.0179074
R5161 vdd.n3728 vdd.n3727 0.0179074
R5162 vdd.n3747 vdd.n3746 0.0179074
R5163 vdd.n3766 vdd.n3765 0.0179074
R5164 vdd.n3785 vdd.n3784 0.0179074
R5165 vdd.n3804 vdd.n3803 0.0179074
R5166 vdd.n3825 vdd.n3822 0.0179074
R5167 vdd.n1691 vdd.n1685 0.0173272
R5168 vdd.n1713 vdd.n57 0.0173272
R5169 vdd.n1715 vdd.n41 0.0173272
R5170 vdd.n1748 vdd.n39 0.0173272
R5171 vdd.n1771 vdd.n23 0.0173272
R5172 vdd.n1856 vdd.n7 0.0173272
R5173 vdd.n3726 vdd.n3717 0.0173272
R5174 vdd.n3745 vdd.n1925 0.0173272
R5175 vdd.n3764 vdd.n1914 0.0173272
R5176 vdd.n3783 vdd.n1903 0.0173272
R5177 vdd.n3802 vdd.n1892 0.0173272
R5178 vdd.n3821 vdd.n1877 0.0173272
R5179 vdd.n660 vdd.n651 0.0172857
R5180 vdd.n2739 vdd.n2730 0.0172857
R5181 vdd vdd.n3834 0.0169115
R5182 vdd.n1858 vdd.n2 0.0168953
R5183 vdd.n1868 vdd.n2 0.0168953
R5184 vdd.n3823 vdd.n1872 0.0168953
R5185 vdd.n3833 vdd.n1872 0.0168953
R5186 vdd.n683 vdd.n682 0.0167579
R5187 vdd vdd.n1869 0.0166033
R5188 vdd.n1834 vdd.n1833 0.016125
R5189 vdd.n2776 vdd.n2760 0.016125
R5190 vdd.n2498 vdd.n2497 0.0161041
R5191 vdd.n2655 vdd.n2558 0.0159756
R5192 vdd.n2547 vdd.n2546 0.0159756
R5193 vdd.n2696 vdd.n2540 0.0159756
R5194 vdd.n2690 vdd.n2544 0.0159756
R5195 vdd.n691 vdd.n611 0.0156071
R5196 vdd.n662 vdd.n650 0.0156071
R5197 vdd.n678 vdd.n646 0.0156071
R5198 vdd.n681 vdd.n639 0.0156071
R5199 vdd.n684 vdd.n628 0.0156071
R5200 vdd.n687 vdd.n624 0.0156071
R5201 vdd.n2514 vdd.n2513 0.0156071
R5202 vdd.n2745 vdd.n2744 0.0156071
R5203 vdd.n2750 vdd.n2510 0.0156071
R5204 vdd.n2818 vdd.n2817 0.0156071
R5205 vdd.n2503 vdd.n2472 0.0156071
R5206 vdd.n2499 vdd.n2477 0.0156071
R5207 vdd.n2496 vdd.n2495 0.0156071
R5208 vdd.n2749 vdd.n2469 0.0153019
R5209 vdd.n1866 vdd.n1865 0.0152558
R5210 vdd.n3831 vdd.n3830 0.0152558
R5211 vdd.n658 vdd.n655 0.0148621
R5212 vdd.n2737 vdd.n2734 0.0148621
R5213 vdd.n680 vdd.n679 0.0148365
R5214 vdd.n2502 vdd.n2500 0.014539
R5215 vdd.n704 vdd.n602 0.0143235
R5216 vdd.n710 vdd.n589 0.0143235
R5217 vdd.n741 vdd.n587 0.0143235
R5218 vdd.n763 vdd.n573 0.0143235
R5219 vdd.n786 vdd.n556 0.0143235
R5220 vdd.n830 vdd.n536 0.0143235
R5221 vdd.n851 vdd.n522 0.0143235
R5222 vdd.n876 vdd.n507 0.0143235
R5223 vdd.n898 vdd.n494 0.0143235
R5224 vdd.n910 vdd.n487 0.0143235
R5225 vdd.n955 vdd.n468 0.0143235
R5226 vdd.n961 vdd.n455 0.0143235
R5227 vdd.n992 vdd.n453 0.0143235
R5228 vdd.n1014 vdd.n439 0.0143235
R5229 vdd.n1037 vdd.n422 0.0143235
R5230 vdd.n1081 vdd.n402 0.0143235
R5231 vdd.n1102 vdd.n388 0.0143235
R5232 vdd.n1127 vdd.n373 0.0143235
R5233 vdd.n1149 vdd.n360 0.0143235
R5234 vdd.n1161 vdd.n353 0.0143235
R5235 vdd.n1206 vdd.n334 0.0143235
R5236 vdd.n1212 vdd.n321 0.0143235
R5237 vdd.n1243 vdd.n319 0.0143235
R5238 vdd.n1265 vdd.n305 0.0143235
R5239 vdd.n1288 vdd.n288 0.0143235
R5240 vdd.n1332 vdd.n268 0.0143235
R5241 vdd.n1353 vdd.n254 0.0143235
R5242 vdd.n1378 vdd.n239 0.0143235
R5243 vdd.n1400 vdd.n226 0.0143235
R5244 vdd.n1412 vdd.n219 0.0143235
R5245 vdd.n1457 vdd.n200 0.0143235
R5246 vdd.n1463 vdd.n187 0.0143235
R5247 vdd.n1494 vdd.n185 0.0143235
R5248 vdd.n1516 vdd.n171 0.0143235
R5249 vdd.n1539 vdd.n154 0.0143235
R5250 vdd.n1579 vdd.n122 0.0143235
R5251 vdd.n1602 vdd.n120 0.0143235
R5252 vdd.n1630 vdd.n1629 0.0143235
R5253 vdd.n1636 vdd.n88 0.0143235
R5254 vdd.n1663 vdd.n86 0.0143235
R5255 vdd.n1694 vdd.n58 0.0143235
R5256 vdd.n1717 vdd.n56 0.0143235
R5257 vdd.n1745 vdd.n1744 0.0143235
R5258 vdd.n1751 vdd.n24 0.0143235
R5259 vdd.n1774 vdd.n8 0.0143235
R5260 vdd.n2827 vdd.n2459 0.0143235
R5261 vdd.n2848 vdd.n2457 0.0143235
R5262 vdd.n2867 vdd.n2445 0.0143235
R5263 vdd.n2889 vdd.n2431 0.0143235
R5264 vdd.n2909 vdd.n2420 0.0143235
R5265 vdd.n2955 vdd.n2953 0.0143235
R5266 vdd.n2961 vdd.n2960 0.0143235
R5267 vdd.n2992 vdd.n2991 0.0143235
R5268 vdd.n2998 vdd.n2352 0.0143235
R5269 vdd.n3019 vdd.n2339 0.0143235
R5270 vdd.n3053 vdd.n2325 0.0143235
R5271 vdd.n3074 vdd.n2323 0.0143235
R5272 vdd.n3093 vdd.n2311 0.0143235
R5273 vdd.n3115 vdd.n2297 0.0143235
R5274 vdd.n3135 vdd.n2286 0.0143235
R5275 vdd.n3181 vdd.n3179 0.0143235
R5276 vdd.n3187 vdd.n3186 0.0143235
R5277 vdd.n3218 vdd.n3217 0.0143235
R5278 vdd.n3224 vdd.n2218 0.0143235
R5279 vdd.n3245 vdd.n2205 0.0143235
R5280 vdd.n3279 vdd.n2191 0.0143235
R5281 vdd.n3300 vdd.n2189 0.0143235
R5282 vdd.n3319 vdd.n2177 0.0143235
R5283 vdd.n3341 vdd.n2163 0.0143235
R5284 vdd.n3361 vdd.n2152 0.0143235
R5285 vdd.n3407 vdd.n3405 0.0143235
R5286 vdd.n3413 vdd.n3412 0.0143235
R5287 vdd.n3444 vdd.n3443 0.0143235
R5288 vdd.n3450 vdd.n2084 0.0143235
R5289 vdd.n3471 vdd.n2071 0.0143235
R5290 vdd.n3505 vdd.n2057 0.0143235
R5291 vdd.n3526 vdd.n2055 0.0143235
R5292 vdd.n3545 vdd.n2043 0.0143235
R5293 vdd.n3567 vdd.n2029 0.0143235
R5294 vdd.n3587 vdd.n2018 0.0143235
R5295 vdd.n3633 vdd.n3631 0.0143235
R5296 vdd.n3639 vdd.n3638 0.0143235
R5297 vdd.n3670 vdd.n3669 0.0143235
R5298 vdd.n3676 vdd.n1950 0.0143235
R5299 vdd.n3701 vdd.n1948 0.0143235
R5300 vdd.n3729 vdd.n1926 0.0143235
R5301 vdd.n3748 vdd.n1915 0.0143235
R5302 vdd.n3767 vdd.n1904 0.0143235
R5303 vdd.n3786 vdd.n1893 0.0143235
R5304 vdd.n3805 vdd.n1878 0.0143235
R5305 vdd.n686 vdd.n685 0.0140975
R5306 vdd.n1819 vdd.n1808 0.0140135
R5307 vdd.n2803 vdd.n2762 0.0140135
R5308 vdd.n716 vdd.n601 0.0137576
R5309 vdd.n734 vdd.n733 0.0137576
R5310 vdd.n758 vdd.n757 0.0137576
R5311 vdd.n769 vdd.n572 0.0137576
R5312 vdd.n795 vdd.n555 0.0137576
R5313 vdd.n832 vdd.n534 0.0137576
R5314 vdd.n849 vdd.n848 0.0137576
R5315 vdd.n874 vdd.n510 0.0137576
R5316 vdd.n896 vdd.n497 0.0137576
R5317 vdd.n908 vdd.n907 0.0137576
R5318 vdd.n916 vdd.n915 0.0137576
R5319 vdd.n918 vdd.n917 0.0137576
R5320 vdd.n967 vdd.n467 0.0137576
R5321 vdd.n985 vdd.n984 0.0137576
R5322 vdd.n1009 vdd.n1008 0.0137576
R5323 vdd.n1020 vdd.n438 0.0137576
R5324 vdd.n1046 vdd.n421 0.0137576
R5325 vdd.n1083 vdd.n400 0.0137576
R5326 vdd.n1100 vdd.n1099 0.0137576
R5327 vdd.n1125 vdd.n376 0.0137576
R5328 vdd.n1147 vdd.n363 0.0137576
R5329 vdd.n1159 vdd.n1158 0.0137576
R5330 vdd.n1167 vdd.n1166 0.0137576
R5331 vdd.n1169 vdd.n1168 0.0137576
R5332 vdd.n1218 vdd.n333 0.0137576
R5333 vdd.n1236 vdd.n1235 0.0137576
R5334 vdd.n1260 vdd.n1259 0.0137576
R5335 vdd.n1271 vdd.n304 0.0137576
R5336 vdd.n1297 vdd.n287 0.0137576
R5337 vdd.n1334 vdd.n266 0.0137576
R5338 vdd.n1351 vdd.n1350 0.0137576
R5339 vdd.n1376 vdd.n242 0.0137576
R5340 vdd.n1398 vdd.n229 0.0137576
R5341 vdd.n1410 vdd.n1409 0.0137576
R5342 vdd.n1418 vdd.n1417 0.0137576
R5343 vdd.n1420 vdd.n1419 0.0137576
R5344 vdd.n1469 vdd.n199 0.0137576
R5345 vdd.n1487 vdd.n1486 0.0137576
R5346 vdd.n1511 vdd.n1510 0.0137576
R5347 vdd.n1522 vdd.n170 0.0137576
R5348 vdd.n1548 vdd.n153 0.0137576
R5349 vdd.n1581 vdd.n133 0.0137576
R5350 vdd.n1604 vdd.n117 0.0137576
R5351 vdd.n1624 vdd.n108 0.0137576
R5352 vdd.n1639 vdd.n1638 0.0137576
R5353 vdd.n1665 vdd.n84 0.0137576
R5354 vdd.n1696 vdd.n69 0.0137576
R5355 vdd.n1719 vdd.n53 0.0137576
R5356 vdd.n1739 vdd.n44 0.0137576
R5357 vdd.n1754 vdd.n1753 0.0137576
R5358 vdd.n1776 vdd.n21 0.0137576
R5359 vdd.n1863 vdd.n5 0.0137576
R5360 vdd.n2841 vdd.n2840 0.0137576
R5361 vdd.n2862 vdd.n2861 0.0137576
R5362 vdd.n2873 vdd.n2444 0.0137576
R5363 vdd.n2895 vdd.n2430 0.0137576
R5364 vdd.n2915 vdd.n2419 0.0137576
R5365 vdd.n2951 vdd.n2386 0.0137576
R5366 vdd.n2966 vdd.n2379 0.0137576
R5367 vdd.n2986 vdd.n2373 0.0137576
R5368 vdd.n3001 vdd.n3000 0.0137576
R5369 vdd.n3021 vdd.n2349 0.0137576
R5370 vdd.n3045 vdd.n2336 0.0137576
R5371 vdd.n3047 vdd.n3046 0.0137576
R5372 vdd.n3067 vdd.n3066 0.0137576
R5373 vdd.n3088 vdd.n3087 0.0137576
R5374 vdd.n3099 vdd.n2310 0.0137576
R5375 vdd.n3121 vdd.n2296 0.0137576
R5376 vdd.n3141 vdd.n2285 0.0137576
R5377 vdd.n3177 vdd.n2252 0.0137576
R5378 vdd.n3192 vdd.n2245 0.0137576
R5379 vdd.n3212 vdd.n2239 0.0137576
R5380 vdd.n3227 vdd.n3226 0.0137576
R5381 vdd.n3247 vdd.n2215 0.0137576
R5382 vdd.n3271 vdd.n2202 0.0137576
R5383 vdd.n3273 vdd.n3272 0.0137576
R5384 vdd.n3293 vdd.n3292 0.0137576
R5385 vdd.n3314 vdd.n3313 0.0137576
R5386 vdd.n3325 vdd.n2176 0.0137576
R5387 vdd.n3347 vdd.n2162 0.0137576
R5388 vdd.n3367 vdd.n2151 0.0137576
R5389 vdd.n3403 vdd.n2118 0.0137576
R5390 vdd.n3418 vdd.n2111 0.0137576
R5391 vdd.n3438 vdd.n2105 0.0137576
R5392 vdd.n3453 vdd.n3452 0.0137576
R5393 vdd.n3473 vdd.n2081 0.0137576
R5394 vdd.n3497 vdd.n2068 0.0137576
R5395 vdd.n3499 vdd.n3498 0.0137576
R5396 vdd.n3519 vdd.n3518 0.0137576
R5397 vdd.n3540 vdd.n3539 0.0137576
R5398 vdd.n3551 vdd.n2042 0.0137576
R5399 vdd.n3573 vdd.n2028 0.0137576
R5400 vdd.n3593 vdd.n2017 0.0137576
R5401 vdd.n3629 vdd.n1984 0.0137576
R5402 vdd.n3644 vdd.n1977 0.0137576
R5403 vdd.n3664 vdd.n1971 0.0137576
R5404 vdd.n3679 vdd.n3678 0.0137576
R5405 vdd.n3703 vdd.n1946 0.0137576
R5406 vdd.n3731 vdd.n1934 0.0137576
R5407 vdd.n3750 vdd.n1923 0.0137576
R5408 vdd.n3769 vdd.n1912 0.0137576
R5409 vdd.n3788 vdd.n1901 0.0137576
R5410 vdd.n3807 vdd.n1890 0.0137576
R5411 vdd.n3828 vdd.n1875 0.0137576
R5412 vdd.n657 vdd.n653 0.0137243
R5413 vdd.n2736 vdd.n2732 0.0137243
R5414 vdd.n1817 vdd.n1816 0.0137188
R5415 vdd.n2802 vdd.n2779 0.0137188
R5416 vdd.n2802 vdd.n2781 0.0137188
R5417 vdd.n2617 vdd.n2616 0.0134151
R5418 vdd.n1801 vdd.n1795 0.0130393
R5419 vdd.n1814 vdd.n1813 0.0130393
R5420 vdd.n2769 vdd.n2768 0.0130393
R5421 vdd.n2785 vdd.n2782 0.0130393
R5422 vdd.n690 vdd.n688 0.0129151
R5423 vdd.n2820 vdd.n2466 0.0125552
R5424 vdd.n706 vdd.n705 0.0125513
R5425 vdd.n709 vdd.n588 0.0125513
R5426 vdd.n740 vdd.n739 0.0125513
R5427 vdd.n765 vdd.n764 0.0125513
R5428 vdd.n788 vdd.n787 0.0125513
R5429 vdd.n829 vdd.n828 0.0125513
R5430 vdd.n853 vdd.n852 0.0125513
R5431 vdd.n878 vdd.n877 0.0125513
R5432 vdd.n900 vdd.n899 0.0125513
R5433 vdd.n912 vdd.n911 0.0125513
R5434 vdd.n957 vdd.n956 0.0125513
R5435 vdd.n960 vdd.n454 0.0125513
R5436 vdd.n991 vdd.n990 0.0125513
R5437 vdd.n1016 vdd.n1015 0.0125513
R5438 vdd.n1039 vdd.n1038 0.0125513
R5439 vdd.n1080 vdd.n1079 0.0125513
R5440 vdd.n1104 vdd.n1103 0.0125513
R5441 vdd.n1129 vdd.n1128 0.0125513
R5442 vdd.n1151 vdd.n1150 0.0125513
R5443 vdd.n1163 vdd.n1162 0.0125513
R5444 vdd.n1208 vdd.n1207 0.0125513
R5445 vdd.n1211 vdd.n320 0.0125513
R5446 vdd.n1242 vdd.n1241 0.0125513
R5447 vdd.n1267 vdd.n1266 0.0125513
R5448 vdd.n1290 vdd.n1289 0.0125513
R5449 vdd.n1331 vdd.n1330 0.0125513
R5450 vdd.n1355 vdd.n1354 0.0125513
R5451 vdd.n1380 vdd.n1379 0.0125513
R5452 vdd.n1402 vdd.n1401 0.0125513
R5453 vdd.n1414 vdd.n1413 0.0125513
R5454 vdd.n1459 vdd.n1458 0.0125513
R5455 vdd.n1462 vdd.n186 0.0125513
R5456 vdd.n1493 vdd.n1492 0.0125513
R5457 vdd.n1518 vdd.n1517 0.0125513
R5458 vdd.n1541 vdd.n1540 0.0125513
R5459 vdd.n1578 vdd.n121 0.0125513
R5460 vdd.n1601 vdd.n1600 0.0125513
R5461 vdd.n1628 vdd.n103 0.0125513
R5462 vdd.n1635 vdd.n87 0.0125513
R5463 vdd.n1662 vdd.n1661 0.0125513
R5464 vdd.n2826 vdd.n2458 0.0125513
R5465 vdd.n2847 vdd.n2846 0.0125513
R5466 vdd.n2869 vdd.n2868 0.0125513
R5467 vdd.n2891 vdd.n2890 0.0125513
R5468 vdd.n2911 vdd.n2910 0.0125513
R5469 vdd.n2956 vdd.n2384 0.0125513
R5470 vdd.n2962 vdd.n2958 0.0125513
R5471 vdd.n2990 vdd.n2368 0.0125513
R5472 vdd.n2997 vdd.n2351 0.0125513
R5473 vdd.n3018 vdd.n2338 0.0125513
R5474 vdd.n3052 vdd.n2324 0.0125513
R5475 vdd.n3073 vdd.n3072 0.0125513
R5476 vdd.n3095 vdd.n3094 0.0125513
R5477 vdd.n3117 vdd.n3116 0.0125513
R5478 vdd.n3137 vdd.n3136 0.0125513
R5479 vdd.n3182 vdd.n2250 0.0125513
R5480 vdd.n3188 vdd.n3184 0.0125513
R5481 vdd.n3216 vdd.n2234 0.0125513
R5482 vdd.n3223 vdd.n2217 0.0125513
R5483 vdd.n3244 vdd.n2204 0.0125513
R5484 vdd.n3278 vdd.n2190 0.0125513
R5485 vdd.n3299 vdd.n3298 0.0125513
R5486 vdd.n3321 vdd.n3320 0.0125513
R5487 vdd.n3343 vdd.n3342 0.0125513
R5488 vdd.n3363 vdd.n3362 0.0125513
R5489 vdd.n3408 vdd.n2116 0.0125513
R5490 vdd.n3414 vdd.n3410 0.0125513
R5491 vdd.n3442 vdd.n2100 0.0125513
R5492 vdd.n3449 vdd.n2083 0.0125513
R5493 vdd.n3470 vdd.n2070 0.0125513
R5494 vdd.n3504 vdd.n2056 0.0125513
R5495 vdd.n3525 vdd.n3524 0.0125513
R5496 vdd.n3547 vdd.n3546 0.0125513
R5497 vdd.n3569 vdd.n3568 0.0125513
R5498 vdd.n3589 vdd.n3588 0.0125513
R5499 vdd.n3634 vdd.n1982 0.0125513
R5500 vdd.n3640 vdd.n3636 0.0125513
R5501 vdd.n3668 vdd.n1966 0.0125513
R5502 vdd.n3675 vdd.n1949 0.0125513
R5503 vdd.n3700 vdd.n3699 0.0125513
R5504 vdd.n2652 vdd 0.0124926
R5505 vdd.n2516 vdd 0.0124382
R5506 vdd.n3834 vdd 0.0122885
R5507 vdd.n1693 vdd.n57 0.0121049
R5508 vdd.n1716 vdd.n1715 0.0121049
R5509 vdd.n1743 vdd.n39 0.0121049
R5510 vdd.n1750 vdd.n23 0.0121049
R5511 vdd.n1773 vdd.n7 0.0121049
R5512 vdd.n3728 vdd.n1925 0.0121049
R5513 vdd.n3747 vdd.n1914 0.0121049
R5514 vdd.n3766 vdd.n1903 0.0121049
R5515 vdd.n3785 vdd.n1892 0.0121049
R5516 vdd.n3804 vdd.n1877 0.0121049
R5517 vdd.n665 vdd 0.0108155
R5518 vdd.n659 vdd.n654 0.0105714
R5519 vdd.n2738 vdd.n2733 0.0105714
R5520 vdd.n693 vdd.n692 0.0103794
R5521 vdd.n645 vdd.n642 0.0103794
R5522 vdd.n638 vdd.n631 0.0103794
R5523 vdd.n633 vdd.n627 0.0103794
R5524 vdd.n623 vdd.n620 0.0103794
R5525 vdd.n2752 vdd.n2751 0.0103794
R5526 vdd.n2816 vdd.n2470 0.0103794
R5527 vdd.n2505 vdd.n2504 0.0103794
R5528 vdd.n2487 vdd.n2476 0.0103794
R5529 vdd.n2494 vdd.n2480 0.0103794
R5530 vdd.n719 vdd.n718 0.0099697
R5531 vdd.n731 vdd.n730 0.0099697
R5532 vdd.n755 vdd.n754 0.0099697
R5533 vdd.n770 vdd.n571 0.0099697
R5534 vdd.n798 vdd.n797 0.0099697
R5535 vdd.n814 vdd.n813 0.0099697
R5536 vdd.n544 vdd.n541 0.0099697
R5537 vdd.n836 vdd.n835 0.0099697
R5538 vdd.n860 vdd.n518 0.0099697
R5539 vdd.n872 vdd.n871 0.0099697
R5540 vdd.n894 vdd.n893 0.0099697
R5541 vdd.n933 vdd.n484 0.0099697
R5542 vdd.n970 vdd.n969 0.0099697
R5543 vdd.n982 vdd.n981 0.0099697
R5544 vdd.n1006 vdd.n1005 0.0099697
R5545 vdd.n1021 vdd.n437 0.0099697
R5546 vdd.n1049 vdd.n1048 0.0099697
R5547 vdd.n1065 vdd.n1064 0.0099697
R5548 vdd.n410 vdd.n407 0.0099697
R5549 vdd.n1087 vdd.n1086 0.0099697
R5550 vdd.n1111 vdd.n384 0.0099697
R5551 vdd.n1123 vdd.n1122 0.0099697
R5552 vdd.n1145 vdd.n1144 0.0099697
R5553 vdd.n1184 vdd.n350 0.0099697
R5554 vdd.n1221 vdd.n1220 0.0099697
R5555 vdd.n1233 vdd.n1232 0.0099697
R5556 vdd.n1257 vdd.n1256 0.0099697
R5557 vdd.n1272 vdd.n303 0.0099697
R5558 vdd.n1300 vdd.n1299 0.0099697
R5559 vdd.n1316 vdd.n1315 0.0099697
R5560 vdd.n276 vdd.n273 0.0099697
R5561 vdd.n1338 vdd.n1337 0.0099697
R5562 vdd.n1362 vdd.n250 0.0099697
R5563 vdd.n1374 vdd.n1373 0.0099697
R5564 vdd.n1396 vdd.n1395 0.0099697
R5565 vdd.n1435 vdd.n216 0.0099697
R5566 vdd.n1472 vdd.n1471 0.0099697
R5567 vdd.n1484 vdd.n1483 0.0099697
R5568 vdd.n1508 vdd.n1507 0.0099697
R5569 vdd.n1523 vdd.n169 0.0099697
R5570 vdd.n1551 vdd.n1550 0.0099697
R5571 vdd.n1567 vdd.n1566 0.0099697
R5572 vdd.n142 vdd.n139 0.0099697
R5573 vdd.n1584 vdd.n1583 0.0099697
R5574 vdd.n1608 vdd.n116 0.0099697
R5575 vdd.n1622 vdd.n1619 0.0099697
R5576 vdd.n99 vdd.n91 0.0099697
R5577 vdd.n1669 vdd.n1668 0.0099697
R5578 vdd.n1699 vdd.n1698 0.0099697
R5579 vdd.n1723 vdd.n52 0.0099697
R5580 vdd.n1737 vdd.n1734 0.0099697
R5581 vdd.n35 vdd.n27 0.0099697
R5582 vdd.n1779 vdd.n1778 0.0099697
R5583 vdd.n2838 vdd.n2837 0.0099697
R5584 vdd.n2859 vdd.n2858 0.0099697
R5585 vdd.n2874 vdd.n2443 0.0099697
R5586 vdd.n2898 vdd.n2897 0.0099697
R5587 vdd.n2918 vdd.n2917 0.0099697
R5588 vdd.n2412 vdd.n2411 0.0099697
R5589 vdd.n2408 vdd.n2407 0.0099697
R5590 vdd.n2949 vdd.n2948 0.0099697
R5591 vdd.n2968 vdd.n2378 0.0099697
R5592 vdd.n2984 vdd.n2981 0.0099697
R5593 vdd.n2364 vdd.n2363 0.0099697
R5594 vdd.n3024 vdd.n3023 0.0099697
R5595 vdd.n3064 vdd.n3063 0.0099697
R5596 vdd.n3085 vdd.n3084 0.0099697
R5597 vdd.n3100 vdd.n2309 0.0099697
R5598 vdd.n3124 vdd.n3123 0.0099697
R5599 vdd.n3144 vdd.n3143 0.0099697
R5600 vdd.n2278 vdd.n2277 0.0099697
R5601 vdd.n2274 vdd.n2273 0.0099697
R5602 vdd.n3175 vdd.n3174 0.0099697
R5603 vdd.n3194 vdd.n2244 0.0099697
R5604 vdd.n3210 vdd.n3207 0.0099697
R5605 vdd.n2230 vdd.n2229 0.0099697
R5606 vdd.n3250 vdd.n3249 0.0099697
R5607 vdd.n3290 vdd.n3289 0.0099697
R5608 vdd.n3311 vdd.n3310 0.0099697
R5609 vdd.n3326 vdd.n2175 0.0099697
R5610 vdd.n3350 vdd.n3349 0.0099697
R5611 vdd.n3370 vdd.n3369 0.0099697
R5612 vdd.n2144 vdd.n2143 0.0099697
R5613 vdd.n2140 vdd.n2139 0.0099697
R5614 vdd.n3401 vdd.n3400 0.0099697
R5615 vdd.n3420 vdd.n2110 0.0099697
R5616 vdd.n3436 vdd.n3433 0.0099697
R5617 vdd.n2096 vdd.n2095 0.0099697
R5618 vdd.n3476 vdd.n3475 0.0099697
R5619 vdd.n3516 vdd.n3515 0.0099697
R5620 vdd.n3537 vdd.n3536 0.0099697
R5621 vdd.n3552 vdd.n2041 0.0099697
R5622 vdd.n3576 vdd.n3575 0.0099697
R5623 vdd.n3596 vdd.n3595 0.0099697
R5624 vdd.n2010 vdd.n2009 0.0099697
R5625 vdd.n2006 vdd.n2005 0.0099697
R5626 vdd.n3627 vdd.n3626 0.0099697
R5627 vdd.n3646 vdd.n1976 0.0099697
R5628 vdd.n3662 vdd.n3659 0.0099697
R5629 vdd.n1962 vdd.n1961 0.0099697
R5630 vdd.n3707 vdd.n3706 0.0099697
R5631 vdd.n3734 vdd.n3733 0.0099697
R5632 vdd.n3753 vdd.n3752 0.0099697
R5633 vdd.n3772 vdd.n3771 0.0099697
R5634 vdd.n3791 vdd.n3790 0.0099697
R5635 vdd.n3810 vdd.n3809 0.0099697
R5636 vdd.n2652 vdd.n2651 0.00926384
R5637 vdd.n676 vdd.n663 0.00907233
R5638 vdd.n1869 vdd.n1 0.00833333
R5639 vdd vdd.n1871 0.00833333
R5640 vdd.n2617 vdd 0.00788007
R5641 vdd.n1835 vdd.n1834 0.00701042
R5642 vdd.n1833 vdd.n1821 0.00701042
R5643 vdd.n2777 vdd.n2776 0.00701042
R5644 vdd.n2805 vdd.n2760 0.00701042
R5645 vdd.n2685 vdd 0.00649631
R5646 vdd.n691 vdd.n612 0.00635126
R5647 vdd.n678 vdd.n641 0.00635126
R5648 vdd.n681 vdd.n630 0.00635126
R5649 vdd.n684 vdd.n626 0.00635126
R5650 vdd.n687 vdd.n619 0.00635126
R5651 vdd.n2750 vdd.n2511 0.00635126
R5652 vdd.n2818 vdd.n2468 0.00635126
R5653 vdd.n2503 vdd.n2473 0.00635126
R5654 vdd.n2499 vdd.n2475 0.00635126
R5655 vdd.n2496 vdd.n2479 0.00635126
R5656 vdd.n2654 vdd.n2653 0.00543007
R5657 vdd.n2654 vdd.n2560 0.00543007
R5658 vdd.n2559 vdd.n2545 0.00543007
R5659 vdd.n2688 vdd.n2545 0.00543007
R5660 vdd.n2689 vdd.n2543 0.00543007
R5661 vdd.n2693 vdd.n2543 0.00543007
R5662 vdd.n2695 vdd.n2694 0.00543007
R5663 vdd.n2695 vdd.n2542 0.00543007
R5664 vdd.n2541 vdd.n2512 0.00543007
R5665 vdd.n2728 vdd.n2512 0.00543007
R5666 vdd.n2820 vdd.n2819 0.00523052
R5667 vdd.n2659 vdd.n2658 0.00511255
R5668 vdd.n2498 vdd.n2474 0.00507792
R5669 vdd.n2500 vdd.n2474 0.00507792
R5670 vdd.n2502 vdd.n2501 0.00507792
R5671 vdd.n2501 vdd.n2466 0.00507792
R5672 vdd.n2819 vdd.n2467 0.00507792
R5673 vdd.n2469 vdd.n2467 0.00507792
R5674 vdd.n2749 vdd.n2748 0.00507792
R5675 vdd.n2748 vdd.n2747 0.00507792
R5676 vdd.n2742 vdd.n2740 0.00507792
R5677 vdd.n661 vdd.n647 0.00493396
R5678 vdd.n663 vdd.n647 0.00493396
R5679 vdd.n677 vdd.n640 0.00493396
R5680 vdd.n679 vdd.n640 0.00493396
R5681 vdd.n680 vdd.n629 0.00493396
R5682 vdd.n682 vdd.n629 0.00493396
R5683 vdd.n683 vdd.n625 0.00493396
R5684 vdd.n685 vdd.n625 0.00493396
R5685 vdd.n686 vdd.n618 0.00493396
R5686 vdd.n688 vdd.n618 0.00493396
R5687 vdd.n690 vdd.n689 0.00493396
R5688 vdd.n689 vdd.n617 0.00493396
R5689 vdd.n2766 vdd.n1870 0.00490305
R5690 vdd.n2742 vdd.n2729 0.00462013
R5691 vdd.n1821 vdd.n1820 0.00440625
R5692 vdd.n2805 vdd.n2804 0.00440625
R5693 vdd.n702 vdd.n606 0.00428788
R5694 vdd.n713 vdd.n712 0.00428788
R5695 vdd.n743 vdd.n585 0.00428788
R5696 vdd.n759 vdd.n569 0.00428788
R5697 vdd.n784 vdd.n560 0.00428788
R5698 vdd.n809 vdd.n545 0.00428788
R5699 vdd.n820 vdd.n540 0.00428788
R5700 vdd.n527 vdd.n525 0.00428788
R5701 vdd.n857 vdd.n521 0.00428788
R5702 vdd.n882 vdd.n506 0.00428788
R5703 vdd.n904 vdd.n491 0.00428788
R5704 vdd.n930 vdd.n486 0.00428788
R5705 vdd.n953 vdd.n472 0.00428788
R5706 vdd.n964 vdd.n963 0.00428788
R5707 vdd.n994 vdd.n451 0.00428788
R5708 vdd.n1010 vdd.n435 0.00428788
R5709 vdd.n1035 vdd.n426 0.00428788
R5710 vdd.n1060 vdd.n411 0.00428788
R5711 vdd.n1071 vdd.n406 0.00428788
R5712 vdd.n393 vdd.n391 0.00428788
R5713 vdd.n1108 vdd.n387 0.00428788
R5714 vdd.n1133 vdd.n372 0.00428788
R5715 vdd.n1155 vdd.n357 0.00428788
R5716 vdd.n1181 vdd.n352 0.00428788
R5717 vdd.n1204 vdd.n338 0.00428788
R5718 vdd.n1215 vdd.n1214 0.00428788
R5719 vdd.n1245 vdd.n317 0.00428788
R5720 vdd.n1261 vdd.n301 0.00428788
R5721 vdd.n1286 vdd.n292 0.00428788
R5722 vdd.n1311 vdd.n277 0.00428788
R5723 vdd.n1322 vdd.n272 0.00428788
R5724 vdd.n259 vdd.n257 0.00428788
R5725 vdd.n1359 vdd.n253 0.00428788
R5726 vdd.n1384 vdd.n238 0.00428788
R5727 vdd.n1406 vdd.n223 0.00428788
R5728 vdd.n1432 vdd.n218 0.00428788
R5729 vdd.n1455 vdd.n204 0.00428788
R5730 vdd.n1466 vdd.n1465 0.00428788
R5731 vdd.n1496 vdd.n183 0.00428788
R5732 vdd.n1512 vdd.n167 0.00428788
R5733 vdd.n1537 vdd.n158 0.00428788
R5734 vdd.n1562 vdd.n143 0.00428788
R5735 vdd.n1573 vdd.n138 0.00428788
R5736 vdd.n1595 vdd.n124 0.00428788
R5737 vdd.n1625 vdd.n107 0.00428788
R5738 vdd.n100 vdd.n98 0.00428788
R5739 vdd.n1653 vdd.n90 0.00428788
R5740 vdd.n75 vdd.n73 0.00428788
R5741 vdd.n1688 vdd.n1687 0.00428788
R5742 vdd.n1710 vdd.n60 0.00428788
R5743 vdd.n1740 vdd.n43 0.00428788
R5744 vdd.n36 vdd.n34 0.00428788
R5745 vdd.n1768 vdd.n26 0.00428788
R5746 vdd.n1853 vdd.n10 0.00428788
R5747 vdd.n2829 vdd.n2464 0.00428788
R5748 vdd.n2850 vdd.n2455 0.00428788
R5749 vdd.n2863 vdd.n2441 0.00428788
R5750 vdd.n2887 vdd.n2434 0.00428788
R5751 vdd.n2907 vdd.n2423 0.00428788
R5752 vdd.n2926 vdd.n2401 0.00428788
R5753 vdd.n2935 vdd.n2397 0.00428788
R5754 vdd.n2965 vdd.n2381 0.00428788
R5755 vdd.n2987 vdd.n2372 0.00428788
R5756 vdd.n2365 vdd.n2361 0.00428788
R5757 vdd.n3013 vdd.n2354 0.00428788
R5758 vdd.n3037 vdd.n2341 0.00428788
R5759 vdd.n3055 vdd.n2332 0.00428788
R5760 vdd.n3076 vdd.n2321 0.00428788
R5761 vdd.n3089 vdd.n2307 0.00428788
R5762 vdd.n3113 vdd.n2300 0.00428788
R5763 vdd.n3133 vdd.n2289 0.00428788
R5764 vdd.n3152 vdd.n2267 0.00428788
R5765 vdd.n3161 vdd.n2263 0.00428788
R5766 vdd.n3191 vdd.n2247 0.00428788
R5767 vdd.n3213 vdd.n2238 0.00428788
R5768 vdd.n2231 vdd.n2227 0.00428788
R5769 vdd.n3239 vdd.n2220 0.00428788
R5770 vdd.n3263 vdd.n2207 0.00428788
R5771 vdd.n3281 vdd.n2198 0.00428788
R5772 vdd.n3302 vdd.n2187 0.00428788
R5773 vdd.n3315 vdd.n2173 0.00428788
R5774 vdd.n3339 vdd.n2166 0.00428788
R5775 vdd.n3359 vdd.n2155 0.00428788
R5776 vdd.n3378 vdd.n2133 0.00428788
R5777 vdd.n3387 vdd.n2129 0.00428788
R5778 vdd.n3417 vdd.n2113 0.00428788
R5779 vdd.n3439 vdd.n2104 0.00428788
R5780 vdd.n2097 vdd.n2093 0.00428788
R5781 vdd.n3465 vdd.n2086 0.00428788
R5782 vdd.n3489 vdd.n2073 0.00428788
R5783 vdd.n3507 vdd.n2064 0.00428788
R5784 vdd.n3528 vdd.n2053 0.00428788
R5785 vdd.n3541 vdd.n2039 0.00428788
R5786 vdd.n3565 vdd.n2032 0.00428788
R5787 vdd.n3585 vdd.n2021 0.00428788
R5788 vdd.n3604 vdd.n1999 0.00428788
R5789 vdd.n3613 vdd.n1995 0.00428788
R5790 vdd.n3643 vdd.n1979 0.00428788
R5791 vdd.n3665 vdd.n1970 0.00428788
R5792 vdd.n1963 vdd.n1959 0.00428788
R5793 vdd.n3691 vdd.n1952 0.00428788
R5794 vdd.n1940 vdd.n1938 0.00428788
R5795 vdd.n3723 vdd.n3718 0.00428788
R5796 vdd.n3742 vdd.n1928 0.00428788
R5797 vdd.n3761 vdd.n1917 0.00428788
R5798 vdd.n3780 vdd.n1906 0.00428788
R5799 vdd.n3799 vdd.n1895 0.00428788
R5800 vdd.n3818 vdd.n1880 0.00428788
R5801 vdd.n1811 vdd.n1810 0.00428087
R5802 vdd.n1800 vdd.n1799 0.00428087
R5803 vdd.n2800 vdd.n2799 0.00428087
R5804 vdd.n2656 vdd.n2655 0.00404637
R5805 vdd.n2687 vdd.n2546 0.00404637
R5806 vdd.n2697 vdd.n2696 0.00404637
R5807 vdd.n2692 vdd.n2544 0.00404637
R5808 vdd.n2727 vdd.n2513 0.00397409
R5809 vdd.n1867 vdd.n1866 0.00391036
R5810 vdd.n3832 vdd.n3831 0.00391036
R5811 vdd vdd.n1868 0.00377907
R5812 vdd vdd.n3833 0.00377907
R5813 vdd.n1813 vdd.n1811 0.00360776
R5814 vdd.n1801 vdd.n1800 0.00360776
R5815 vdd.n2769 vdd.n1870 0.00360776
R5816 vdd.n2800 vdd.n2782 0.00360776
R5817 vdd.n659 vdd.n652 0.00351641
R5818 vdd.n2738 vdd.n2731 0.00351641
R5819 vdd.n2497 vdd.n2478 0.00328896
R5820 vdd.n831 vdd.n830 0.00326471
R5821 vdd.n851 vdd.n850 0.00326471
R5822 vdd.n876 vdd.n875 0.00326471
R5823 vdd.n898 vdd.n897 0.00326471
R5824 vdd.n910 vdd.n909 0.00326471
R5825 vdd.n924 vdd.n913 0.00326471
R5826 vdd.n1082 vdd.n1081 0.00326471
R5827 vdd.n1102 vdd.n1101 0.00326471
R5828 vdd.n1127 vdd.n1126 0.00326471
R5829 vdd.n1149 vdd.n1148 0.00326471
R5830 vdd.n1161 vdd.n1160 0.00326471
R5831 vdd.n1175 vdd.n1164 0.00326471
R5832 vdd.n1333 vdd.n1332 0.00326471
R5833 vdd.n1353 vdd.n1352 0.00326471
R5834 vdd.n1378 vdd.n1377 0.00326471
R5835 vdd.n1400 vdd.n1399 0.00326471
R5836 vdd.n1412 vdd.n1411 0.00326471
R5837 vdd.n1426 vdd.n1415 0.00326471
R5838 vdd.n1580 vdd.n1579 0.00326471
R5839 vdd.n1603 vdd.n1602 0.00326471
R5840 vdd.n1629 vdd.n104 0.00326471
R5841 vdd.n1637 vdd.n1636 0.00326471
R5842 vdd.n1664 vdd.n1663 0.00326471
R5843 vdd.n1695 vdd.n1694 0.00326471
R5844 vdd.n1718 vdd.n1717 0.00326471
R5845 vdd.n1744 vdd.n40 0.00326471
R5846 vdd.n1752 vdd.n1751 0.00326471
R5847 vdd.n1775 vdd.n1774 0.00326471
R5848 vdd.n1862 vdd.n1861 0.00326471
R5849 vdd.n2953 vdd.n2952 0.00326471
R5850 vdd.n2961 vdd.n2383 0.00326471
R5851 vdd.n2991 vdd.n2369 0.00326471
R5852 vdd.n2999 vdd.n2998 0.00326471
R5853 vdd.n3020 vdd.n3019 0.00326471
R5854 vdd.n3044 vdd.n3043 0.00326471
R5855 vdd.n3179 vdd.n3178 0.00326471
R5856 vdd.n3187 vdd.n2249 0.00326471
R5857 vdd.n3217 vdd.n2235 0.00326471
R5858 vdd.n3225 vdd.n3224 0.00326471
R5859 vdd.n3246 vdd.n3245 0.00326471
R5860 vdd.n3270 vdd.n3269 0.00326471
R5861 vdd.n3405 vdd.n3404 0.00326471
R5862 vdd.n3413 vdd.n2115 0.00326471
R5863 vdd.n3443 vdd.n2101 0.00326471
R5864 vdd.n3451 vdd.n3450 0.00326471
R5865 vdd.n3472 vdd.n3471 0.00326471
R5866 vdd.n3496 vdd.n3495 0.00326471
R5867 vdd.n3631 vdd.n3630 0.00326471
R5868 vdd.n3639 vdd.n1981 0.00326471
R5869 vdd.n3669 vdd.n1967 0.00326471
R5870 vdd.n3677 vdd.n3676 0.00326471
R5871 vdd.n3702 vdd.n3701 0.00326471
R5872 vdd.n3730 vdd.n3729 0.00326471
R5873 vdd.n3749 vdd.n3748 0.00326471
R5874 vdd.n3768 vdd.n3767 0.00326471
R5875 vdd.n3787 vdd.n3786 0.00326471
R5876 vdd.n3806 vdd.n3805 0.00326471
R5877 vdd.n3827 vdd.n3826 0.00326471
R5878 vdd.n675 vdd.n674 0.00292718
R5879 vdd.n715 vdd.n602 0.00257353
R5880 vdd.n735 vdd.n589 0.00257353
R5881 vdd.n587 vdd.n575 0.00257353
R5882 vdd.n768 vdd.n573 0.00257353
R5883 vdd.n794 vdd.n556 0.00257353
R5884 vdd.n923 vdd.n919 0.00257353
R5885 vdd.n966 vdd.n468 0.00257353
R5886 vdd.n986 vdd.n455 0.00257353
R5887 vdd.n453 vdd.n441 0.00257353
R5888 vdd.n1019 vdd.n439 0.00257353
R5889 vdd.n1045 vdd.n422 0.00257353
R5890 vdd.n1174 vdd.n1170 0.00257353
R5891 vdd.n1217 vdd.n334 0.00257353
R5892 vdd.n1237 vdd.n321 0.00257353
R5893 vdd.n319 vdd.n307 0.00257353
R5894 vdd.n1270 vdd.n305 0.00257353
R5895 vdd.n1296 vdd.n288 0.00257353
R5896 vdd.n1425 vdd.n1421 0.00257353
R5897 vdd.n1468 vdd.n200 0.00257353
R5898 vdd.n1488 vdd.n187 0.00257353
R5899 vdd.n185 vdd.n173 0.00257353
R5900 vdd.n1521 vdd.n171 0.00257353
R5901 vdd.n1547 vdd.n154 0.00257353
R5902 vdd.n2842 vdd.n2459 0.00257353
R5903 vdd.n2457 vdd.n2447 0.00257353
R5904 vdd.n2872 vdd.n2445 0.00257353
R5905 vdd.n2894 vdd.n2431 0.00257353
R5906 vdd.n2914 vdd.n2420 0.00257353
R5907 vdd.n3048 vdd.n2335 0.00257353
R5908 vdd.n3068 vdd.n2325 0.00257353
R5909 vdd.n2323 vdd.n2313 0.00257353
R5910 vdd.n3098 vdd.n2311 0.00257353
R5911 vdd.n3120 vdd.n2297 0.00257353
R5912 vdd.n3140 vdd.n2286 0.00257353
R5913 vdd.n3274 vdd.n2201 0.00257353
R5914 vdd.n3294 vdd.n2191 0.00257353
R5915 vdd.n2189 vdd.n2179 0.00257353
R5916 vdd.n3324 vdd.n2177 0.00257353
R5917 vdd.n3346 vdd.n2163 0.00257353
R5918 vdd.n3366 vdd.n2152 0.00257353
R5919 vdd.n3500 vdd.n2067 0.00257353
R5920 vdd.n3520 vdd.n2057 0.00257353
R5921 vdd.n2055 vdd.n2045 0.00257353
R5922 vdd.n3550 vdd.n2043 0.00257353
R5923 vdd.n3572 vdd.n2029 0.00257353
R5924 vdd.n3592 vdd.n2018 0.00257353
R5925 vdd.n701 vdd.n598 0.00239394
R5926 vdd.n593 vdd.n591 0.00239394
R5927 vdd.n744 vdd.n578 0.00239394
R5928 vdd.n774 vdd.n773 0.00239394
R5929 vdd.n783 vdd.n553 0.00239394
R5930 vdd.n808 vdd.n543 0.00239394
R5931 vdd.n819 vdd.n818 0.00239394
R5932 vdd.n846 vdd.n526 0.00239394
R5933 vdd.n859 vdd.n519 0.00239394
R5934 vdd.n883 vdd.n504 0.00239394
R5935 vdd.n905 vdd.n492 0.00239394
R5936 vdd.n932 vdd.n479 0.00239394
R5937 vdd.n952 vdd.n464 0.00239394
R5938 vdd.n459 vdd.n457 0.00239394
R5939 vdd.n995 vdd.n444 0.00239394
R5940 vdd.n1025 vdd.n1024 0.00239394
R5941 vdd.n1034 vdd.n419 0.00239394
R5942 vdd.n1059 vdd.n409 0.00239394
R5943 vdd.n1070 vdd.n1069 0.00239394
R5944 vdd.n1097 vdd.n392 0.00239394
R5945 vdd.n1110 vdd.n385 0.00239394
R5946 vdd.n1134 vdd.n370 0.00239394
R5947 vdd.n1156 vdd.n358 0.00239394
R5948 vdd.n1183 vdd.n345 0.00239394
R5949 vdd.n1203 vdd.n330 0.00239394
R5950 vdd.n325 vdd.n323 0.00239394
R5951 vdd.n1246 vdd.n310 0.00239394
R5952 vdd.n1276 vdd.n1275 0.00239394
R5953 vdd.n1285 vdd.n285 0.00239394
R5954 vdd.n1310 vdd.n275 0.00239394
R5955 vdd.n1321 vdd.n1320 0.00239394
R5956 vdd.n1348 vdd.n258 0.00239394
R5957 vdd.n1361 vdd.n251 0.00239394
R5958 vdd.n1385 vdd.n236 0.00239394
R5959 vdd.n1407 vdd.n224 0.00239394
R5960 vdd.n1434 vdd.n211 0.00239394
R5961 vdd.n1454 vdd.n196 0.00239394
R5962 vdd.n191 vdd.n189 0.00239394
R5963 vdd.n1497 vdd.n176 0.00239394
R5964 vdd.n1527 vdd.n1526 0.00239394
R5965 vdd.n1536 vdd.n151 0.00239394
R5966 vdd.n1561 vdd.n141 0.00239394
R5967 vdd.n1572 vdd.n1571 0.00239394
R5968 vdd.n1594 vdd.n125 0.00239394
R5969 vdd.n1607 vdd.n109 0.00239394
R5970 vdd.n1641 vdd.n97 0.00239394
R5971 vdd.n1652 vdd.n1651 0.00239394
R5972 vdd.n1681 vdd.n74 0.00239394
R5973 vdd.n702 vdd.n600 0.00239394
R5974 vdd.n712 vdd.n590 0.00239394
R5975 vdd.n743 vdd.n577 0.00239394
R5976 vdd.n772 vdd.n569 0.00239394
R5977 vdd.n784 vdd.n554 0.00239394
R5978 vdd.n810 vdd.n809 0.00239394
R5979 vdd.n820 vdd.n539 0.00239394
R5980 vdd.n833 vdd.n527 0.00239394
R5981 vdd.n858 vdd.n857 0.00239394
R5982 vdd.n882 vdd.n505 0.00239394
R5983 vdd.n904 vdd.n493 0.00239394
R5984 vdd.n931 vdd.n930 0.00239394
R5985 vdd.n953 vdd.n466 0.00239394
R5986 vdd.n963 vdd.n456 0.00239394
R5987 vdd.n994 vdd.n443 0.00239394
R5988 vdd.n1023 vdd.n435 0.00239394
R5989 vdd.n1035 vdd.n420 0.00239394
R5990 vdd.n1061 vdd.n1060 0.00239394
R5991 vdd.n1071 vdd.n405 0.00239394
R5992 vdd.n1084 vdd.n393 0.00239394
R5993 vdd.n1109 vdd.n1108 0.00239394
R5994 vdd.n1133 vdd.n371 0.00239394
R5995 vdd.n1155 vdd.n359 0.00239394
R5996 vdd.n1182 vdd.n1181 0.00239394
R5997 vdd.n1204 vdd.n332 0.00239394
R5998 vdd.n1214 vdd.n322 0.00239394
R5999 vdd.n1245 vdd.n309 0.00239394
R6000 vdd.n1274 vdd.n301 0.00239394
R6001 vdd.n1286 vdd.n286 0.00239394
R6002 vdd.n1312 vdd.n1311 0.00239394
R6003 vdd.n1322 vdd.n271 0.00239394
R6004 vdd.n1335 vdd.n259 0.00239394
R6005 vdd.n1360 vdd.n1359 0.00239394
R6006 vdd.n1384 vdd.n237 0.00239394
R6007 vdd.n1406 vdd.n225 0.00239394
R6008 vdd.n1433 vdd.n1432 0.00239394
R6009 vdd.n1455 vdd.n198 0.00239394
R6010 vdd.n1465 vdd.n188 0.00239394
R6011 vdd.n1496 vdd.n175 0.00239394
R6012 vdd.n1525 vdd.n167 0.00239394
R6013 vdd.n1537 vdd.n152 0.00239394
R6014 vdd.n1563 vdd.n1562 0.00239394
R6015 vdd.n1573 vdd.n137 0.00239394
R6016 vdd.n1595 vdd.n123 0.00239394
R6017 vdd.n1606 vdd.n107 0.00239394
R6018 vdd.n1620 vdd.n98 0.00239394
R6019 vdd.n1653 vdd.n89 0.00239394
R6020 vdd.n1666 vdd.n75 0.00239394
R6021 vdd.n1709 vdd.n61 0.00239394
R6022 vdd.n1722 vdd.n45 0.00239394
R6023 vdd.n1756 vdd.n33 0.00239394
R6024 vdd.n1767 vdd.n1766 0.00239394
R6025 vdd.n1852 vdd.n11 0.00239394
R6026 vdd.n1710 vdd.n59 0.00239394
R6027 vdd.n1721 vdd.n43 0.00239394
R6028 vdd.n1735 vdd.n34 0.00239394
R6029 vdd.n1768 vdd.n25 0.00239394
R6030 vdd.n1853 vdd.n9 0.00239394
R6031 vdd.n2830 vdd.n2461 0.00239394
R6032 vdd.n2851 vdd.n2450 0.00239394
R6033 vdd.n2878 vdd.n2877 0.00239394
R6034 vdd.n2886 vdd.n2428 0.00239394
R6035 vdd.n2906 vdd.n2417 0.00239394
R6036 vdd.n2925 vdd.n2404 0.00239394
R6037 vdd.n2936 vdd.n2395 0.00239394
R6038 vdd.n2389 vdd.n2380 0.00239394
R6039 vdd.n2971 vdd.n2374 0.00239394
R6040 vdd.n3003 vdd.n2360 0.00239394
R6041 vdd.n3012 vdd.n2355 0.00239394
R6042 vdd.n3036 vdd.n2342 0.00239394
R6043 vdd.n3056 vdd.n2327 0.00239394
R6044 vdd.n3077 vdd.n2316 0.00239394
R6045 vdd.n3104 vdd.n3103 0.00239394
R6046 vdd.n3112 vdd.n2294 0.00239394
R6047 vdd.n3132 vdd.n2283 0.00239394
R6048 vdd.n3151 vdd.n2270 0.00239394
R6049 vdd.n3162 vdd.n2261 0.00239394
R6050 vdd.n2255 vdd.n2246 0.00239394
R6051 vdd.n3197 vdd.n2240 0.00239394
R6052 vdd.n3229 vdd.n2226 0.00239394
R6053 vdd.n3238 vdd.n2221 0.00239394
R6054 vdd.n3262 vdd.n2208 0.00239394
R6055 vdd.n3282 vdd.n2193 0.00239394
R6056 vdd.n3303 vdd.n2182 0.00239394
R6057 vdd.n3330 vdd.n3329 0.00239394
R6058 vdd.n3338 vdd.n2160 0.00239394
R6059 vdd.n3358 vdd.n2149 0.00239394
R6060 vdd.n3377 vdd.n2136 0.00239394
R6061 vdd.n3388 vdd.n2127 0.00239394
R6062 vdd.n2121 vdd.n2112 0.00239394
R6063 vdd.n3423 vdd.n2106 0.00239394
R6064 vdd.n3455 vdd.n2092 0.00239394
R6065 vdd.n3464 vdd.n2087 0.00239394
R6066 vdd.n3488 vdd.n2074 0.00239394
R6067 vdd.n3508 vdd.n2059 0.00239394
R6068 vdd.n3529 vdd.n2048 0.00239394
R6069 vdd.n3556 vdd.n3555 0.00239394
R6070 vdd.n3564 vdd.n2026 0.00239394
R6071 vdd.n3584 vdd.n2015 0.00239394
R6072 vdd.n3603 vdd.n2002 0.00239394
R6073 vdd.n3614 vdd.n1993 0.00239394
R6074 vdd.n1987 vdd.n1978 0.00239394
R6075 vdd.n3649 vdd.n1972 0.00239394
R6076 vdd.n3681 vdd.n1958 0.00239394
R6077 vdd.n3690 vdd.n1953 0.00239394
R6078 vdd.n3713 vdd.n1939 0.00239394
R6079 vdd.n2829 vdd.n2460 0.00239394
R6080 vdd.n2850 vdd.n2449 0.00239394
R6081 vdd.n2876 vdd.n2441 0.00239394
R6082 vdd.n2887 vdd.n2429 0.00239394
R6083 vdd.n2907 vdd.n2418 0.00239394
R6084 vdd.n2926 vdd.n2402 0.00239394
R6085 vdd.n2935 vdd.n2396 0.00239394
R6086 vdd.n2387 vdd.n2381 0.00239394
R6087 vdd.n2970 vdd.n2372 0.00239394
R6088 vdd.n2982 vdd.n2361 0.00239394
R6089 vdd.n3013 vdd.n2353 0.00239394
R6090 vdd.n3037 vdd.n2340 0.00239394
R6091 vdd.n3055 vdd.n2326 0.00239394
R6092 vdd.n3076 vdd.n2315 0.00239394
R6093 vdd.n3102 vdd.n2307 0.00239394
R6094 vdd.n3113 vdd.n2295 0.00239394
R6095 vdd.n3133 vdd.n2284 0.00239394
R6096 vdd.n3152 vdd.n2268 0.00239394
R6097 vdd.n3161 vdd.n2262 0.00239394
R6098 vdd.n2253 vdd.n2247 0.00239394
R6099 vdd.n3196 vdd.n2238 0.00239394
R6100 vdd.n3208 vdd.n2227 0.00239394
R6101 vdd.n3239 vdd.n2219 0.00239394
R6102 vdd.n3263 vdd.n2206 0.00239394
R6103 vdd.n3281 vdd.n2192 0.00239394
R6104 vdd.n3302 vdd.n2181 0.00239394
R6105 vdd.n3328 vdd.n2173 0.00239394
R6106 vdd.n3339 vdd.n2161 0.00239394
R6107 vdd.n3359 vdd.n2150 0.00239394
R6108 vdd.n3378 vdd.n2134 0.00239394
R6109 vdd.n3387 vdd.n2128 0.00239394
R6110 vdd.n2119 vdd.n2113 0.00239394
R6111 vdd.n3422 vdd.n2104 0.00239394
R6112 vdd.n3434 vdd.n2093 0.00239394
R6113 vdd.n3465 vdd.n2085 0.00239394
R6114 vdd.n3489 vdd.n2072 0.00239394
R6115 vdd.n3507 vdd.n2058 0.00239394
R6116 vdd.n3528 vdd.n2047 0.00239394
R6117 vdd.n3554 vdd.n2039 0.00239394
R6118 vdd.n3565 vdd.n2027 0.00239394
R6119 vdd.n3585 vdd.n2016 0.00239394
R6120 vdd.n3604 vdd.n2000 0.00239394
R6121 vdd.n3613 vdd.n1994 0.00239394
R6122 vdd.n1985 vdd.n1979 0.00239394
R6123 vdd.n3648 vdd.n1970 0.00239394
R6124 vdd.n3660 vdd.n1959 0.00239394
R6125 vdd.n3691 vdd.n1951 0.00239394
R6126 vdd.n3704 vdd.n1940 0.00239394
R6127 vdd.n3741 vdd.n1929 0.00239394
R6128 vdd.n3760 vdd.n1918 0.00239394
R6129 vdd.n3779 vdd.n1907 0.00239394
R6130 vdd.n3798 vdd.n1896 0.00239394
R6131 vdd.n3817 vdd.n1881 0.00239394
R6132 vdd.n3742 vdd.n1927 0.00239394
R6133 vdd.n3761 vdd.n1916 0.00239394
R6134 vdd.n3780 vdd.n1905 0.00239394
R6135 vdd.n3799 vdd.n1894 0.00239394
R6136 vdd.n3818 vdd.n1879 0.00239394
R6137 vdd.n1860 vdd.n1859 0.00224074
R6138 vdd.n3825 vdd.n3824 0.00224074
R6139 vdd.n662 vdd.n648 0.0021514
R6140 vdd.n2745 vdd.n2741 0.0021514
R6141 vdd.n1865 vdd.n4 0.00213953
R6142 vdd.n3830 vdd.n1874 0.00213953
R6143 vdd.n1816 vdd.n1815 0.00196875
R6144 vdd.n1794 vdd.n1793 0.00196875
R6145 vdd.n2779 vdd.n2764 0.00196875
R6146 vdd.n2784 vdd.n2781 0.00196875
R6147 vdd vdd.n616 0.00170513
R6148 vdd.n922 vdd 0.00170513
R6149 vdd.n1173 vdd 0.00170513
R6150 vdd.n1424 vdd 0.00170513
R6151 vdd.n2821 vdd 0.00170513
R6152 vdd vdd.n2334 0.00170513
R6153 vdd vdd.n2200 0.00170513
R6154 vdd vdd.n2066 0.00170513
R6155 vdd.n2754 vdd.t62 0.00166424
R6156 vdd.n2685 vdd.n2684 0.00142251
R6157 vdd.n614 vdd.n605 0.00119118
R6158 vdd.n703 vdd.n605 0.00119118
R6159 vdd.n714 vdd.n603 0.00119118
R6160 vdd.n711 vdd.n603 0.00119118
R6161 vdd.n736 vdd.n586 0.00119118
R6162 vdd.n742 vdd.n586 0.00119118
R6163 vdd.n761 vdd.n760 0.00119118
R6164 vdd.n762 vdd.n761 0.00119118
R6165 vdd.n767 vdd.n559 0.00119118
R6166 vdd.n785 vdd.n559 0.00119118
R6167 vdd.n793 vdd.n557 0.00119118
R6168 vdd.n557 vdd.n546 0.00119118
R6169 vdd.n822 vdd.n821 0.00119118
R6170 vdd.n822 vdd.n535 0.00119118
R6171 vdd.n826 vdd.n825 0.00119118
R6172 vdd.n826 vdd.n524 0.00119118
R6173 vdd.n856 vdd.n855 0.00119118
R6174 vdd.n855 vdd.n509 0.00119118
R6175 vdd.n881 vdd.n880 0.00119118
R6176 vdd.n880 vdd.n496 0.00119118
R6177 vdd.n903 vdd.n902 0.00119118
R6178 vdd.n902 vdd.n490 0.00119118
R6179 vdd.n929 vdd.n928 0.00119118
R6180 vdd.n928 vdd.n488 0.00119118
R6181 vdd.n920 vdd.n471 0.00119118
R6182 vdd.n954 vdd.n471 0.00119118
R6183 vdd.n965 vdd.n469 0.00119118
R6184 vdd.n962 vdd.n469 0.00119118
R6185 vdd.n987 vdd.n452 0.00119118
R6186 vdd.n993 vdd.n452 0.00119118
R6187 vdd.n1012 vdd.n1011 0.00119118
R6188 vdd.n1013 vdd.n1012 0.00119118
R6189 vdd.n1018 vdd.n425 0.00119118
R6190 vdd.n1036 vdd.n425 0.00119118
R6191 vdd.n1044 vdd.n423 0.00119118
R6192 vdd.n423 vdd.n412 0.00119118
R6193 vdd.n1073 vdd.n1072 0.00119118
R6194 vdd.n1073 vdd.n401 0.00119118
R6195 vdd.n1077 vdd.n1076 0.00119118
R6196 vdd.n1077 vdd.n390 0.00119118
R6197 vdd.n1107 vdd.n1106 0.00119118
R6198 vdd.n1106 vdd.n375 0.00119118
R6199 vdd.n1132 vdd.n1131 0.00119118
R6200 vdd.n1131 vdd.n362 0.00119118
R6201 vdd.n1154 vdd.n1153 0.00119118
R6202 vdd.n1153 vdd.n356 0.00119118
R6203 vdd.n1180 vdd.n1179 0.00119118
R6204 vdd.n1179 vdd.n354 0.00119118
R6205 vdd.n1171 vdd.n337 0.00119118
R6206 vdd.n1205 vdd.n337 0.00119118
R6207 vdd.n1216 vdd.n335 0.00119118
R6208 vdd.n1213 vdd.n335 0.00119118
R6209 vdd.n1238 vdd.n318 0.00119118
R6210 vdd.n1244 vdd.n318 0.00119118
R6211 vdd.n1263 vdd.n1262 0.00119118
R6212 vdd.n1264 vdd.n1263 0.00119118
R6213 vdd.n1269 vdd.n291 0.00119118
R6214 vdd.n1287 vdd.n291 0.00119118
R6215 vdd.n1295 vdd.n289 0.00119118
R6216 vdd.n289 vdd.n278 0.00119118
R6217 vdd.n1324 vdd.n1323 0.00119118
R6218 vdd.n1324 vdd.n267 0.00119118
R6219 vdd.n1328 vdd.n1327 0.00119118
R6220 vdd.n1328 vdd.n256 0.00119118
R6221 vdd.n1358 vdd.n1357 0.00119118
R6222 vdd.n1357 vdd.n241 0.00119118
R6223 vdd.n1383 vdd.n1382 0.00119118
R6224 vdd.n1382 vdd.n228 0.00119118
R6225 vdd.n1405 vdd.n1404 0.00119118
R6226 vdd.n1404 vdd.n222 0.00119118
R6227 vdd.n1431 vdd.n1430 0.00119118
R6228 vdd.n1430 vdd.n220 0.00119118
R6229 vdd.n1422 vdd.n203 0.00119118
R6230 vdd.n1456 vdd.n203 0.00119118
R6231 vdd.n1467 vdd.n201 0.00119118
R6232 vdd.n1464 vdd.n201 0.00119118
R6233 vdd.n1489 vdd.n184 0.00119118
R6234 vdd.n1495 vdd.n184 0.00119118
R6235 vdd.n1514 vdd.n1513 0.00119118
R6236 vdd.n1515 vdd.n1514 0.00119118
R6237 vdd.n1520 vdd.n157 0.00119118
R6238 vdd.n1538 vdd.n157 0.00119118
R6239 vdd.n1546 vdd.n155 0.00119118
R6240 vdd.n155 vdd.n144 0.00119118
R6241 vdd.n1575 vdd.n1574 0.00119118
R6242 vdd.n1575 vdd.n134 0.00119118
R6243 vdd.n1597 vdd.n1596 0.00119118
R6244 vdd.n1597 vdd.n118 0.00119118
R6245 vdd.n119 vdd.n106 0.00119118
R6246 vdd.n1626 vdd.n106 0.00119118
R6247 vdd.n1632 vdd.n1631 0.00119118
R6248 vdd.n1632 vdd.n102 0.00119118
R6249 vdd.n1655 vdd.n1654 0.00119118
R6250 vdd.n1655 vdd.n85 0.00119118
R6251 vdd.n1659 vdd.n1658 0.00119118
R6252 vdd.n1659 vdd.n72 0.00119118
R6253 vdd.n1690 vdd.n1689 0.00119118
R6254 vdd.n1690 vdd.n70 0.00119118
R6255 vdd.n1712 vdd.n1711 0.00119118
R6256 vdd.n1712 vdd.n54 0.00119118
R6257 vdd.n55 vdd.n42 0.00119118
R6258 vdd.n1741 vdd.n42 0.00119118
R6259 vdd.n1747 vdd.n1746 0.00119118
R6260 vdd.n1747 vdd.n38 0.00119118
R6261 vdd.n1770 vdd.n1769 0.00119118
R6262 vdd.n1770 vdd.n22 0.00119118
R6263 vdd.n1855 vdd.n1854 0.00119118
R6264 vdd.n1855 vdd.n6 0.00119118
R6265 vdd.n2823 vdd.n2465 0.00119118
R6266 vdd.n2828 vdd.n2465 0.00119118
R6267 vdd.n2843 vdd.n2456 0.00119118
R6268 vdd.n2849 vdd.n2456 0.00119118
R6269 vdd.n2865 vdd.n2864 0.00119118
R6270 vdd.n2866 vdd.n2865 0.00119118
R6271 vdd.n2871 vdd.n2433 0.00119118
R6272 vdd.n2888 vdd.n2433 0.00119118
R6273 vdd.n2893 vdd.n2422 0.00119118
R6274 vdd.n2908 vdd.n2422 0.00119118
R6275 vdd.n2913 vdd.n2400 0.00119118
R6276 vdd.n2927 vdd.n2400 0.00119118
R6277 vdd.n2934 vdd.n2933 0.00119118
R6278 vdd.n2933 vdd.n2385 0.00119118
R6279 vdd.n2954 vdd.n2382 0.00119118
R6280 vdd.n2964 vdd.n2382 0.00119118
R6281 vdd.n2959 vdd.n2371 0.00119118
R6282 vdd.n2988 vdd.n2371 0.00119118
R6283 vdd.n2994 vdd.n2993 0.00119118
R6284 vdd.n2994 vdd.n2367 0.00119118
R6285 vdd.n3015 vdd.n3014 0.00119118
R6286 vdd.n3015 vdd.n2350 0.00119118
R6287 vdd.n3039 vdd.n3038 0.00119118
R6288 vdd.n3039 vdd.n2337 0.00119118
R6289 vdd.n3049 vdd.n2333 0.00119118
R6290 vdd.n3054 vdd.n2333 0.00119118
R6291 vdd.n3069 vdd.n2322 0.00119118
R6292 vdd.n3075 vdd.n2322 0.00119118
R6293 vdd.n3091 vdd.n3090 0.00119118
R6294 vdd.n3092 vdd.n3091 0.00119118
R6295 vdd.n3097 vdd.n2299 0.00119118
R6296 vdd.n3114 vdd.n2299 0.00119118
R6297 vdd.n3119 vdd.n2288 0.00119118
R6298 vdd.n3134 vdd.n2288 0.00119118
R6299 vdd.n3139 vdd.n2266 0.00119118
R6300 vdd.n3153 vdd.n2266 0.00119118
R6301 vdd.n3160 vdd.n3159 0.00119118
R6302 vdd.n3159 vdd.n2251 0.00119118
R6303 vdd.n3180 vdd.n2248 0.00119118
R6304 vdd.n3190 vdd.n2248 0.00119118
R6305 vdd.n3185 vdd.n2237 0.00119118
R6306 vdd.n3214 vdd.n2237 0.00119118
R6307 vdd.n3220 vdd.n3219 0.00119118
R6308 vdd.n3220 vdd.n2233 0.00119118
R6309 vdd.n3241 vdd.n3240 0.00119118
R6310 vdd.n3241 vdd.n2216 0.00119118
R6311 vdd.n3265 vdd.n3264 0.00119118
R6312 vdd.n3265 vdd.n2203 0.00119118
R6313 vdd.n3275 vdd.n2199 0.00119118
R6314 vdd.n3280 vdd.n2199 0.00119118
R6315 vdd.n3295 vdd.n2188 0.00119118
R6316 vdd.n3301 vdd.n2188 0.00119118
R6317 vdd.n3317 vdd.n3316 0.00119118
R6318 vdd.n3318 vdd.n3317 0.00119118
R6319 vdd.n3323 vdd.n2165 0.00119118
R6320 vdd.n3340 vdd.n2165 0.00119118
R6321 vdd.n3345 vdd.n2154 0.00119118
R6322 vdd.n3360 vdd.n2154 0.00119118
R6323 vdd.n3365 vdd.n2132 0.00119118
R6324 vdd.n3379 vdd.n2132 0.00119118
R6325 vdd.n3386 vdd.n3385 0.00119118
R6326 vdd.n3385 vdd.n2117 0.00119118
R6327 vdd.n3406 vdd.n2114 0.00119118
R6328 vdd.n3416 vdd.n2114 0.00119118
R6329 vdd.n3411 vdd.n2103 0.00119118
R6330 vdd.n3440 vdd.n2103 0.00119118
R6331 vdd.n3446 vdd.n3445 0.00119118
R6332 vdd.n3446 vdd.n2099 0.00119118
R6333 vdd.n3467 vdd.n3466 0.00119118
R6334 vdd.n3467 vdd.n2082 0.00119118
R6335 vdd.n3491 vdd.n3490 0.00119118
R6336 vdd.n3491 vdd.n2069 0.00119118
R6337 vdd.n3501 vdd.n2065 0.00119118
R6338 vdd.n3506 vdd.n2065 0.00119118
R6339 vdd.n3521 vdd.n2054 0.00119118
R6340 vdd.n3527 vdd.n2054 0.00119118
R6341 vdd.n3543 vdd.n3542 0.00119118
R6342 vdd.n3544 vdd.n3543 0.00119118
R6343 vdd.n3549 vdd.n2031 0.00119118
R6344 vdd.n3566 vdd.n2031 0.00119118
R6345 vdd.n3571 vdd.n2020 0.00119118
R6346 vdd.n3586 vdd.n2020 0.00119118
R6347 vdd.n3591 vdd.n1998 0.00119118
R6348 vdd.n3605 vdd.n1998 0.00119118
R6349 vdd.n3612 vdd.n3611 0.00119118
R6350 vdd.n3611 vdd.n1983 0.00119118
R6351 vdd.n3632 vdd.n1980 0.00119118
R6352 vdd.n3642 vdd.n1980 0.00119118
R6353 vdd.n3637 vdd.n1969 0.00119118
R6354 vdd.n3666 vdd.n1969 0.00119118
R6355 vdd.n3672 vdd.n3671 0.00119118
R6356 vdd.n3672 vdd.n1965 0.00119118
R6357 vdd.n3693 vdd.n3692 0.00119118
R6358 vdd.n3693 vdd.n1947 0.00119118
R6359 vdd.n3697 vdd.n3696 0.00119118
R6360 vdd.n3697 vdd.n1937 0.00119118
R6361 vdd.n3725 vdd.n3724 0.00119118
R6362 vdd.n3725 vdd.n1935 0.00119118
R6363 vdd.n3744 vdd.n3743 0.00119118
R6364 vdd.n3744 vdd.n1924 0.00119118
R6365 vdd.n3763 vdd.n3762 0.00119118
R6366 vdd.n3763 vdd.n1913 0.00119118
R6367 vdd.n3782 vdd.n3781 0.00119118
R6368 vdd.n3782 vdd.n1902 0.00119118
R6369 vdd.n3801 vdd.n3800 0.00119118
R6370 vdd.n3801 vdd.n1891 0.00119118
R6371 vdd.n3820 vdd.n3819 0.00119118
R6372 vdd.n3820 vdd.n1876 0.00119118
R6373 vdd.n655 vdd.n653 0.0011215
R6374 vdd.n2734 vdd.n2732 0.0011215
R6375 vdd.n613 vdd.n604 0.00110256
R6376 vdd.n708 vdd.n707 0.00110256
R6377 vdd.n738 vdd.n737 0.00110256
R6378 vdd.n576 vdd.n574 0.00110256
R6379 vdd.n766 vdd.n558 0.00110256
R6380 vdd.n792 vdd.n791 0.00110256
R6381 vdd.n824 vdd.n823 0.00110256
R6382 vdd.n827 vdd.n523 0.00110256
R6383 vdd.n854 vdd.n508 0.00110256
R6384 vdd.n879 vdd.n495 0.00110256
R6385 vdd.n901 vdd.n489 0.00110256
R6386 vdd.n927 vdd.n926 0.00110256
R6387 vdd.n921 vdd.n470 0.00110256
R6388 vdd.n959 vdd.n958 0.00110256
R6389 vdd.n989 vdd.n988 0.00110256
R6390 vdd.n442 vdd.n440 0.00110256
R6391 vdd.n1017 vdd.n424 0.00110256
R6392 vdd.n1043 vdd.n1042 0.00110256
R6393 vdd.n1075 vdd.n1074 0.00110256
R6394 vdd.n1078 vdd.n389 0.00110256
R6395 vdd.n1105 vdd.n374 0.00110256
R6396 vdd.n1130 vdd.n361 0.00110256
R6397 vdd.n1152 vdd.n355 0.00110256
R6398 vdd.n1178 vdd.n1177 0.00110256
R6399 vdd.n1172 vdd.n336 0.00110256
R6400 vdd.n1210 vdd.n1209 0.00110256
R6401 vdd.n1240 vdd.n1239 0.00110256
R6402 vdd.n308 vdd.n306 0.00110256
R6403 vdd.n1268 vdd.n290 0.00110256
R6404 vdd.n1294 vdd.n1293 0.00110256
R6405 vdd.n1326 vdd.n1325 0.00110256
R6406 vdd.n1329 vdd.n255 0.00110256
R6407 vdd.n1356 vdd.n240 0.00110256
R6408 vdd.n1381 vdd.n227 0.00110256
R6409 vdd.n1403 vdd.n221 0.00110256
R6410 vdd.n1429 vdd.n1428 0.00110256
R6411 vdd.n1423 vdd.n202 0.00110256
R6412 vdd.n1461 vdd.n1460 0.00110256
R6413 vdd.n1491 vdd.n1490 0.00110256
R6414 vdd.n174 vdd.n172 0.00110256
R6415 vdd.n1519 vdd.n156 0.00110256
R6416 vdd.n1545 vdd.n1544 0.00110256
R6417 vdd.n1577 vdd.n1576 0.00110256
R6418 vdd.n1599 vdd.n1598 0.00110256
R6419 vdd.n1627 vdd.n105 0.00110256
R6420 vdd.n1634 vdd.n1633 0.00110256
R6421 vdd.n1657 vdd.n1656 0.00110256
R6422 vdd.n1660 vdd.n71 0.00110256
R6423 vdd.n2825 vdd.n2824 0.00110256
R6424 vdd.n2845 vdd.n2844 0.00110256
R6425 vdd.n2448 vdd.n2446 0.00110256
R6426 vdd.n2870 vdd.n2432 0.00110256
R6427 vdd.n2892 vdd.n2421 0.00110256
R6428 vdd.n2912 vdd.n2399 0.00110256
R6429 vdd.n2932 vdd.n2931 0.00110256
R6430 vdd.n2963 vdd.n2957 0.00110256
R6431 vdd.n2989 vdd.n2370 0.00110256
R6432 vdd.n2996 vdd.n2995 0.00110256
R6433 vdd.n3017 vdd.n3016 0.00110256
R6434 vdd.n3041 vdd.n3040 0.00110256
R6435 vdd.n3051 vdd.n3050 0.00110256
R6436 vdd.n3071 vdd.n3070 0.00110256
R6437 vdd.n2314 vdd.n2312 0.00110256
R6438 vdd.n3096 vdd.n2298 0.00110256
R6439 vdd.n3118 vdd.n2287 0.00110256
R6440 vdd.n3138 vdd.n2265 0.00110256
R6441 vdd.n3158 vdd.n3157 0.00110256
R6442 vdd.n3189 vdd.n3183 0.00110256
R6443 vdd.n3215 vdd.n2236 0.00110256
R6444 vdd.n3222 vdd.n3221 0.00110256
R6445 vdd.n3243 vdd.n3242 0.00110256
R6446 vdd.n3267 vdd.n3266 0.00110256
R6447 vdd.n3277 vdd.n3276 0.00110256
R6448 vdd.n3297 vdd.n3296 0.00110256
R6449 vdd.n2180 vdd.n2178 0.00110256
R6450 vdd.n3322 vdd.n2164 0.00110256
R6451 vdd.n3344 vdd.n2153 0.00110256
R6452 vdd.n3364 vdd.n2131 0.00110256
R6453 vdd.n3384 vdd.n3383 0.00110256
R6454 vdd.n3415 vdd.n3409 0.00110256
R6455 vdd.n3441 vdd.n2102 0.00110256
R6456 vdd.n3448 vdd.n3447 0.00110256
R6457 vdd.n3469 vdd.n3468 0.00110256
R6458 vdd.n3493 vdd.n3492 0.00110256
R6459 vdd.n3503 vdd.n3502 0.00110256
R6460 vdd.n3523 vdd.n3522 0.00110256
R6461 vdd.n2046 vdd.n2044 0.00110256
R6462 vdd.n3548 vdd.n2030 0.00110256
R6463 vdd.n3570 vdd.n2019 0.00110256
R6464 vdd.n3590 vdd.n1997 0.00110256
R6465 vdd.n3610 vdd.n3609 0.00110256
R6466 vdd.n3641 vdd.n3635 0.00110256
R6467 vdd.n3667 vdd.n1968 0.00110256
R6468 vdd.n3674 vdd.n3673 0.00110256
R6469 vdd.n3695 vdd.n3694 0.00110256
R6470 vdd.n3698 vdd.n1936 0.00110256
R6471 vdd.n1692 vdd.n1691 0.00108025
R6472 vdd.n1714 vdd.n1713 0.00108025
R6473 vdd.n1742 vdd.n41 0.00108025
R6474 vdd.n1749 vdd.n1748 0.00108025
R6475 vdd.n1772 vdd.n1771 0.00108025
R6476 vdd.n1857 vdd.n1856 0.00108025
R6477 vdd.n3727 vdd.n3726 0.00108025
R6478 vdd.n3746 vdd.n3745 0.00108025
R6479 vdd.n3765 vdd.n3764 0.00108025
R6480 vdd.n3784 vdd.n3783 0.00108025
R6481 vdd.n3803 vdd.n3802 0.00108025
R6482 vdd.n3822 vdd.n3821 0.00108025
R6483 vdd.n2651 vdd.n2561 0.000961255
R6484 vdd.n2630 vdd.n2629 0.000961255
R6485 vdd.n2639 vdd.n2638 0.000961255
R6486 vdd.n2640 vdd.n2557 0.000961255
R6487 vdd.n2660 vdd.n2659 0.000961255
R6488 vdd.n2664 vdd.n2555 0.000961255
R6489 vdd.n2672 vdd.n2671 0.000961255
R6490 vdd.n2670 vdd.n2665 0.000961255
R6491 vdd.n2684 vdd.n2548 0.000961255
R6492 vdd.n2746 vdd.n2729 0.000957792
R6493 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[2].t2 140.387
R6494 async_setb_delay_ctrl_code[2].n2 async_setb_delay_ctrl_code[2].t1 140.34
R6495 async_setb_delay_ctrl_code[2].n1 async_setb_delay_ctrl_code[2].t0 140.34
R6496 async_setb_delay_ctrl_code[2].n0 async_setb_delay_ctrl_code[2].t3 140.34
R6497 async_setb_delay_ctrl_code[2].n2 async_setb_delay_ctrl_code[2] 2.83
R6498 async_setb_delay_ctrl_code[2].n1 async_setb_delay_ctrl_code[2] 0.285826
R6499 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[2].n0 0.264087
R6500 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[2].n1 0.0466957
R6501 async_setb_delay_ctrl_code[2].n0 async_setb_delay_ctrl_code[2] 0.0466957
R6502 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[2].n2 0.0022562
R6503 vss vss.n1625 1.2997e+06
R6504 vss.n232 vss 1.15644e+06
R6505 vss.n1627 vss.n1626 21533.3
R6506 vss vss.n231 735.562
R6507 vss.n1626 vss 735.562
R6508 vss.n1409 vss.n1408 709.212
R6509 vss.n201 vss.t55 641.946
R6510 vss.n31 vss.t80 641.946
R6511 vss.n1628 vss.n5 626.532
R6512 vss.n1629 vss.n1628 626.365
R6513 vss.t77 vss.t3 611.288
R6514 vss.t28 vss.t22 611.288
R6515 vss.n1628 vss.n4 569.942
R6516 vss.t11 vss.n1487 536.975
R6517 vss.n1012 vss.t59 534.08
R6518 vss.t62 vss.n1572 415.149
R6519 vss.n94 vss.t31 391.634
R6520 vss.n99 vss.t46 338.432
R6521 vss.n122 vss.t48 338.432
R6522 vss.n201 vss 320.974
R6523 vss.n31 vss 320.974
R6524 vss.n231 vss.n230 307.599
R6525 vss.n1626 vss.n75 307.599
R6526 vss.n479 vss.n478 292.964
R6527 vss.n148 vss.n147 292.5
R6528 vss.n149 vss.n148 292.5
R6529 vss.n142 vss.n141 292.5
R6530 vss.n141 vss.n140 292.5
R6531 vss.n138 vss.n137 292.5
R6532 vss.n137 vss.n136 292.5
R6533 vss.n133 vss.n132 292.5
R6534 vss.n132 vss.n131 292.5
R6535 vss.n252 vss.n251 292.5
R6536 vss.n251 vss.n250 292.5
R6537 vss.n256 vss.n255 292.5
R6538 vss.n255 vss.n254 292.5
R6539 vss.n262 vss.n261 292.5
R6540 vss.n263 vss.n262 292.5
R6541 vss.n266 vss.n265 292.5
R6542 vss.n265 vss.n264 292.5
R6543 vss.n119 vss.n118 292.5
R6544 vss.n118 vss.n117 292.5
R6545 vss.n115 vss.n114 292.5
R6546 vss.n114 vss.n113 292.5
R6547 vss.n104 vss.n103 292.5
R6548 vss.n103 vss.n102 292.5
R6549 vss.n234 vss.n233 292.5
R6550 vss.n233 vss.n232 292.5
R6551 vss.n203 vss.n202 292.5
R6552 vss.n202 vss.n201 292.5
R6553 vss.n1593 vss.n1592 292.5
R6554 vss.n287 vss.n286 292.5
R6555 vss.n286 vss.n285 292.5
R6556 vss.n301 vss.n300 292.5
R6557 vss.n300 vss.n299 292.5
R6558 vss.n307 vss.n306 292.5
R6559 vss.n306 vss.n305 292.5
R6560 vss.n312 vss.n311 292.5
R6561 vss.n333 vss.n332 292.5
R6562 vss.n329 vss.n328 292.5
R6563 vss.n361 vss.n360 292.5
R6564 vss.n357 vss.n356 292.5
R6565 vss.n373 vss.n372 292.5
R6566 vss.n378 vss.n377 292.5
R6567 vss.n386 vss.n385 292.5
R6568 vss.n381 vss.n380 292.5
R6569 vss.n82 vss.n81 292.5
R6570 vss.n89 vss.n88 292.5
R6571 vss.n1615 vss.n1614 292.5
R6572 vss.n400 vss.n399 292.5
R6573 vss.n403 vss.n402 292.5
R6574 vss.n409 vss.n408 292.5
R6575 vss.n418 vss.n417 292.5
R6576 vss.n1585 vss.n1584 292.5
R6577 vss.n1589 vss.n1588 292.5
R6578 vss.n1597 vss.n1596 292.5
R6579 vss.n486 vss.n485 292.5
R6580 vss.n482 vss.n481 292.5
R6581 vss.n33 vss.n32 292.5
R6582 vss.n32 vss.n31 292.5
R6583 vss.n264 vss.t78 280.175
R6584 vss.t5 vss.n149 280.175
R6585 vss.n1628 vss.t1 278.445
R6586 vss.t0 vss.n1627 247.989
R6587 vss vss.n263 241.969
R6588 vss.n232 vss 241.969
R6589 vss.n181 vss.n180 227.357
R6590 vss.n42 vss.n41 227.357
R6591 vss.n99 vss.t87 224.35
R6592 vss.n122 vss.t86 224.35
R6593 vss.n423 vss.t14 211.167
R6594 vss.n371 vss.t10 184.713
R6595 vss vss.t34 183.873
R6596 vss.n117 vss.t26 178.292
R6597 vss.n1464 vss.t2 178.026
R6598 vss.n1310 vss.t69 178.026
R6599 vss.n1429 vss.t40 178.026
R6600 vss.n1219 vss.t42 178.026
R6601 vss.n853 vss.t41 178.026
R6602 vss.n962 vss.t39 178.026
R6603 vss.t59 vss.n948 178.026
R6604 vss.n1549 vss.t11 177.907
R6605 vss.n229 vss.n228 173.861
R6606 vss.n74 vss.n73 173.861
R6607 vss.n140 vss.t60 171.925
R6608 vss.t64 vss.t21 152.269
R6609 vss.n228 vss.t50 147.113
R6610 vss.n73 vss.t83 147.113
R6611 vss.n113 vss.t47 146.454
R6612 vss.n136 vss.t49 146.454
R6613 vss.n307 vss.t58 141.861
R6614 vss.t34 vss.t35 137.905
R6615 vss.n349 vss.n348 132.159
R6616 vss.n77 vss.n76 132.159
R6617 vss.n79 vss.n78 132.159
R6618 vss.t35 vss.t62 132.159
R6619 vss.n351 vss.t72 130.722
R6620 vss.n1577 vss.n1576 130.722
R6621 vss.t37 vss.n1574 126.412
R6622 vss.n348 vss.t9 124.977
R6623 vss.t73 vss.n346 119.231
R6624 vss.n350 vss.t29 119.231
R6625 vss.t75 vss.n1622 114.921
R6626 vss.n327 vss.n326 113.207
R6627 vss.n203 vss.t56 107.195
R6628 vss.n33 vss.t81 107.195
R6629 vss.n223 vss.t51 107.195
R6630 vss.n1591 vss.t38 107.195
R6631 vss.n480 vss.t45 107.195
R6632 vss.n68 vss.t84 107.195
R6633 vss.t12 vss.n1623 106.302
R6634 vss.n87 vss.n86 106.038
R6635 vss.n421 vss.n420 105.3
R6636 vss.t1 vss.t0 104.418
R6637 vss.n260 vss.n259 103.942
R6638 vss.n281 vss.n280 103.942
R6639 vss.n407 vss.n406 103.942
R6640 vss.n146 vss.n145 103.942
R6641 vss.n1579 vss.n1578 99.119
R6642 vss.n95 vss.t4 94.2521
R6643 vss.n125 vss.t23 94.1942
R6644 vss.t7 vss.n345 93.373
R6645 vss.n182 vss.n179 93.0283
R6646 vss.n43 vss.n40 93.0283
R6647 vss.t30 vss.n79 89.0635
R6648 vss.t85 vss.n80 77.5715
R6649 vss.n462 vss.t36 77.3934
R6650 vss.n462 vss.t33 77.3934
R6651 vss.n491 vss.t44 77.3934
R6652 vss.n491 vss.t43 77.3934
R6653 vss.n326 vss.t8 75.7148
R6654 vss.n259 vss.t27 74.2862
R6655 vss.n145 vss.t61 74.2862
R6656 vss.n1580 vss.t16 73.262
R6657 vss.n125 vss.t67 71.5727
R6658 vss.n95 vss.t32 71.5126
R6659 vss.n227 vss.n151 71.1394
R6660 vss.n72 vss.n7 71.1394
R6661 vss.n344 vss.t57 68.9525
R6662 vss.t52 vss.n1579 68.9525
R6663 vss.t21 vss.n344 67.516
R6664 vss.n1625 vss.t20 64.643
R6665 vss.n102 vss.t77 63.6763
R6666 vss.t78 vss 63.6763
R6667 vss.n131 vss.t28 63.6763
R6668 vss vss.t5 63.6763
R6669 vss.n285 vss.t70 63.2065
R6670 vss.n1580 vss.t52 63.2065
R6671 vss.n100 vss 62.5322
R6672 vss.n123 vss 62.5149
R6673 vss.t16 vss.n423 58.897
R6674 vss.n285 vss.t18 57.4605
R6675 vss.n1622 vss.t85 54.5875
R6676 vss.n406 vss.t25 54.2862
R6677 vss.n420 vss.t17 54.2862
R6678 vss.n230 vss.n229 53.4959
R6679 vss.n75 vss.n74 53.4959
R6680 vss.t14 vss.n422 53.151
R6681 vss.n78 vss.t24 48.8415
R6682 vss.n1625 vss.n1624 45.9685
R6683 vss.n345 vss.t64 44.532
R6684 vss.n473 vss.t68 43.7547
R6685 vss.n502 vss.t63 43.7547
R6686 vss.t70 vss 43.0955
R6687 vss.n80 vss.t30 43.0955
R6688 vss.n1629 vss.t82 41.4448
R6689 vss.n5 vss.t54 41.4448
R6690 vss.n86 vss.t13 41.4291
R6691 vss.n346 vss.t7 38.786
R6692 vss.n280 vss.t71 38.5719
R6693 vss.n280 vss.t19 38.5719
R6694 vss.n326 vss.t74 38.5719
R6695 vss.n86 vss.t76 38.5719
R6696 vss.n126 vss.n125 34.4596
R6697 vss.n96 vss.n95 34.4551
R6698 vss.n406 vss.t15 25.9346
R6699 vss.n420 vss.t53 25.9346
R6700 vss.n1624 vss.t12 25.8575
R6701 vss.n259 vss.t79 25.4291
R6702 vss.n145 vss.t6 25.4291
R6703 vss.n1573 vss 24.421
R6704 vss.n506 vss.n489 22.2971
R6705 vss.n151 vss.n150 21.8894
R6706 vss.n7 vss.n6 21.8894
R6707 vss.t20 vss.n77 21.548
R6708 vss vss.n99 18.19
R6709 vss vss.n122 18.19
R6710 vss.n1623 vss.t75 17.2385
R6711 vss.n477 vss.n397 17.0403
R6712 vss.n97 vss.n96 13.2928
R6713 vss.n204 vss.n203 13.1351
R6714 vss.n34 vss.n33 13.1351
R6715 vss.n127 vss.n126 13.042
R6716 vss.n351 vss.t73 12.929
R6717 vss.t29 vss.n349 12.929
R6718 vss vss.n281 12.8005
R6719 vss.n250 vss.t66 12.7357
R6720 vss vss.n284 10.4504
R6721 vss.n189 vss.n188 9.3005
R6722 vss.n187 vss.n186 9.3005
R6723 vss.n227 vss.n226 9.3005
R6724 vss.n228 vss.n227 9.3005
R6725 vss.n72 vss.n71 9.3005
R6726 vss.n73 vss.n72 9.3005
R6727 vss.n933 vss.n932 9.15497
R6728 vss.n932 vss.n931 9.15497
R6729 vss.n898 vss.n897 9.15497
R6730 vss.n897 vss.n4 9.15497
R6731 vss.n1069 vss.n1068 9.15497
R6732 vss.n1074 vss.n1073 9.15497
R6733 vss.n1073 vss.n4 9.15497
R6734 vss.n947 vss.n946 9.15497
R6735 vss.n948 vss.n947 9.15497
R6736 vss.n940 vss.n939 9.15497
R6737 vss.n939 vss.n938 9.15497
R6738 vss.n970 vss.n969 9.15497
R6739 vss.n976 vss.n975 9.15497
R6740 vss.n1011 vss.n1010 9.15497
R6741 vss.n1012 vss.n1011 9.15497
R6742 vss.n964 vss.n963 9.15497
R6743 vss.n963 vss.n962 9.15497
R6744 vss.n1116 vss.n1115 9.15497
R6745 vss.n1123 vss.n1122 9.15497
R6746 vss.n1122 vss.n1121 9.15497
R6747 vss.n1129 vss.n1128 9.15497
R6748 vss.n1110 vss.n1109 9.15497
R6749 vss.n1213 vss.n1212 9.15497
R6750 vss.n1190 vss.n1189 9.15497
R6751 vss.n1189 vss.n1188 9.15497
R6752 vss.n1173 vss.n1172 9.15497
R6753 vss.n1221 vss.n1220 9.15497
R6754 vss.n1220 vss.n1219 9.15497
R6755 vss.n1424 vss.n1423 9.15497
R6756 vss.n1423 vss.n1422 9.15497
R6757 vss.n1431 vss.n1430 9.15497
R6758 vss.n1430 vss.n1429 9.15497
R6759 vss.n1411 vss.n1410 9.15497
R6760 vss.n1410 vss.n1409 9.15497
R6761 vss.n1417 vss.n1416 9.15497
R6762 vss.n1365 vss.n1364 9.15497
R6763 vss.n1364 vss.n1363 9.15497
R6764 vss.n1372 vss.n1371 9.15497
R6765 vss.n1371 vss.n1370 9.15497
R6766 vss.n1407 vss.n1406 9.15497
R6767 vss.n1408 vss.n1407 9.15497
R6768 vss.n1358 vss.n1357 9.15497
R6769 vss.n1472 vss.n1471 9.15497
R6770 vss.n1466 vss.n1465 9.15497
R6771 vss.n1465 vss.n1464 9.15497
R6772 vss.n1486 vss.n1485 9.15497
R6773 vss.n1487 vss.n1486 9.15497
R6774 vss.n1479 vss.n1478 9.15497
R6775 vss.n1478 vss.n1477 9.15497
R6776 vss.n1057 vss.n1056 9.15497
R6777 vss.n1063 vss.n1062 9.15497
R6778 vss.n875 vss.n874 9.15497
R6779 vss.n874 vss.n873 9.15497
R6780 vss.n882 vss.n881 9.15497
R6781 vss.n881 vss.n880 9.15497
R6782 vss.n1014 vss.n1013 9.15497
R6783 vss.n1013 vss.n1012 9.15497
R6784 vss.n868 vss.n867 9.15497
R6785 vss.n842 vss.n841 9.15497
R6786 vss.n841 vss.n840 9.15497
R6787 vss.n848 vss.n847 9.15497
R6788 vss.n855 vss.n854 9.15497
R6789 vss.n854 vss.n853 9.15497
R6790 vss.n835 vss.n834 9.15497
R6791 vss.n834 vss.n833 9.15497
R6792 vss.n716 vss.n715 9.15497
R6793 vss.n715 vss.n714 9.15497
R6794 vss.n751 vss.n750 9.15497
R6795 vss.n789 vss.n788 9.15497
R6796 vss.n788 vss.n787 9.15497
R6797 vss.n723 vss.n722 9.15497
R6798 vss.n699 vss.n698 9.15497
R6799 vss.n705 vss.n704 9.15497
R6800 vss.n686 vss.n685 9.15497
R6801 vss.n693 vss.n692 9.15497
R6802 vss.n692 vss.n691 9.15497
R6803 vss.n1318 vss.n1317 9.15497
R6804 vss.n1324 vss.n1323 9.15497
R6805 vss.n1343 vss.n1342 9.15497
R6806 vss.n1408 vss.n1343 9.15497
R6807 vss.n1312 vss.n1311 9.15497
R6808 vss.n1311 vss.n1310 9.15497
R6809 vss.n1292 vss.n1291 9.15497
R6810 vss.n1291 vss.n1290 9.15497
R6811 vss.n1298 vss.n1297 9.15497
R6812 vss.n1279 vss.n1278 9.15497
R6813 vss.n1285 vss.n1284 9.15497
R6814 vss.n1502 vss.n1501 9.15497
R6815 vss.n1501 vss.n1500 9.15497
R6816 vss.n1548 vss.n1547 9.15497
R6817 vss.n1549 vss.n1548 9.15497
R6818 vss.n1489 vss.n1488 9.15497
R6819 vss.n1495 vss.n1494 9.15497
R6820 vss.n1557 vss.n1556 9.15497
R6821 vss.n1551 vss.n1550 9.15497
R6822 vss.n1550 vss.n1549 9.15497
R6823 vss.n1571 vss.n1570 9.15497
R6824 vss.n1572 vss.n1571 9.15497
R6825 vss.n1564 vss.n1563 9.15497
R6826 vss.n1563 vss.n1562 9.15497
R6827 vss.n183 vss.n182 9.01392
R6828 vss.n182 vss.n181 9.01392
R6829 vss.n1621 vss.n1620 9.01392
R6830 vss.n353 vss.n352 9.01392
R6831 vss.n284 vss.n283 9.01392
R6832 vss.n44 vss.n43 9.01392
R6833 vss.n43 vss.n42 9.01392
R6834 vss.n1582 vss.n1581 9.01392
R6835 vss.n1581 vss.n1580 9.01392
R6836 vss.n1622 vss.n1621 9.01392
R6837 vss.n352 vss.n351 9.01392
R6838 vss.n373 vss.n371 8.0005
R6839 vss.n203 vss 7.93155
R6840 vss.n33 vss 7.93155
R6841 vss.n224 vss.n223 7.52991
R6842 vss.n69 vss.n68 7.52991
R6843 vss.n329 vss.n327 7.28939
R6844 vss.n1593 vss.n1591 7.28939
R6845 vss.t9 vss.n347 7.183
R6846 vss.n89 vss.n87 6.93383
R6847 vss.n482 vss.n480 6.16917
R6848 vss.n484 vss.n482 4.80472
R6849 vss.n489 vss.n479 4.68956
R6850 vss.n205 vss.n204 4.6505
R6851 vss.n1616 vss.n1615 4.6505
R6852 vss.n1598 vss.n1597 4.6505
R6853 vss.n1590 vss.n1589 4.6505
R6854 vss.n1586 vss.n1585 4.6505
R6855 vss.n419 vss.n418 4.6505
R6856 vss.n416 vss.n415 4.6505
R6857 vss.n410 vss.n409 4.6505
R6858 vss.n404 vss.n403 4.6505
R6859 vss.n401 vss.n400 4.6505
R6860 vss.n1594 vss.n1593 4.6505
R6861 vss.n288 vss.n287 4.6505
R6862 vss.n302 vss.n301 4.6505
R6863 vss.n313 vss.n312 4.6505
R6864 vss.n308 vss.n307 4.6505
R6865 vss.n324 vss.n323 4.6505
R6866 vss.n334 vss.n333 4.6505
R6867 vss.n330 vss.n329 4.6505
R6868 vss.n362 vss.n361 4.6505
R6869 vss.n374 vss.n373 4.6505
R6870 vss.n358 vss.n357 4.6505
R6871 vss.n387 vss.n386 4.6505
R6872 vss.n379 vss.n378 4.6505
R6873 vss.n83 vss.n82 4.6505
R6874 vss.n382 vss.n381 4.6505
R6875 vss.n90 vss.n89 4.6505
R6876 vss.n488 vss.n487 4.6505
R6877 vss.n98 vss.n97 4.6505
R6878 vss.n101 vss.n100 4.6505
R6879 vss.n105 vss.n104 4.6505
R6880 vss.n116 vss.n115 4.6505
R6881 vss.n121 vss.n120 4.6505
R6882 vss.n267 vss.n266 4.6505
R6883 vss.n261 vss.n258 4.6505
R6884 vss.n257 vss.n256 4.6505
R6885 vss.n253 vss.n252 4.6505
R6886 vss.n128 vss.n127 4.6505
R6887 vss.n124 vss.n123 4.6505
R6888 vss.n235 vss.n234 4.6505
R6889 vss.n134 vss.n133 4.6505
R6890 vss.n139 vss.n138 4.6505
R6891 vss.n143 vss.n142 4.6505
R6892 vss.n147 vss.n144 4.6505
R6893 vss.n35 vss.n34 4.6505
R6894 vss.n222 vss.n221 4.5005
R6895 vss vss.n199 4.5005
R6896 vss vss.n30 4.5005
R6897 vss.n67 vss.n66 4.5005
R6898 vss.n1578 vss.n1577 4.31
R6899 vss.n1575 vss.t37 4.31
R6900 vss.n222 vss.n152 3.76521
R6901 vss.n67 vss.n10 3.76521
R6902 vss.n183 vss.n178 3.45447
R6903 vss.n44 vss.n39 3.45447
R6904 vss vss.n55 3.4105
R6905 vss.n225 vss.n224 3.38874
R6906 vss.n70 vss.n69 3.38874
R6907 vss.n184 vss.n177 3.25129
R6908 vss.n45 vss.n38 3.25129
R6909 vss.n283 vss 3.2005
R6910 vss.n237 vss.n236 3.1686
R6911 vss.n283 vss.n282 3.1005
R6912 vss.n1583 vss.n1582 3.1005
R6913 vss.n1620 vss.n1619 3.1005
R6914 vss.n354 vss.n353 3.1005
R6915 vss.n282 vss 3.09901
R6916 vss.n185 vss.n184 3.03311
R6917 vss.n1570 vss.n1569 3.03311
R6918 vss.n1490 vss.n1489 3.03311
R6919 vss.n1280 vss.n1279 3.03311
R6920 vss.n1319 vss.n1318 3.03311
R6921 vss.n1485 vss.n1484 3.03311
R6922 vss.n1366 vss.n1365 3.03311
R6923 vss.n687 vss.n686 3.03311
R6924 vss.n718 vss.n716 3.03311
R6925 vss.n843 vss.n842 3.03311
R6926 vss.n876 vss.n875 3.03311
R6927 vss.n1412 vss.n1411 3.03311
R6928 vss.n1215 vss.n1213 3.03311
R6929 vss.n1117 vss.n1116 3.03311
R6930 vss.n971 vss.n970 3.03311
R6931 vss.n1058 vss.n1057 3.03311
R6932 vss.n946 vss.n945 3.03311
R6933 vss.n934 vss.n933 3.03311
R6934 vss.n899 vss.n898 3.03311
R6935 vss.n1070 vss.n1069 3.03311
R6936 vss.n1075 vss.n1074 3.03311
R6937 vss.n941 vss.n940 3.03311
R6938 vss.n977 vss.n976 3.03311
R6939 vss.n1010 vss.n1009 3.03311
R6940 vss.n965 vss.n964 3.03311
R6941 vss.n1124 vss.n1123 3.03311
R6942 vss.n1130 vss.n1129 3.03311
R6943 vss.n1111 vss.n1110 3.03311
R6944 vss.n1191 vss.n1190 3.03311
R6945 vss.n1174 vss.n1173 3.03311
R6946 vss.n1222 vss.n1221 3.03311
R6947 vss.n1425 vss.n1424 3.03311
R6948 vss.n1432 vss.n1431 3.03311
R6949 vss.n1418 vss.n1417 3.03311
R6950 vss.n1373 vss.n1372 3.03311
R6951 vss.n1406 vss.n1405 3.03311
R6952 vss.n1359 vss.n1358 3.03311
R6953 vss.n1473 vss.n1472 3.03311
R6954 vss.n1467 vss.n1466 3.03311
R6955 vss.n1480 vss.n1479 3.03311
R6956 vss.n1064 vss.n1063 3.03311
R6957 vss.n883 vss.n882 3.03311
R6958 vss.n1015 vss.n1014 3.03311
R6959 vss.n869 vss.n868 3.03311
R6960 vss.n849 vss.n848 3.03311
R6961 vss.n856 vss.n855 3.03311
R6962 vss.n836 vss.n835 3.03311
R6963 vss.n752 vss.n751 3.03311
R6964 vss.n790 vss.n789 3.03311
R6965 vss.n724 vss.n723 3.03311
R6966 vss.n700 vss.n699 3.03311
R6967 vss.n706 vss.n705 3.03311
R6968 vss.n694 vss.n693 3.03311
R6969 vss.n1325 vss.n1324 3.03311
R6970 vss.n1342 vss.n1341 3.03311
R6971 vss.n1313 vss.n1312 3.03311
R6972 vss.n1293 vss.n1292 3.03311
R6973 vss.n1299 vss.n1298 3.03311
R6974 vss.n1286 vss.n1285 3.03311
R6975 vss.n1503 vss.n1502 3.03311
R6976 vss.n1547 vss.n1546 3.03311
R6977 vss.n1496 vss.n1495 3.03311
R6978 vss.n1558 vss.n1557 3.03311
R6979 vss.n1552 vss.n1551 3.03311
R6980 vss.n1565 vss.n1564 3.03311
R6981 vss.n46 vss.n45 3.03311
R6982 vss.n226 vss.n225 3.01226
R6983 vss.n71 vss.n70 3.01226
R6984 vss.n483 vss 3.0005
R6985 vss.n278 vss 2.98902
R6986 vss.n76 vss.t65 2.8735
R6987 vss.n303 vss 2.71795
R6988 vss.n98 vss.n94 2.68183
R6989 vss.n304 vss 2.63181
R6990 vss.n309 vss 2.47651
R6991 vss.n325 vss 2.41977
R6992 vss.n165 vss.n164 2.24031
R6993 vss.n343 vss 2.11899
R6994 vss.n355 vss 2.04132
R6995 vss.n166 vss 1.94963
R6996 vss.n1600 vss.n1599 1.94045
R6997 vss.n413 vss.n412 1.94045
R6998 vss.n290 vss.n289 1.94045
R6999 vss.n315 vss.n314 1.94045
R7000 vss.n336 vss.n335 1.94045
R7001 vss.n364 vss.n363 1.94045
R7002 vss.n389 vss.n388 1.94045
R7003 vss.n1613 vss.n1612 1.94045
R7004 vss.n107 vss.n106 1.94045
R7005 vss.n269 vss.n268 1.94045
R7006 vss.n249 vss.n248 1.94045
R7007 vss.n375 vss 1.63982
R7008 vss.n376 vss 1.58131
R7009 vss.n279 vss 1.57072
R7010 vss.n226 vss.n222 1.50638
R7011 vss.n9 vss.n8 1.50638
R7012 vss.n71 vss.n67 1.50638
R7013 vss.t72 vss.n350 1.437
R7014 vss.n1576 vss.n1575 1.437
R7015 vss.n1574 vss.n1573 1.437
R7016 vss.n383 vss 1.43106
R7017 vss.n310 vss 1.41264
R7018 vss.n219 vss.n218 1.35607
R7019 vss.n193 vss.n191 1.35607
R7020 vss.n64 vss.n63 1.35607
R7021 vss.n208 vss.n207 1.35607
R7022 vss.n1340 vss.n1339 1.35607
R7023 vss.n1404 vss.n1403 1.35607
R7024 vss.n1018 vss.n1016 1.35607
R7025 vss.n756 vss.n753 1.35607
R7026 vss.n793 vss.n791 1.35607
R7027 vss.n1008 vss.n1007 1.35607
R7028 vss.n1195 vss.n1192 1.35607
R7029 vss.n1177 vss.n1175 1.35607
R7030 vss.n1078 vss.n1076 1.35607
R7031 vss.n928 vss.n927 1.35607
R7032 vss.n29 vss.n24 1.35607
R7033 vss.n52 vss.n50 1.35607
R7034 vss.n331 vss 1.25121
R7035 vss.n84 vss 1.16066
R7036 vss.n504 vss.n503 1.13981
R7037 vss.n475 vss.n474 1.13981
R7038 vss.n170 vss.n169 1.13462
R7039 vss.n1639 vss.n1638 1.13462
R7040 vss.n10 vss.n9 1.12991
R7041 vss.n85 vss 1.10656
R7042 vss.n359 vss 1.10479
R7043 vss.n1582 vss.n421 1.06717
R7044 vss.n1634 vss.n1633 1.04173
R7045 vss.n1552 vss.n424 1.04008
R7046 vss.n1546 vss.n1545 1.04008
R7047 vss.n1300 vss.n1299 1.04008
R7048 vss.n1467 vss.n1463 1.04008
R7049 vss.n707 vss.n706 1.04008
R7050 vss.n857 vss.n856 1.04008
R7051 vss.n1433 vss.n1432 1.04008
R7052 vss.n1131 vss.n1130 1.04008
R7053 vss.n1313 vss.n1309 1.03985
R7054 vss.n1359 vss.n1356 1.03985
R7055 vss.n725 vss.n724 1.03985
R7056 vss.n869 vss.n866 1.03985
R7057 vss.n1223 vss.n1222 1.03985
R7058 vss.n965 vss.n961 1.03985
R7059 vss.n1058 vss.n1055 1.03984
R7060 vss.n945 vss.n896 1.03984
R7061 vss.n1617 vss 0.976265
R7062 vss.n409 vss.n407 0.889389
R7063 vss.n1637 vss.n1636 0.853
R7064 vss.n168 vss.n166 0.853
R7065 vss.n218 vss.n217 0.853
R7066 vss.n194 vss.n193 0.853
R7067 vss.n209 vss.n208 0.853
R7068 vss.n242 vss.n241 0.853
R7069 vss.n246 vss.n245 0.853
R7070 vss.n467 vss.n465 0.853
R7071 vss.n555 vss.n554 0.853
R7072 vss.n1544 vss.n1543 0.853
R7073 vss.n1339 vss.n583 0.853
R7074 vss.n1403 vss.n1402 0.853
R7075 vss.n1019 vss.n1018 0.853
R7076 vss.n1007 vss.n1006 0.853
R7077 vss.n1079 vss.n1078 0.853
R7078 vss.n927 vss.n926 0.853
R7079 vss.n895 vss.n894 0.853
R7080 vss.n1080 vss.n1079 0.853
R7081 vss.n1054 vss.n1053 0.853
R7082 vss.n589 vss.n588 0.853
R7083 vss.n960 vss.n959 0.853
R7084 vss.n1144 vss.n1143 0.853
R7085 vss.n1133 vss.n1104 0.853
R7086 vss.n1133 vss.n1132 0.853
R7087 vss.n1155 vss.n1154 0.853
R7088 vss.n1163 vss.n1162 0.853
R7089 vss.n1196 vss.n1195 0.853
R7090 vss.n1178 vss.n1177 0.853
R7091 vss.n1207 vss.n1206 0.853
R7092 vss.n1227 vss.n1226 0.853
R7093 vss.n611 vss.n610 0.853
R7094 vss.n1436 vss.n1435 0.853
R7095 vss.n1435 vss.n1434 0.853
R7096 vss.n600 vss.n599 0.853
R7097 vss.n1092 vss.n1019 0.853
R7098 vss.n654 vss.n653 0.853
R7099 vss.n865 vss.n864 0.853
R7100 vss.n824 vss.n823 0.853
R7101 vss.n859 vss.n858 0.853
R7102 vss.n813 vss.n812 0.853
R7103 vss.n802 vss.n801 0.853
R7104 vss.n757 vss.n756 0.853
R7105 vss.n794 vss.n782 0.853
R7106 vss.n794 vss.n793 0.853
R7107 vss.n740 vss.n739 0.853
R7108 vss.n729 vss.n728 0.853
R7109 vss.n676 vss.n675 0.853
R7110 vss.n709 vss.n708 0.853
R7111 vss.n665 vss.n664 0.853
R7112 vss.n433 vss.n432 0.853
R7113 vss.n1355 vss.n1354 0.853
R7114 vss.n455 vss.n454 0.853
R7115 vss.n1461 vss.n1460 0.853
R7116 vss.n1462 vss.n1461 0.853
R7117 vss.n444 vss.n443 0.853
R7118 vss.n1448 vss.n583 0.853
R7119 vss.n1247 vss.n1246 0.853
R7120 vss.n1308 vss.n1307 0.853
R7121 vss.n1269 vss.n1268 0.853
R7122 vss.n1302 vss.n1301 0.853
R7123 vss.n1258 vss.n1257 0.853
R7124 vss.n556 vss.n555 0.853
R7125 vss.n496 vss.n494 0.853
R7126 vss.n1610 vss.n1609 0.853
R7127 vss.n392 vss.n391 0.853
R7128 vss.n367 vss.n366 0.853
R7129 vss.n1606 vss.n396 0.853
R7130 vss.n1603 vss.n1602 0.853
R7131 vss.n339 vss.n338 0.853
R7132 vss.n318 vss.n317 0.853
R7133 vss.n293 vss.n292 0.853
R7134 vss.n273 vss.n272 0.853
R7135 vss.n110 vss.n109 0.853
R7136 vss.n63 vss.n61 0.853
R7137 vss.n29 vss.n28 0.853
R7138 vss.n53 vss.n52 0.853
R7139 vss.n384 vss 0.847393
R7140 vss.n216 vss.n215 0.699777
R7141 vss.n26 vss.n16 0.699777
R7142 vss.n211 vss.n210 0.699516
R7143 vss.n60 vss.n59 0.699516
R7144 vss.n469 vss.n468 0.698382
R7145 vss.n498 vss.n497 0.698382
R7146 vss.n474 vss.n473 0.684595
R7147 vss.n503 vss.n502 0.684595
R7148 vss.n248 vss.n247 0.682957
R7149 vss.n240 vss.n239 0.682957
R7150 vss.n108 vss.n107 0.682697
R7151 vss.n390 vss.n389 0.682668
R7152 vss.n365 vss.n364 0.682668
R7153 vss.n337 vss.n336 0.682668
R7154 vss.n316 vss.n315 0.682668
R7155 vss.n291 vss.n290 0.682668
R7156 vss.n412 vss.n411 0.682668
R7157 vss.n1601 vss.n1600 0.682668
R7158 vss.n1612 vss.n1611 0.682668
R7159 vss.n270 vss.n269 0.682657
R7160 vss.n1618 vss 0.59755
R7161 vss.n405 vss 0.59425
R7162 vss.n147 vss.n146 0.361063
R7163 vss.n287 vss.n281 0.356056
R7164 vss.n266 vss.n260 0.351185
R7165 vss.n470 vss.n469 0.319741
R7166 vss.n499 vss.n498 0.315296
R7167 vss.n1587 vss 0.30649
R7168 vss.n414 vss 0.254134
R7169 vss.n1305 vss.n1304 0.212
R7170 vss.n1352 vss.n1351 0.212
R7171 vss.n712 vss.n711 0.212
R7172 vss.n797 vss.n796 0.212
R7173 vss.n862 vss.n861 0.212
R7174 vss.n1230 vss.n1229 0.212
R7175 vss.n1166 vss.n1165 0.212
R7176 vss.n957 vss.n956 0.212
R7177 vss.n184 vss.n183 0.203675
R7178 vss.n45 vss.n44 0.203675
R7179 vss.n120 vss.n119 0.175842
R7180 vss.n212 vss.n172 0.170375
R7181 vss vss.n56 0.170375
R7182 vss.n487 vss.n486 0.154717
R7183 vss.n321 vss.n275 0.135899
R7184 vss.n419 vss.n416 0.120292
R7185 vss.n1583 vss.n419 0.120292
R7186 vss.n1586 vss.n1583 0.120292
R7187 vss.n404 vss.n401 0.120292
R7188 vss.n130 vss.n112 0.11645
R7189 vss.n1595 vss.n1594 0.107271
R7190 vss.n507 vss.n506 0.105976
R7191 vss.n507 vss.n477 0.105385
R7192 vss.n163 vss 0.104812
R7193 vss.n1617 vss.n1616 0.0981562
R7194 vss.n303 vss.n302 0.0981562
R7195 vss.n375 vss.n374 0.0981562
R7196 vss.n383 vss.n382 0.0981562
R7197 vss.n84 vss.n83 0.0981562
R7198 vss.n244 vss.n243 0.0971283
R7199 vss.n296 vss.n295 0.0959178
R7200 vss.n1595 vss 0.0935233
R7201 vss.n36 vss.n35 0.0929479
R7202 vss.n359 vss.n358 0.0877396
R7203 vss.n101 vss.n98 0.0798104
R7204 vss.n121 vss.n116 0.0798104
R7205 vss.n267 vss.n258 0.0798104
R7206 vss.n257 vss.n253 0.0798104
R7207 vss.n128 vss.n124 0.0798104
R7208 vss.n143 vss.n139 0.0798104
R7209 vss.n144 vss.n143 0.0798104
R7210 vss.n1605 vss.n1604 0.0761718
R7211 vss.n106 vss.n105 0.0737759
R7212 vss.n155 vss.n154 0.0734167
R7213 vss.n13 vss.n12 0.0734167
R7214 vss.n1567 vss.n1566 0.0685147
R7215 vss.n1560 vss.n1559 0.0685147
R7216 vss.n1554 vss.n1553 0.0685147
R7217 vss.n1493 vss.n1492 0.0685147
R7218 vss.n1499 vss.n1498 0.0685147
R7219 vss.n1506 vss.n1505 0.0685147
R7220 vss.n1283 vss.n1282 0.0685147
R7221 vss.n1289 vss.n1288 0.0685147
R7222 vss.n1296 vss.n1295 0.0685147
R7223 vss.n1315 vss.n1314 0.0685147
R7224 vss.n1321 vss.n1320 0.0685147
R7225 vss.n1327 vss.n1326 0.0685147
R7226 vss.n1482 vss.n1481 0.0685147
R7227 vss.n1475 vss.n1474 0.0685147
R7228 vss.n1469 vss.n1468 0.0685147
R7229 vss.n1361 vss.n1360 0.0685147
R7230 vss.n1368 vss.n1367 0.0685147
R7231 vss.n1375 vss.n1374 0.0685147
R7232 vss.n690 vss.n689 0.0685147
R7233 vss.n697 vss.n696 0.0685147
R7234 vss.n703 vss.n702 0.0685147
R7235 vss.n721 vss.n720 0.0685147
R7236 vss.n839 vss.n838 0.0685147
R7237 vss.n846 vss.n845 0.0685147
R7238 vss.n852 vss.n851 0.0685147
R7239 vss.n871 vss.n870 0.0685147
R7240 vss.n878 vss.n877 0.0685147
R7241 vss.n885 vss.n884 0.0685147
R7242 vss.n1415 vss.n1414 0.0685147
R7243 vss.n1421 vss.n1420 0.0685147
R7244 vss.n1428 vss.n1427 0.0685147
R7245 vss.n1218 vss.n1217 0.0685147
R7246 vss.n1114 vss.n1113 0.0685147
R7247 vss.n1120 vss.n1119 0.0685147
R7248 vss.n1127 vss.n1126 0.0685147
R7249 vss.n967 vss.n966 0.0685147
R7250 vss.n973 vss.n972 0.0685147
R7251 vss.n979 vss.n978 0.0685147
R7252 vss.n1060 vss.n1059 0.0685147
R7253 vss.n1066 vss.n1065 0.0685147
R7254 vss.n1072 vss.n1071 0.0685147
R7255 vss.n944 vss.n943 0.0685147
R7256 vss.n937 vss.n936 0.0685147
R7257 vss.n930 vss.n929 0.0685147
R7258 vss.n56 vss 0.0678766
R7259 vss.n1608 vss.n1607 0.0658282
R7260 vss.n405 vss.n404 0.0656042
R7261 vss.n206 vss.n205 0.0643021
R7262 vss.n331 vss.n330 0.0643021
R7263 vss.n236 vss.n235 0.062569
R7264 vss vss.n1586 0.0603958
R7265 vss.n394 vss.n393 0.0578436
R7266 vss.n249 vss.n128 0.0565345
R7267 vss.n488 vss.n484 0.0557885
R7268 vss.n477 vss.n476 0.0550615
R7269 vss.n1630 vss 0.0548478
R7270 vss.n506 vss.n505 0.0544685
R7271 vss.n369 vss.n368 0.0527625
R7272 vss vss.n189 0.0512812
R7273 vss vss.n48 0.0512812
R7274 vss.n212 vss.n211 0.0498797
R7275 vss vss.n16 0.0498797
R7276 vss.n539 vss.n538 0.0482941
R7277 vss.n545 vss.n544 0.0482941
R7278 vss.n551 vss.n550 0.0482941
R7279 vss.n1511 vss.n1510 0.0482941
R7280 vss.n1517 vss.n1516 0.0482941
R7281 vss.n1523 vss.n1522 0.0482941
R7282 vss.n1253 vss.n1252 0.0482941
R7283 vss.n1264 vss.n1263 0.0482941
R7284 vss.n1275 vss.n1274 0.0482941
R7285 vss.n1240 vss.n1239 0.0482941
R7286 vss.n1330 vss.n1329 0.0482941
R7287 vss.n1336 vss.n1335 0.0482941
R7288 vss.n439 vss.n438 0.0482941
R7289 vss.n450 vss.n449 0.0482941
R7290 vss.n426 vss.n425 0.0482941
R7291 vss.n1348 vss.n1347 0.0482941
R7292 vss.n1378 vss.n1377 0.0482941
R7293 vss.n1384 vss.n1383 0.0482941
R7294 vss.n660 vss.n659 0.0482941
R7295 vss.n671 vss.n670 0.0482941
R7296 vss.n682 vss.n681 0.0482941
R7297 vss.n735 vss.n734 0.0482941
R7298 vss.n746 vss.n745 0.0482941
R7299 vss.n784 vss.n783 0.0482941
R7300 vss.n808 vss.n807 0.0482941
R7301 vss.n819 vss.n818 0.0482941
R7302 vss.n830 vss.n829 0.0482941
R7303 vss.n647 vss.n646 0.0482941
R7304 vss.n635 vss.n634 0.0482941
R7305 vss.n641 vss.n640 0.0482941
R7306 vss.n595 vss.n594 0.0482941
R7307 vss.n606 vss.n605 0.0482941
R7308 vss.n1233 vss.n1232 0.0482941
R7309 vss.n1202 vss.n1201 0.0482941
R7310 vss.n1184 vss.n1183 0.0482941
R7311 vss.n1169 vss.n1168 0.0482941
R7312 vss.n1150 vss.n1149 0.0482941
R7313 vss.n1139 vss.n1138 0.0482941
R7314 vss.n1106 vss.n1105 0.0482941
R7315 vss.n953 vss.n952 0.0482941
R7316 vss.n982 vss.n981 0.0482941
R7317 vss.n988 vss.n987 0.0482941
R7318 vss.n1049 vss.n1048 0.0482941
R7319 vss.n1037 vss.n1036 0.0482941
R7320 vss.n1043 vss.n1042 0.0482941
R7321 vss.n890 vss.n889 0.0482941
R7322 vss.n902 vss.n901 0.0482941
R7323 vss.n908 vss.n907 0.0482941
R7324 vss.n414 vss.n413 0.0455581
R7325 vss.n314 vss.n313 0.0440714
R7326 vss.n268 vss.n121 0.0436034
R7327 vss.n1636 vss.n1635 0.0434688
R7328 vss.n30 vss.n29 0.0427297
R7329 vss.n208 vss.n199 0.0427297
R7330 vss.n388 vss.n387 0.0426598
R7331 vss.n135 vss.n134 0.0418793
R7332 vss.n166 vss.n162 0.0415156
R7333 vss.n465 vss.n461 0.0415156
R7334 vss.n494 vss.n490 0.0415156
R7335 vss.n197 vss.n196 0.0411354
R7336 vss.n55 vss.n17 0.0411354
R7337 vss vss.n257 0.0392931
R7338 vss.n1568 vss.n1567 0.0391029
R7339 vss.n1566 vss.n1565 0.0391029
R7340 vss.n1561 vss.n1560 0.0391029
R7341 vss.n1559 vss.n1558 0.0391029
R7342 vss.n1555 vss.n1554 0.0391029
R7343 vss.n1553 vss.n1552 0.0391029
R7344 vss.n537 vss.n536 0.0391029
R7345 vss.n541 vss.n540 0.0391029
R7346 vss.n543 vss.n542 0.0391029
R7347 vss.n547 vss.n546 0.0391029
R7348 vss.n549 vss.n548 0.0391029
R7349 vss.n553 vss.n552 0.0391029
R7350 vss.n1492 vss.n1491 0.0391029
R7351 vss.n1496 vss.n1493 0.0391029
R7352 vss.n1498 vss.n1497 0.0391029
R7353 vss.n1503 vss.n1499 0.0391029
R7354 vss.n1505 vss.n1504 0.0391029
R7355 vss.n1546 vss.n1506 0.0391029
R7356 vss.n1509 vss.n1508 0.0391029
R7357 vss.n1513 vss.n1512 0.0391029
R7358 vss.n1515 vss.n1514 0.0391029
R7359 vss.n1519 vss.n1518 0.0391029
R7360 vss.n1521 vss.n1520 0.0391029
R7361 vss.n1525 vss.n1524 0.0391029
R7362 vss.n1282 vss.n1281 0.0391029
R7363 vss.n1286 vss.n1283 0.0391029
R7364 vss.n1288 vss.n1287 0.0391029
R7365 vss.n1293 vss.n1289 0.0391029
R7366 vss.n1295 vss.n1294 0.0391029
R7367 vss.n1299 vss.n1296 0.0391029
R7368 vss.n1246 vss.n1245 0.0391029
R7369 vss.n1255 vss.n1254 0.0391029
R7370 vss.n1257 vss.n1256 0.0391029
R7371 vss.n1266 vss.n1265 0.0391029
R7372 vss.n1268 vss.n1267 0.0391029
R7373 vss.n1277 vss.n1276 0.0391029
R7374 vss.n1314 vss.n1313 0.0391029
R7375 vss.n1316 vss.n1315 0.0391029
R7376 vss.n1320 vss.n1319 0.0391029
R7377 vss.n1322 vss.n1321 0.0391029
R7378 vss.n1326 vss.n1325 0.0391029
R7379 vss.n1340 vss.n1327 0.0391029
R7380 vss.n1242 vss.n1241 0.0391029
R7381 vss.n1238 vss.n1237 0.0391029
R7382 vss.n1332 vss.n1331 0.0391029
R7383 vss.n1334 vss.n1333 0.0391029
R7384 vss.n1339 vss.n1337 0.0391029
R7385 vss.n1483 vss.n1482 0.0391029
R7386 vss.n1481 vss.n1480 0.0391029
R7387 vss.n1476 vss.n1475 0.0391029
R7388 vss.n1474 vss.n1473 0.0391029
R7389 vss.n1470 vss.n1469 0.0391029
R7390 vss.n1468 vss.n1467 0.0391029
R7391 vss.n432 vss.n431 0.0391029
R7392 vss.n441 vss.n440 0.0391029
R7393 vss.n443 vss.n442 0.0391029
R7394 vss.n452 vss.n451 0.0391029
R7395 vss.n454 vss.n453 0.0391029
R7396 vss.n428 vss.n427 0.0391029
R7397 vss.n1360 vss.n1359 0.0391029
R7398 vss.n1362 vss.n1361 0.0391029
R7399 vss.n1367 vss.n1366 0.0391029
R7400 vss.n1369 vss.n1368 0.0391029
R7401 vss.n1374 vss.n1373 0.0391029
R7402 vss.n1404 vss.n1375 0.0391029
R7403 vss.n1350 vss.n1349 0.0391029
R7404 vss.n1346 vss.n1345 0.0391029
R7405 vss.n1380 vss.n1379 0.0391029
R7406 vss.n1382 vss.n1381 0.0391029
R7407 vss.n1403 vss.n1385 0.0391029
R7408 vss.n689 vss.n688 0.0391029
R7409 vss.n694 vss.n690 0.0391029
R7410 vss.n696 vss.n695 0.0391029
R7411 vss.n700 vss.n697 0.0391029
R7412 vss.n702 vss.n701 0.0391029
R7413 vss.n706 vss.n703 0.0391029
R7414 vss.n653 vss.n652 0.0391029
R7415 vss.n662 vss.n661 0.0391029
R7416 vss.n664 vss.n663 0.0391029
R7417 vss.n673 vss.n672 0.0391029
R7418 vss.n675 vss.n674 0.0391029
R7419 vss.n684 vss.n683 0.0391029
R7420 vss.n724 vss.n721 0.0391029
R7421 vss.n720 vss.n719 0.0391029
R7422 vss.n718 vss.n717 0.0391029
R7423 vss.n753 vss.n748 0.0391029
R7424 vss.n752 vss.n749 0.0391029
R7425 vss.n791 vss.n786 0.0391029
R7426 vss.n727 vss.n726 0.0391029
R7427 vss.n739 vss.n736 0.0391029
R7428 vss.n738 vss.n737 0.0391029
R7429 vss.n756 vss.n747 0.0391029
R7430 vss.n755 vss.n754 0.0391029
R7431 vss.n793 vss.n785 0.0391029
R7432 vss.n838 vss.n837 0.0391029
R7433 vss.n843 vss.n839 0.0391029
R7434 vss.n845 vss.n844 0.0391029
R7435 vss.n849 vss.n846 0.0391029
R7436 vss.n851 vss.n850 0.0391029
R7437 vss.n856 vss.n852 0.0391029
R7438 vss.n801 vss.n800 0.0391029
R7439 vss.n810 vss.n809 0.0391029
R7440 vss.n812 vss.n811 0.0391029
R7441 vss.n821 vss.n820 0.0391029
R7442 vss.n823 vss.n822 0.0391029
R7443 vss.n832 vss.n831 0.0391029
R7444 vss.n870 vss.n869 0.0391029
R7445 vss.n872 vss.n871 0.0391029
R7446 vss.n877 vss.n876 0.0391029
R7447 vss.n879 vss.n878 0.0391029
R7448 vss.n884 vss.n883 0.0391029
R7449 vss.n1016 vss.n885 0.0391029
R7450 vss.n649 vss.n648 0.0391029
R7451 vss.n645 vss.n644 0.0391029
R7452 vss.n637 vss.n636 0.0391029
R7453 vss.n639 vss.n638 0.0391029
R7454 vss.n1018 vss.n642 0.0391029
R7455 vss.n1414 vss.n1413 0.0391029
R7456 vss.n1418 vss.n1415 0.0391029
R7457 vss.n1420 vss.n1419 0.0391029
R7458 vss.n1425 vss.n1421 0.0391029
R7459 vss.n1427 vss.n1426 0.0391029
R7460 vss.n1432 vss.n1428 0.0391029
R7461 vss.n588 vss.n587 0.0391029
R7462 vss.n597 vss.n596 0.0391029
R7463 vss.n599 vss.n598 0.0391029
R7464 vss.n608 vss.n607 0.0391029
R7465 vss.n610 vss.n609 0.0391029
R7466 vss.n1235 vss.n1234 0.0391029
R7467 vss.n1222 vss.n1218 0.0391029
R7468 vss.n1217 vss.n1216 0.0391029
R7469 vss.n1215 vss.n1214 0.0391029
R7470 vss.n1192 vss.n1186 0.0391029
R7471 vss.n1191 vss.n1187 0.0391029
R7472 vss.n1175 vss.n1171 0.0391029
R7473 vss.n1225 vss.n1224 0.0391029
R7474 vss.n1206 vss.n1203 0.0391029
R7475 vss.n1205 vss.n1204 0.0391029
R7476 vss.n1195 vss.n1185 0.0391029
R7477 vss.n1194 vss.n1193 0.0391029
R7478 vss.n1177 vss.n1170 0.0391029
R7479 vss.n1113 vss.n1112 0.0391029
R7480 vss.n1117 vss.n1114 0.0391029
R7481 vss.n1119 vss.n1118 0.0391029
R7482 vss.n1124 vss.n1120 0.0391029
R7483 vss.n1126 vss.n1125 0.0391029
R7484 vss.n1130 vss.n1127 0.0391029
R7485 vss.n1162 vss.n1161 0.0391029
R7486 vss.n1152 vss.n1151 0.0391029
R7487 vss.n1154 vss.n1153 0.0391029
R7488 vss.n1141 vss.n1140 0.0391029
R7489 vss.n1143 vss.n1142 0.0391029
R7490 vss.n1108 vss.n1107 0.0391029
R7491 vss.n966 vss.n965 0.0391029
R7492 vss.n968 vss.n967 0.0391029
R7493 vss.n972 vss.n971 0.0391029
R7494 vss.n974 vss.n973 0.0391029
R7495 vss.n978 vss.n977 0.0391029
R7496 vss.n1008 vss.n979 0.0391029
R7497 vss.n955 vss.n954 0.0391029
R7498 vss.n951 vss.n950 0.0391029
R7499 vss.n984 vss.n983 0.0391029
R7500 vss.n986 vss.n985 0.0391029
R7501 vss.n1007 vss.n989 0.0391029
R7502 vss.n1059 vss.n1058 0.0391029
R7503 vss.n1061 vss.n1060 0.0391029
R7504 vss.n1065 vss.n1064 0.0391029
R7505 vss.n1067 vss.n1066 0.0391029
R7506 vss.n1071 vss.n1070 0.0391029
R7507 vss.n1076 vss.n1072 0.0391029
R7508 vss.n1051 vss.n1050 0.0391029
R7509 vss.n1047 vss.n1046 0.0391029
R7510 vss.n1039 vss.n1038 0.0391029
R7511 vss.n1041 vss.n1040 0.0391029
R7512 vss.n1078 vss.n1044 0.0391029
R7513 vss.n945 vss.n944 0.0391029
R7514 vss.n943 vss.n942 0.0391029
R7515 vss.n941 vss.n937 0.0391029
R7516 vss.n936 vss.n935 0.0391029
R7517 vss.n934 vss.n930 0.0391029
R7518 vss.n929 vss.n928 0.0391029
R7519 vss.n892 vss.n891 0.0391029
R7520 vss.n888 vss.n887 0.0391029
R7521 vss.n904 vss.n903 0.0391029
R7522 vss.n906 vss.n905 0.0391029
R7523 vss.n927 vss.n909 0.0391029
R7524 vss.n1619 vss.n1613 0.0385435
R7525 vss.n139 vss.n135 0.038431
R7526 vss.n1599 vss.n1598 0.0382907
R7527 vss.n325 vss.n324 0.0369583
R7528 vss.n268 vss.n267 0.0367069
R7529 vss.n215 vss.n214 0.0361962
R7530 vss.n59 vss.n58 0.0361962
R7531 vss.n174 vss.n173 0.035973
R7532 vss.n193 vss.n192 0.035973
R7533 vss.n22 vss.n21 0.035973
R7534 vss.n52 vss.n51 0.035973
R7535 vss.n416 vss.n414 0.0356562
R7536 vss.n1613 vss.n90 0.0338851
R7537 vss.n363 vss.n355 0.033784
R7538 vss.n207 vss 0.0330521
R7539 vss vss.n24 0.0330521
R7540 vss.n335 vss.n325 0.0326429
R7541 vss.n63 vss.n14 0.0325946
R7542 vss.n218 vss.n156 0.0325946
R7543 vss.n289 vss.n278 0.0321011
R7544 vss.n190 vss 0.03175
R7545 vss.n49 vss 0.03175
R7546 vss.n289 vss.n288 0.0313989
R7547 vss.n341 vss.n340 0.0313585
R7548 vss.n334 vss.n331 0.0312143
R7549 vss.n410 vss.n405 0.0310233
R7550 vss.n160 vss.n159 0.029875
R7551 vss.n19 vss.n18 0.029875
R7552 vss.n1599 vss.n1590 0.0295698
R7553 vss.n1631 vss 0.0285374
R7554 vss.n363 vss.n362 0.0278669
R7555 vss.n191 vss.n190 0.0278438
R7556 vss.n1587 vss 0.0278438
R7557 vss.n50 vss.n49 0.0278438
R7558 vss.n388 vss.n379 0.0263876
R7559 vss.n164 vss.n163 0.0257686
R7560 vss.n1633 vss.n1632 0.0241592
R7561 vss.n463 vss.n462 0.024008
R7562 vss.n492 vss.n491 0.024008
R7563 vss.n253 vss.n249 0.0237759
R7564 vss.n558 vss 0.022851
R7565 vss vss.n1090 0.0226702
R7566 vss vss.n1446 0.0226702
R7567 vss.n314 vss.n308 0.0226429
R7568 vss.n154 vss 0.0226354
R7569 vss.n1594 vss 0.0226354
R7570 vss.n12 vss 0.0226354
R7571 vss.n166 vss.n165 0.0223823
R7572 vss.n354 vss.n343 0.0221837
R7573 vss.n536 vss.n535 0.0219755
R7574 vss.n1508 vss.n1507 0.0219755
R7575 vss.n1246 vss.n1244 0.0219755
R7576 vss.n1339 vss.n1338 0.0219755
R7577 vss.n432 vss.n430 0.0219755
R7578 vss.n1403 vss.n1386 0.0219755
R7579 vss.n653 vss.n651 0.0219755
R7580 vss.n793 vss.n792 0.0219755
R7581 vss.n801 vss.n799 0.0219755
R7582 vss.n1018 vss.n1017 0.0219755
R7583 vss.n588 vss.n586 0.0219755
R7584 vss.n1177 vss.n1176 0.0219755
R7585 vss.n1162 vss.n1160 0.0219755
R7586 vss.n1007 vss.n990 0.0219755
R7587 vss.n1078 vss.n1077 0.0219755
R7588 vss.n927 vss.n910 0.0219755
R7589 vss.n185 vss.n176 0.0213333
R7590 vss.n46 vss.n37 0.0213333
R7591 vss.n310 vss.n309 0.020702
R7592 vss.n220 vss.n219 0.0200312
R7593 vss.n65 vss.n64 0.0200312
R7594 vss.n275 vss.n111 0.0198586
R7595 vss.n85 vss.n84 0.0194394
R7596 vss.n519 vss.n518 0.0191618
R7597 vss.n520 vss.n519 0.0191618
R7598 vss.n524 vss.n523 0.0191618
R7599 vss.n525 vss.n524 0.0191618
R7600 vss.n529 vss.n528 0.0191618
R7601 vss.n530 vss.n529 0.0191618
R7602 vss.n555 vss.n533 0.0191618
R7603 vss.n555 vss.n534 0.0191618
R7604 vss.n1527 vss.n1526 0.0191618
R7605 vss.n1528 vss.n1527 0.0191618
R7606 vss.n1532 vss.n1531 0.0191618
R7607 vss.n1533 vss.n1532 0.0191618
R7608 vss.n1537 vss.n1536 0.0191618
R7609 vss.n1538 vss.n1537 0.0191618
R7610 vss.n1543 vss.n1541 0.0191618
R7611 vss.n1543 vss.n1542 0.0191618
R7612 vss.n1247 vss.n1243 0.0191618
R7613 vss.n1248 vss.n1247 0.0191618
R7614 vss.n1258 vss.n1251 0.0191618
R7615 vss.n1259 vss.n1258 0.0191618
R7616 vss.n1269 vss.n1262 0.0191618
R7617 vss.n1270 vss.n1269 0.0191618
R7618 vss.n1302 vss.n1273 0.0191618
R7619 vss.n1303 vss.n1302 0.0191618
R7620 vss.n1307 vss.n1306 0.0191618
R7621 vss.n572 vss.n571 0.0191618
R7622 vss.n573 vss.n572 0.0191618
R7623 vss.n577 vss.n576 0.0191618
R7624 vss.n578 vss.n577 0.0191618
R7625 vss.n583 vss.n581 0.0191618
R7626 vss.n583 vss.n582 0.0191618
R7627 vss.n433 vss.n429 0.0191618
R7628 vss.n434 vss.n433 0.0191618
R7629 vss.n444 vss.n437 0.0191618
R7630 vss.n445 vss.n444 0.0191618
R7631 vss.n455 vss.n448 0.0191618
R7632 vss.n456 vss.n455 0.0191618
R7633 vss.n1461 vss.n459 0.0191618
R7634 vss.n1461 vss.n460 0.0191618
R7635 vss.n1354 vss.n1353 0.0191618
R7636 vss.n1391 vss.n1390 0.0191618
R7637 vss.n1392 vss.n1391 0.0191618
R7638 vss.n1396 vss.n1395 0.0191618
R7639 vss.n1397 vss.n1396 0.0191618
R7640 vss.n1402 vss.n1400 0.0191618
R7641 vss.n1402 vss.n1401 0.0191618
R7642 vss.n654 vss.n650 0.0191618
R7643 vss.n655 vss.n654 0.0191618
R7644 vss.n665 vss.n658 0.0191618
R7645 vss.n666 vss.n665 0.0191618
R7646 vss.n676 vss.n669 0.0191618
R7647 vss.n677 vss.n676 0.0191618
R7648 vss.n709 vss.n680 0.0191618
R7649 vss.n710 vss.n709 0.0191618
R7650 vss.n729 vss.n713 0.0191618
R7651 vss.n730 vss.n729 0.0191618
R7652 vss.n740 vss.n733 0.0191618
R7653 vss.n741 vss.n740 0.0191618
R7654 vss.n757 vss.n744 0.0191618
R7655 vss.n758 vss.n757 0.0191618
R7656 vss.n794 vss.n761 0.0191618
R7657 vss.n795 vss.n794 0.0191618
R7658 vss.n802 vss.n798 0.0191618
R7659 vss.n803 vss.n802 0.0191618
R7660 vss.n813 vss.n806 0.0191618
R7661 vss.n814 vss.n813 0.0191618
R7662 vss.n824 vss.n817 0.0191618
R7663 vss.n825 vss.n824 0.0191618
R7664 vss.n859 vss.n828 0.0191618
R7665 vss.n860 vss.n859 0.0191618
R7666 vss.n864 vss.n863 0.0191618
R7667 vss.n622 vss.n621 0.0191618
R7668 vss.n623 vss.n622 0.0191618
R7669 vss.n627 vss.n626 0.0191618
R7670 vss.n628 vss.n627 0.0191618
R7671 vss.n1019 vss.n631 0.0191618
R7672 vss.n1019 vss.n632 0.0191618
R7673 vss.n589 vss.n585 0.0191618
R7674 vss.n590 vss.n589 0.0191618
R7675 vss.n600 vss.n593 0.0191618
R7676 vss.n601 vss.n600 0.0191618
R7677 vss.n611 vss.n604 0.0191618
R7678 vss.n612 vss.n611 0.0191618
R7679 vss.n1435 vss.n615 0.0191618
R7680 vss.n1435 vss.n1231 0.0191618
R7681 vss.n1228 vss.n1227 0.0191618
R7682 vss.n1227 vss.n1211 0.0191618
R7683 vss.n1208 vss.n1207 0.0191618
R7684 vss.n1207 vss.n1200 0.0191618
R7685 vss.n1197 vss.n1196 0.0191618
R7686 vss.n1196 vss.n1182 0.0191618
R7687 vss.n1179 vss.n1178 0.0191618
R7688 vss.n1178 vss.n1167 0.0191618
R7689 vss.n1164 vss.n1163 0.0191618
R7690 vss.n1163 vss.n1159 0.0191618
R7691 vss.n1156 vss.n1155 0.0191618
R7692 vss.n1155 vss.n1148 0.0191618
R7693 vss.n1145 vss.n1144 0.0191618
R7694 vss.n1144 vss.n1137 0.0191618
R7695 vss.n1134 vss.n1133 0.0191618
R7696 vss.n1133 vss.n616 0.0191618
R7697 vss.n959 vss.n958 0.0191618
R7698 vss.n995 vss.n994 0.0191618
R7699 vss.n996 vss.n995 0.0191618
R7700 vss.n1000 vss.n999 0.0191618
R7701 vss.n1001 vss.n1000 0.0191618
R7702 vss.n1006 vss.n1004 0.0191618
R7703 vss.n1006 vss.n1005 0.0191618
R7704 vss.n1053 vss.n1052 0.0191618
R7705 vss.n1024 vss.n1023 0.0191618
R7706 vss.n1025 vss.n1024 0.0191618
R7707 vss.n1029 vss.n1028 0.0191618
R7708 vss.n1030 vss.n1029 0.0191618
R7709 vss.n1079 vss.n1033 0.0191618
R7710 vss.n1079 vss.n1034 0.0191618
R7711 vss.n894 vss.n893 0.0191618
R7712 vss.n915 vss.n914 0.0191618
R7713 vss.n916 vss.n915 0.0191618
R7714 vss.n920 vss.n919 0.0191618
R7715 vss.n921 vss.n920 0.0191618
R7716 vss.n926 vss.n924 0.0191618
R7717 vss.n926 vss.n925 0.0191618
R7718 vss.n362 vss.n359 0.0189911
R7719 vss.n213 vss.n212 0.0183481
R7720 vss.n214 vss.n213 0.0183481
R7721 vss.n57 vss 0.0183481
R7722 vss.n58 vss.n57 0.0183481
R7723 vss.n236 vss.n144 0.0177414
R7724 vss.n1632 vss.n1629 0.0173735
R7725 vss vss.n1 0.0172471
R7726 vss vss.n584 0.0172471
R7727 vss.n781 vss 0.0172471
R7728 vss.n1103 vss 0.0172471
R7729 vss.n1091 vss 0.0172471
R7730 vss.n1459 vss 0.0172471
R7731 vss.n1447 vss 0.0172471
R7732 vss.n508 vss.n507 0.0172471
R7733 vss vss.n557 0.0172471
R7734 vss.n489 vss.n488 0.016726
R7735 vss vss.n483 0.016726
R7736 vss.n391 vss.n370 0.0157892
R7737 vss.n366 vss.n342 0.0157892
R7738 vss.n338 vss.n322 0.0157892
R7739 vss.n317 vss.n298 0.0157892
R7740 vss.n292 vss.n277 0.0157892
R7741 vss.n396 vss.n395 0.0157892
R7742 vss.n1602 vss.n398 0.0157892
R7743 vss.n1610 vss.n91 0.0157892
R7744 vss.n384 vss.n383 0.0156515
R7745 vss.n1637 vss.n3 0.0156071
R7746 vss.n168 vss.n167 0.0156071
R7747 vss.n272 vss.n271 0.0156071
R7748 vss.n246 vss.n129 0.0156071
R7749 vss.n241 vss.n238 0.0156071
R7750 vss.n472 vss.n471 0.0156071
R7751 vss.n467 vss.n466 0.0156071
R7752 vss.n501 vss.n500 0.0156071
R7753 vss.n496 vss.n495 0.0156071
R7754 vss.n109 vss.n93 0.0156071
R7755 vss.n522 vss.n521 0.0143235
R7756 vss.n527 vss.n526 0.0143235
R7757 vss.n532 vss.n531 0.0143235
R7758 vss.n1530 vss.n1529 0.0143235
R7759 vss.n1535 vss.n1534 0.0143235
R7760 vss.n1540 vss.n1539 0.0143235
R7761 vss.n1250 vss.n1249 0.0143235
R7762 vss.n1261 vss.n1260 0.0143235
R7763 vss.n1272 vss.n1271 0.0143235
R7764 vss.n570 vss.n569 0.0143235
R7765 vss.n575 vss.n574 0.0143235
R7766 vss.n580 vss.n579 0.0143235
R7767 vss.n436 vss.n435 0.0143235
R7768 vss.n447 vss.n446 0.0143235
R7769 vss.n458 vss.n457 0.0143235
R7770 vss.n1389 vss.n1388 0.0143235
R7771 vss.n1394 vss.n1393 0.0143235
R7772 vss.n1399 vss.n1398 0.0143235
R7773 vss.n657 vss.n656 0.0143235
R7774 vss.n668 vss.n667 0.0143235
R7775 vss.n679 vss.n678 0.0143235
R7776 vss.n732 vss.n731 0.0143235
R7777 vss.n743 vss.n742 0.0143235
R7778 vss.n760 vss.n759 0.0143235
R7779 vss.n805 vss.n804 0.0143235
R7780 vss.n816 vss.n815 0.0143235
R7781 vss.n827 vss.n826 0.0143235
R7782 vss.n620 vss.n619 0.0143235
R7783 vss.n625 vss.n624 0.0143235
R7784 vss.n630 vss.n629 0.0143235
R7785 vss.n592 vss.n591 0.0143235
R7786 vss.n603 vss.n602 0.0143235
R7787 vss.n614 vss.n613 0.0143235
R7788 vss.n1210 vss.n1209 0.0143235
R7789 vss.n1199 vss.n1198 0.0143235
R7790 vss.n1181 vss.n1180 0.0143235
R7791 vss.n1158 vss.n1157 0.0143235
R7792 vss.n1147 vss.n1146 0.0143235
R7793 vss.n1136 vss.n1135 0.0143235
R7794 vss.n993 vss.n992 0.0143235
R7795 vss.n998 vss.n997 0.0143235
R7796 vss.n1003 vss.n1002 0.0143235
R7797 vss.n1022 vss.n1021 0.0143235
R7798 vss.n1027 vss.n1026 0.0143235
R7799 vss.n1032 vss.n1031 0.0143235
R7800 vss.n913 vss.n912 0.0143235
R7801 vss.n918 vss.n917 0.0143235
R7802 vss.n923 vss.n922 0.0143235
R7803 vss.n163 vss.n5 0.0142993
R7804 vss.n258 vss 0.0142931
R7805 vss.n235 vss 0.0142931
R7806 vss.n335 vss.n334 0.0140714
R7807 vss.n464 vss.n463 0.0137243
R7808 vss.n493 vss.n492 0.0137243
R7809 vss.n209 vss.n198 0.0137188
R7810 vss.n195 vss.n194 0.0137188
R7811 vss.n217 vss.n161 0.0137188
R7812 vss.n28 vss.n27 0.0137188
R7813 vss.n54 vss.n53 0.0137188
R7814 vss.n53 vss.n20 0.0137188
R7815 vss.n61 vss.n15 0.0137188
R7816 vss.n221 vss.n153 0.0135208
R7817 vss.n66 vss.n11 0.0135208
R7818 vss.n355 vss.n354 0.0132551
R7819 vss.n288 vss.n279 0.0131404
R7820 vss.n320 vss.n319 0.0127097
R7821 vss.n243 vss.n242 0.0126552
R7822 vss.n242 vss.n237 0.0126552
R7823 vss.n245 vss.n130 0.0126552
R7824 vss.n245 vss.n244 0.0126552
R7825 vss.n63 vss.n62 0.0123243
R7826 vss.n218 vss.n157 0.0123243
R7827 vss.n164 vss 0.0121822
R7828 vss.n538 vss.n537 0.0115294
R7829 vss.n544 vss.n543 0.0115294
R7830 vss.n550 vss.n549 0.0115294
R7831 vss.n1510 vss.n1509 0.0115294
R7832 vss.n1516 vss.n1515 0.0115294
R7833 vss.n1522 vss.n1521 0.0115294
R7834 vss.n1239 vss.n1238 0.0115294
R7835 vss.n1331 vss.n1330 0.0115294
R7836 vss.n1337 vss.n1336 0.0115294
R7837 vss.n1347 vss.n1346 0.0115294
R7838 vss.n1379 vss.n1378 0.0115294
R7839 vss.n1385 vss.n1384 0.0115294
R7840 vss.n736 vss.n735 0.0115294
R7841 vss.n747 vss.n746 0.0115294
R7842 vss.n785 vss.n784 0.0115294
R7843 vss.n646 vss.n645 0.0115294
R7844 vss.n636 vss.n635 0.0115294
R7845 vss.n642 vss.n641 0.0115294
R7846 vss.n1203 vss.n1202 0.0115294
R7847 vss.n1185 vss.n1184 0.0115294
R7848 vss.n1170 vss.n1169 0.0115294
R7849 vss.n952 vss.n951 0.0115294
R7850 vss.n983 vss.n982 0.0115294
R7851 vss.n989 vss.n988 0.0115294
R7852 vss.n1048 vss.n1047 0.0115294
R7853 vss.n1038 vss.n1037 0.0115294
R7854 vss.n1044 vss.n1043 0.0115294
R7855 vss.n889 vss.n888 0.0115294
R7856 vss.n903 vss.n902 0.0115294
R7857 vss.n909 vss.n908 0.0115294
R7858 vss.n1631 vss.n1630 0.0113696
R7859 vss.n762 vss 0.0113046
R7860 vss vss.n780 0.0113046
R7861 vss vss.n1102 0.0113046
R7862 vss vss.n1458 0.0113046
R7863 vss.n297 vss.n296 0.0107238
R7864 vss.n484 vss 0.0107163
R7865 vss.n1636 vss.n1634 0.010716
R7866 vss.n1619 vss.n1618 0.0105932
R7867 vss.n308 vss.n304 0.0105
R7868 vss.n554 vss.n424 0.0104679
R7869 vss.n1545 vss.n1544 0.0104679
R7870 vss.n1301 vss.n1300 0.0104679
R7871 vss.n1463 vss.n1462 0.0104679
R7872 vss.n708 vss.n707 0.0104679
R7873 vss.n858 vss.n857 0.0104679
R7874 vss.n1434 vss.n1433 0.0104679
R7875 vss.n1132 vss.n1131 0.0104679
R7876 vss.n273 vss.n112 0.0102618
R7877 vss.n172 vss 0.01025
R7878 vss.n1055 vss.n1054 0.0100486
R7879 vss.n896 vss.n895 0.0100486
R7880 vss.n1309 vss.n1308 0.0098203
R7881 vss.n1356 vss.n1355 0.0098203
R7882 vss.n866 vss.n865 0.0098203
R7883 vss.n728 vss.n725 0.0098203
R7884 vss.n961 vss.n960 0.0098203
R7885 vss.n1226 vss.n1223 0.0098203
R7886 vss.n540 vss.n539 0.00969118
R7887 vss.n546 vss.n545 0.00969118
R7888 vss.n552 vss.n551 0.00969118
R7889 vss.n1512 vss.n1511 0.00969118
R7890 vss.n1518 vss.n1517 0.00969118
R7891 vss.n1524 vss.n1523 0.00969118
R7892 vss.n1254 vss.n1253 0.00969118
R7893 vss.n1265 vss.n1264 0.00969118
R7894 vss.n1276 vss.n1275 0.00969118
R7895 vss.n1241 vss.n1240 0.00969118
R7896 vss.n1329 vss.n1328 0.00969118
R7897 vss.n1335 vss.n1334 0.00969118
R7898 vss.n440 vss.n439 0.00969118
R7899 vss.n451 vss.n450 0.00969118
R7900 vss.n427 vss.n426 0.00969118
R7901 vss.n1349 vss.n1348 0.00969118
R7902 vss.n1377 vss.n1376 0.00969118
R7903 vss.n1383 vss.n1382 0.00969118
R7904 vss.n661 vss.n660 0.00969118
R7905 vss.n672 vss.n671 0.00969118
R7906 vss.n683 vss.n682 0.00969118
R7907 vss.n809 vss.n808 0.00969118
R7908 vss.n820 vss.n819 0.00969118
R7909 vss.n831 vss.n830 0.00969118
R7910 vss.n648 vss.n647 0.00969118
R7911 vss.n634 vss.n633 0.00969118
R7912 vss.n640 vss.n639 0.00969118
R7913 vss.n596 vss.n595 0.00969118
R7914 vss.n607 vss.n606 0.00969118
R7915 vss.n1234 vss.n1233 0.00969118
R7916 vss.n1151 vss.n1150 0.00969118
R7917 vss.n1140 vss.n1139 0.00969118
R7918 vss.n1107 vss.n1106 0.00969118
R7919 vss.n954 vss.n953 0.00969118
R7920 vss.n981 vss.n980 0.00969118
R7921 vss.n987 vss.n986 0.00969118
R7922 vss.n1050 vss.n1049 0.00969118
R7923 vss.n1036 vss.n1035 0.00969118
R7924 vss.n1042 vss.n1041 0.00969118
R7925 vss.n891 vss.n890 0.00969118
R7926 vss.n901 vss.n900 0.00969118
R7927 vss.n907 vss.n906 0.00969118
R7928 vss.n219 vss.n155 0.00961458
R7929 vss.n64 vss.n13 0.00961458
R7930 vss.n376 vss.n375 0.00933838
R7931 vss.n1632 vss.n1631 0.00809436
R7932 vss.n379 vss.n376 0.00789645
R7933 vss.n1598 vss.n1595 0.00776744
R7934 vss.n176 vss.n175 0.00701042
R7935 vss.n37 vss.n36 0.00701042
R7936 vss.n106 vss.n101 0.00653448
R7937 vss.n1638 vss.n1637 0.00635126
R7938 vss.n169 vss.n168 0.00635126
R7939 vss.n275 vss.n274 0.00608607
R7940 vss.n367 vss.n341 0.00594402
R7941 vss.n368 vss.n367 0.00594402
R7942 vss.n392 vss.n369 0.00594402
R7943 vss.n393 vss.n392 0.00594402
R7944 vss.n1609 vss.n394 0.00594402
R7945 vss.n1609 vss.n1608 0.00594402
R7946 vss.n1607 vss.n1606 0.00594402
R7947 vss.n1606 vss.n1605 0.00594402
R7948 vss.n1604 vss.n1603 0.00594402
R7949 vss.n1603 vss.n397 0.00594402
R7950 vss.n189 vss.n187 0.00570833
R7951 vss.n221 vss.n220 0.00570833
R7952 vss.n48 vss.n47 0.00570833
R7953 vss.n66 vss.n65 0.00570833
R7954 vss.n1618 vss.n1617 0.00560204
R7955 vss.n505 vss.n504 0.00494795
R7956 vss.n504 vss.n499 0.00494795
R7957 vss.n475 vss.n470 0.00494795
R7958 vss.n476 vss.n475 0.00494795
R7959 vss.n296 vss.n294 0.00491315
R7960 vss.n468 vss.n467 0.00489326
R7961 vss.n497 vss.n496 0.00489326
R7962 vss.n247 vss.n246 0.00486839
R7963 vss.n241 vss.n240 0.00486839
R7964 vss vss.n1640 0.00481329
R7965 vss.n217 vss.n216 0.00451955
R7966 vss.n28 vss.n26 0.00451955
R7967 vss.n187 vss.n153 0.00440625
R7968 vss.n47 vss.n11 0.00440625
R7969 vss.n282 vss.n278 0.00432653
R7970 vss.n304 vss.n303 0.00428788
R7971 vss.n387 vss.n384 0.00419822
R7972 vss.n272 vss.n270 0.00417181
R7973 vss.n1590 vss.n1587 0.00413372
R7974 vss.n391 vss.n390 0.0040098
R7975 vss.n366 vss.n365 0.0040098
R7976 vss.n338 vss.n337 0.0040098
R7977 vss.n317 vss.n316 0.0040098
R7978 vss.n292 vss.n291 0.0040098
R7979 vss.n411 vss.n396 0.0040098
R7980 vss.n1602 vss.n1601 0.0040098
R7981 vss.n1611 vss.n1610 0.0040098
R7982 vss.n109 vss.n108 0.00397409
R7983 vss.n210 vss.n209 0.00362372
R7984 vss.n61 vss.n60 0.00362372
R7985 vss.n110 vss.n92 0.00338934
R7986 vss.n111 vss.n110 0.00338934
R7987 vss.n274 vss.n273 0.00338934
R7988 vss.n1090 vss.n1089 0.00320115
R7989 vss.n1089 vss.n1088 0.00320115
R7990 vss.n1087 vss.n1086 0.00320115
R7991 vss.n1086 vss.n1085 0.00320115
R7992 vss.n1084 vss.n1083 0.00320115
R7993 vss.n1083 vss.n1082 0.00320115
R7994 vss.n1081 vss.n1080 0.00320115
R7995 vss.n1080 vss.n1 0.00320115
R7996 vss.n1446 vss.n1445 0.00320115
R7997 vss.n1445 vss.n1444 0.00320115
R7998 vss.n1443 vss.n1442 0.00320115
R7999 vss.n1442 vss.n1441 0.00320115
R8000 vss.n1440 vss.n1439 0.00320115
R8001 vss.n1439 vss.n1438 0.00320115
R8002 vss.n1437 vss.n1436 0.00320115
R8003 vss.n1436 vss.n584 0.00320115
R8004 vss.n763 vss.n762 0.00320115
R8005 vss.n764 vss.n763 0.00320115
R8006 vss.n766 vss.n765 0.00320115
R8007 vss.n767 vss.n766 0.00320115
R8008 vss.n769 vss.n768 0.00320115
R8009 vss.n770 vss.n769 0.00320115
R8010 vss.n782 vss.n771 0.00320115
R8011 vss.n782 vss.n781 0.00320115
R8012 vss.n780 vss.n779 0.00320115
R8013 vss.n779 vss.n778 0.00320115
R8014 vss.n777 vss.n776 0.00320115
R8015 vss.n776 vss.n775 0.00320115
R8016 vss.n774 vss.n773 0.00320115
R8017 vss.n773 vss.n772 0.00320115
R8018 vss.n1104 vss.n617 0.00320115
R8019 vss.n1104 vss.n1103 0.00320115
R8020 vss.n1102 vss.n1101 0.00320115
R8021 vss.n1101 vss.n1100 0.00320115
R8022 vss.n1099 vss.n1098 0.00320115
R8023 vss.n1098 vss.n1097 0.00320115
R8024 vss.n1096 vss.n1095 0.00320115
R8025 vss.n1095 vss.n1094 0.00320115
R8026 vss.n1093 vss.n1092 0.00320115
R8027 vss.n1092 vss.n1091 0.00320115
R8028 vss.n559 vss.n558 0.00320115
R8029 vss.n560 vss.n559 0.00320115
R8030 vss.n562 vss.n561 0.00320115
R8031 vss.n563 vss.n562 0.00320115
R8032 vss.n565 vss.n564 0.00320115
R8033 vss.n566 vss.n565 0.00320115
R8034 vss.n1460 vss.n567 0.00320115
R8035 vss.n1460 vss.n1459 0.00320115
R8036 vss.n1458 vss.n1457 0.00320115
R8037 vss.n1457 vss.n1456 0.00320115
R8038 vss.n1455 vss.n1454 0.00320115
R8039 vss.n1454 vss.n1453 0.00320115
R8040 vss.n1452 vss.n1451 0.00320115
R8041 vss.n1451 vss.n1450 0.00320115
R8042 vss.n1449 vss.n1448 0.00320115
R8043 vss.n1448 vss.n1447 0.00320115
R8044 vss.n509 vss.n508 0.00320115
R8045 vss.n510 vss.n509 0.00320115
R8046 vss.n512 vss.n511 0.00320115
R8047 vss.n513 vss.n512 0.00320115
R8048 vss.n515 vss.n514 0.00320115
R8049 vss.n516 vss.n515 0.00320115
R8050 vss.n556 vss.n517 0.00320115
R8051 vss.n557 vss.n556 0.00320115
R8052 vss.n293 vss.n276 0.00270657
R8053 vss.n294 vss.n293 0.00270657
R8054 vss.n318 vss.n297 0.00270657
R8055 vss.n319 vss.n318 0.00270657
R8056 vss.n340 vss.n339 0.00270657
R8057 vss.n413 vss.n410 0.00268023
R8058 vss.n521 vss.n520 0.00257353
R8059 vss.n523 vss.n522 0.00257353
R8060 vss.n526 vss.n525 0.00257353
R8061 vss.n528 vss.n527 0.00257353
R8062 vss.n531 vss.n530 0.00257353
R8063 vss.n533 vss.n532 0.00257353
R8064 vss.n1529 vss.n1528 0.00257353
R8065 vss.n1531 vss.n1530 0.00257353
R8066 vss.n1534 vss.n1533 0.00257353
R8067 vss.n1536 vss.n1535 0.00257353
R8068 vss.n1539 vss.n1538 0.00257353
R8069 vss.n1541 vss.n1540 0.00257353
R8070 vss.n1249 vss.n1248 0.00257353
R8071 vss.n1251 vss.n1250 0.00257353
R8072 vss.n1260 vss.n1259 0.00257353
R8073 vss.n1262 vss.n1261 0.00257353
R8074 vss.n1271 vss.n1270 0.00257353
R8075 vss.n1273 vss.n1272 0.00257353
R8076 vss.n1304 vss.n1303 0.00257353
R8077 vss.n1306 vss.n1305 0.00257353
R8078 vss.n569 vss.n568 0.00257353
R8079 vss.n571 vss.n570 0.00257353
R8080 vss.n574 vss.n573 0.00257353
R8081 vss.n576 vss.n575 0.00257353
R8082 vss.n579 vss.n578 0.00257353
R8083 vss.n581 vss.n580 0.00257353
R8084 vss.n435 vss.n434 0.00257353
R8085 vss.n437 vss.n436 0.00257353
R8086 vss.n446 vss.n445 0.00257353
R8087 vss.n448 vss.n447 0.00257353
R8088 vss.n457 vss.n456 0.00257353
R8089 vss.n459 vss.n458 0.00257353
R8090 vss.n1351 vss.n460 0.00257353
R8091 vss.n1353 vss.n1352 0.00257353
R8092 vss.n1388 vss.n1387 0.00257353
R8093 vss.n1390 vss.n1389 0.00257353
R8094 vss.n1393 vss.n1392 0.00257353
R8095 vss.n1395 vss.n1394 0.00257353
R8096 vss.n1398 vss.n1397 0.00257353
R8097 vss.n1400 vss.n1399 0.00257353
R8098 vss.n656 vss.n655 0.00257353
R8099 vss.n658 vss.n657 0.00257353
R8100 vss.n667 vss.n666 0.00257353
R8101 vss.n669 vss.n668 0.00257353
R8102 vss.n678 vss.n677 0.00257353
R8103 vss.n680 vss.n679 0.00257353
R8104 vss.n711 vss.n710 0.00257353
R8105 vss.n713 vss.n712 0.00257353
R8106 vss.n731 vss.n730 0.00257353
R8107 vss.n733 vss.n732 0.00257353
R8108 vss.n742 vss.n741 0.00257353
R8109 vss.n744 vss.n743 0.00257353
R8110 vss.n759 vss.n758 0.00257353
R8111 vss.n761 vss.n760 0.00257353
R8112 vss.n796 vss.n795 0.00257353
R8113 vss.n798 vss.n797 0.00257353
R8114 vss.n804 vss.n803 0.00257353
R8115 vss.n806 vss.n805 0.00257353
R8116 vss.n815 vss.n814 0.00257353
R8117 vss.n817 vss.n816 0.00257353
R8118 vss.n826 vss.n825 0.00257353
R8119 vss.n828 vss.n827 0.00257353
R8120 vss.n861 vss.n860 0.00257353
R8121 vss.n863 vss.n862 0.00257353
R8122 vss.n619 vss.n618 0.00257353
R8123 vss.n621 vss.n620 0.00257353
R8124 vss.n624 vss.n623 0.00257353
R8125 vss.n626 vss.n625 0.00257353
R8126 vss.n629 vss.n628 0.00257353
R8127 vss.n631 vss.n630 0.00257353
R8128 vss.n591 vss.n590 0.00257353
R8129 vss.n593 vss.n592 0.00257353
R8130 vss.n602 vss.n601 0.00257353
R8131 vss.n604 vss.n603 0.00257353
R8132 vss.n613 vss.n612 0.00257353
R8133 vss.n615 vss.n614 0.00257353
R8134 vss.n1231 vss.n1230 0.00257353
R8135 vss.n1229 vss.n1228 0.00257353
R8136 vss.n1211 vss.n1210 0.00257353
R8137 vss.n1209 vss.n1208 0.00257353
R8138 vss.n1200 vss.n1199 0.00257353
R8139 vss.n1198 vss.n1197 0.00257353
R8140 vss.n1182 vss.n1181 0.00257353
R8141 vss.n1180 vss.n1179 0.00257353
R8142 vss.n1167 vss.n1166 0.00257353
R8143 vss.n1165 vss.n1164 0.00257353
R8144 vss.n1159 vss.n1158 0.00257353
R8145 vss.n1157 vss.n1156 0.00257353
R8146 vss.n1148 vss.n1147 0.00257353
R8147 vss.n1146 vss.n1145 0.00257353
R8148 vss.n1137 vss.n1136 0.00257353
R8149 vss.n1135 vss.n1134 0.00257353
R8150 vss.n956 vss.n616 0.00257353
R8151 vss.n958 vss.n957 0.00257353
R8152 vss.n992 vss.n991 0.00257353
R8153 vss.n994 vss.n993 0.00257353
R8154 vss.n997 vss.n996 0.00257353
R8155 vss.n999 vss.n998 0.00257353
R8156 vss.n1002 vss.n1001 0.00257353
R8157 vss.n1004 vss.n1003 0.00257353
R8158 vss.n1021 vss.n1020 0.00257353
R8159 vss.n1023 vss.n1022 0.00257353
R8160 vss.n1026 vss.n1025 0.00257353
R8161 vss.n1028 vss.n1027 0.00257353
R8162 vss.n1031 vss.n1030 0.00257353
R8163 vss.n1033 vss.n1032 0.00257353
R8164 vss.n912 vss.n911 0.00257353
R8165 vss.n914 vss.n913 0.00257353
R8166 vss.n917 vss.n916 0.00257353
R8167 vss.n919 vss.n918 0.00257353
R8168 vss.n922 vss.n921 0.00257353
R8169 vss.n924 vss.n923 0.00257353
R8170 vss.n1569 vss.n1568 0.00233824
R8171 vss.n1565 vss.n1561 0.00233824
R8172 vss.n1558 vss.n1555 0.00233824
R8173 vss.n542 vss.n541 0.00233824
R8174 vss.n548 vss.n547 0.00233824
R8175 vss.n554 vss.n553 0.00233824
R8176 vss.n1491 vss.n1490 0.00233824
R8177 vss.n1497 vss.n1496 0.00233824
R8178 vss.n1504 vss.n1503 0.00233824
R8179 vss.n1514 vss.n1513 0.00233824
R8180 vss.n1520 vss.n1519 0.00233824
R8181 vss.n1544 vss.n1525 0.00233824
R8182 vss.n1281 vss.n1280 0.00233824
R8183 vss.n1287 vss.n1286 0.00233824
R8184 vss.n1294 vss.n1293 0.00233824
R8185 vss.n1257 vss.n1255 0.00233824
R8186 vss.n1268 vss.n1266 0.00233824
R8187 vss.n1301 vss.n1277 0.00233824
R8188 vss.n1319 vss.n1316 0.00233824
R8189 vss.n1325 vss.n1322 0.00233824
R8190 vss.n1341 vss.n1340 0.00233824
R8191 vss.n1308 vss.n1242 0.00233824
R8192 vss.n1237 vss.n1236 0.00233824
R8193 vss.n1333 vss.n1332 0.00233824
R8194 vss.n1484 vss.n1483 0.00233824
R8195 vss.n1480 vss.n1476 0.00233824
R8196 vss.n1473 vss.n1470 0.00233824
R8197 vss.n443 vss.n441 0.00233824
R8198 vss.n454 vss.n452 0.00233824
R8199 vss.n1462 vss.n428 0.00233824
R8200 vss.n1366 vss.n1362 0.00233824
R8201 vss.n1373 vss.n1369 0.00233824
R8202 vss.n1405 vss.n1404 0.00233824
R8203 vss.n1355 vss.n1350 0.00233824
R8204 vss.n1345 vss.n1344 0.00233824
R8205 vss.n1381 vss.n1380 0.00233824
R8206 vss.n688 vss.n687 0.00233824
R8207 vss.n695 vss.n694 0.00233824
R8208 vss.n701 vss.n700 0.00233824
R8209 vss.n664 vss.n662 0.00233824
R8210 vss.n675 vss.n673 0.00233824
R8211 vss.n708 vss.n684 0.00233824
R8212 vss.n719 vss.n718 0.00233824
R8213 vss.n753 vss.n752 0.00233824
R8214 vss.n791 vss.n790 0.00233824
R8215 vss.n728 vss.n727 0.00233824
R8216 vss.n739 vss.n738 0.00233824
R8217 vss.n756 vss.n755 0.00233824
R8218 vss.n837 vss.n836 0.00233824
R8219 vss.n844 vss.n843 0.00233824
R8220 vss.n850 vss.n849 0.00233824
R8221 vss.n812 vss.n810 0.00233824
R8222 vss.n823 vss.n821 0.00233824
R8223 vss.n858 vss.n832 0.00233824
R8224 vss.n876 vss.n872 0.00233824
R8225 vss.n883 vss.n879 0.00233824
R8226 vss.n1016 vss.n1015 0.00233824
R8227 vss.n865 vss.n649 0.00233824
R8228 vss.n644 vss.n643 0.00233824
R8229 vss.n638 vss.n637 0.00233824
R8230 vss.n1413 vss.n1412 0.00233824
R8231 vss.n1419 vss.n1418 0.00233824
R8232 vss.n1426 vss.n1425 0.00233824
R8233 vss.n599 vss.n597 0.00233824
R8234 vss.n610 vss.n608 0.00233824
R8235 vss.n1434 vss.n1235 0.00233824
R8236 vss.n1216 vss.n1215 0.00233824
R8237 vss.n1192 vss.n1191 0.00233824
R8238 vss.n1175 vss.n1174 0.00233824
R8239 vss.n1226 vss.n1225 0.00233824
R8240 vss.n1206 vss.n1205 0.00233824
R8241 vss.n1195 vss.n1194 0.00233824
R8242 vss.n1112 vss.n1111 0.00233824
R8243 vss.n1118 vss.n1117 0.00233824
R8244 vss.n1125 vss.n1124 0.00233824
R8245 vss.n1154 vss.n1152 0.00233824
R8246 vss.n1143 vss.n1141 0.00233824
R8247 vss.n1132 vss.n1108 0.00233824
R8248 vss.n971 vss.n968 0.00233824
R8249 vss.n977 vss.n974 0.00233824
R8250 vss.n1009 vss.n1008 0.00233824
R8251 vss.n960 vss.n955 0.00233824
R8252 vss.n950 vss.n949 0.00233824
R8253 vss.n985 vss.n984 0.00233824
R8254 vss.n1064 vss.n1061 0.00233824
R8255 vss.n1070 vss.n1067 0.00233824
R8256 vss.n1076 vss.n1075 0.00233824
R8257 vss.n1054 vss.n1051 0.00233824
R8258 vss.n1046 vss.n1045 0.00233824
R8259 vss.n1040 vss.n1039 0.00233824
R8260 vss.n942 vss.n941 0.00233824
R8261 vss.n935 vss.n934 0.00233824
R8262 vss.n928 vss.n899 0.00233824
R8263 vss.n895 vss.n892 0.00233824
R8264 vss.n887 vss.n886 0.00233824
R8265 vss.n905 vss.n904 0.00233824
R8266 vss.n1088 vss.n1087 0.00230077
R8267 vss.n1085 vss.n1084 0.00230077
R8268 vss.n1082 vss.n1081 0.00230077
R8269 vss.n1444 vss.n1443 0.00230077
R8270 vss.n1441 vss.n1440 0.00230077
R8271 vss.n1438 vss.n1437 0.00230077
R8272 vss.n765 vss.n764 0.00230077
R8273 vss.n768 vss.n767 0.00230077
R8274 vss.n771 vss.n770 0.00230077
R8275 vss.n778 vss.n777 0.00230077
R8276 vss.n775 vss.n774 0.00230077
R8277 vss.n772 vss.n617 0.00230077
R8278 vss.n1100 vss.n1099 0.00230077
R8279 vss.n1097 vss.n1096 0.00230077
R8280 vss.n1094 vss.n1093 0.00230077
R8281 vss.n561 vss.n560 0.00230077
R8282 vss.n564 vss.n563 0.00230077
R8283 vss.n567 vss.n566 0.00230077
R8284 vss.n1456 vss.n1455 0.00230077
R8285 vss.n1453 vss.n1452 0.00230077
R8286 vss.n1450 vss.n1449 0.00230077
R8287 vss.n511 vss.n510 0.00230077
R8288 vss.n514 vss.n513 0.00230077
R8289 vss.n517 vss.n516 0.00230077
R8290 vss.n29 vss.n25 0.00218919
R8291 vss.n193 vss.n174 0.00218919
R8292 vss.n208 vss.n200 0.00218919
R8293 vss.n52 vss.n22 0.00218919
R8294 vss.n503 vss.n501 0.0021514
R8295 vss.n474 vss.n472 0.0021514
R8296 vss.n90 vss.n85 0.0020528
R8297 vss.n171 vss.n170 0.00198734
R8298 vss.n170 vss.n0 0.00198734
R8299 vss.n1640 vss.n1639 0.00198734
R8300 vss.n1639 vss.n2 0.00198734
R8301 vss.n198 vss.n197 0.00196875
R8302 vss.n196 vss.n195 0.00196875
R8303 vss.n159 vss.n158 0.00196875
R8304 vss.n161 vss.n160 0.00196875
R8305 vss.n27 vss.n17 0.00196875
R8306 vss.n55 vss.n54 0.00196875
R8307 vss.n20 vss.n19 0.00196875
R8308 vss.n18 vss.n15 0.00196875
R8309 vss.n339 vss.n321 0.0018975
R8310 vss.n207 vss.n206 0.00180208
R8311 vss.n191 vss.n185 0.00180208
R8312 vss.n24 vss.n23 0.00180208
R8313 vss.n50 vss.n46 0.00180208
R8314 vss.n483 vss 0.00170192
R8315 vss.n321 vss.n320 0.00130908
R8316 vss.n313 vss.n310 0.00121429
R8317 vss.n465 vss.n464 0.0011215
R8318 vss.n494 vss.n493 0.0011215
R8319 vss vss.n0 0.00109494
R8320 vss.n172 vss.n171 0.000797468
R8321 vss.n56 vss.n2 0.000797468
R8322 async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[1].t0 140.387
R8323 async_resetb_delay_ctrl_code[1].n0 async_resetb_delay_ctrl_code[1].t1 140.34
R8324 async_resetb_delay_ctrl_code[1].n0 async_resetb_delay_ctrl_code[1] 0.204648
R8325 async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[1].n0 0.00217851
R8326 eob eob.n9 352.005
R8327 eob.n6 eob.t3 329.01
R8328 eob.n9 eob.t2 272.062
R8329 eob.n9 eob.t1 206.19
R8330 eob.n5 eob.t0 140.888
R8331 eob.n10 eob 26.2742
R8332 eob.n7 eob.n6 9.3005
R8333 eob.n6 eob.n5 7.71392
R8334 eob.n1 eob 4.94565
R8335 eob eob.n10 4.71629
R8336 eob.n7 eob.n4 2.84654
R8337 eob.n3 eob.n1 1.12162
R8338 eob eob.n8 0.674184
R8339 eob.n8 eob.n7 0.337342
R8340 eob.n1 eob.n0 0.00956032
R8341 eob.n4 eob.n3 0.00699236
R8342 eob.n3 eob.n2 0.00269298
R8343 sample_clk sample_clk.n6 352.005
R8344 sample_clk.n3 sample_clk.t5 329.767
R8345 sample_clk.n6 sample_clk.t4 272.062
R8346 sample_clk.n11 sample_clk.t1 269.921
R8347 sample_clk.n11 sample_clk.t2 234.573
R8348 sample_clk.n6 sample_clk.t3 206.19
R8349 sample_clk.n3 sample_clk.t0 147.18
R8350 sample_clk.n12 sample_clk.n11 76.0005
R8351 sample_clk.n7 sample_clk 25.6005
R8352 sample_clk sample_clk.n10 12.5496
R8353 sample_clk.n5 sample_clk.n4 9.30195
R8354 sample_clk.n8 sample_clk.n7 9.3005
R8355 sample_clk sample_clk.n12 7.57233
R8356 sample_clk.n5 sample_clk.n3 7.16864
R8357 sample_clk.n7 sample_clk 5.38997
R8358 sample_clk.n12 sample_clk 4.68782
R8359 sample_clk sample_clk.n2 3.03311
R8360 sample_clk.n10 sample_clk.n9 2.24192
R8361 sample_clk.n0 sample_clk 1.66492
R8362 sample_clk sample_clk.n5 0.337342
R8363 sample_clk.n1 sample_clk.n0 0.0369583
R8364 sample_clk.n9 sample_clk.n8 0.0213333
R8365 sample_clk.n10 sample_clk.n1 0.0208917
R8366 sample_clk.n9 sample_clk.n2 0.0099697
R8367 sample_clk.n4 sample_clk.n2 0.0019432
R8368 ready.t10 ready.t19 221.72
R8369 ready.t3 ready.t10 221.72
R8370 ready.t16 ready.t3 221.72
R8371 ready.t4 ready.t16 221.72
R8372 ready.t21 ready.t4 221.72
R8373 ready.t12 ready.t21 221.72
R8374 ready.t8 ready.t12 221.72
R8375 ready.t14 ready.t1 221.72
R8376 ready.t5 ready.t14 221.72
R8377 ready.t17 ready.t5 221.72
R8378 ready.t7 ready.t17 221.72
R8379 ready.t0 ready.t7 221.72
R8380 ready.t15 ready.t0 221.72
R8381 ready.t9 ready.t15 221.72
R8382 ready.t20 ready.t11 221.72
R8383 ready.t2 ready.t20 221.72
R8384 ready.t13 ready.t2 221.72
R8385 ready.t18 ready.t13 221.72
R8386 ready.t6 ready.t18 221.72
R8387 ready.n4 ready.t6 154.8
R8388 ready.n2 ready.t9 98.5385
R8389 ready.n0 ready 89.9738
R8390 ready.n0 ready.t8 74.8959
R8391 ready.n1 ready 40.1672
R8392 ready.n3 ready.n0 21.3003
R8393 ready.n3 ready.n2 19.0526
R8394 ready.n5 ready.n3 13.9039
R8395 ready.n1 ready 11.8854
R8396 ready.n2 ready.n1 2.56597
R8397 ready ready.n5 1.64944
R8398 ready ready.n4 1.10206
R8399 ready.n4 ready 0.10169
R8400 ready.n5 ready 0.0603958
R8401 ready.n4 ready 0.0447708
R8402 async_clk_sar async_clk_sar.n0 294.219
R8403 async_clk_sar.n2 async_clk_sar.n0 292.5
R8404 async_clk_sar.n1 async_clk_sar.n0 292.5
R8405 async_clk_sar.t2 async_clk_sar.t18 221.72
R8406 async_clk_sar.t16 async_clk_sar.t2 221.72
R8407 async_clk_sar.t21 async_clk_sar.t16 221.72
R8408 async_clk_sar.t7 async_clk_sar.t21 221.72
R8409 async_clk_sar.t12 async_clk_sar.t7 221.72
R8410 async_clk_sar.t13 async_clk_sar.t8 221.72
R8411 async_clk_sar.t5 async_clk_sar.t13 221.72
R8412 async_clk_sar.t17 async_clk_sar.t5 221.72
R8413 async_clk_sar.t11 async_clk_sar.t17 221.72
R8414 async_clk_sar.t23 async_clk_sar.t11 221.72
R8415 async_clk_sar.t19 async_clk_sar.t23 221.72
R8416 async_clk_sar.t6 async_clk_sar.t19 221.72
R8417 async_clk_sar.t9 async_clk_sar.t3 221.72
R8418 async_clk_sar.t14 async_clk_sar.t9 221.72
R8419 async_clk_sar.t20 async_clk_sar.t14 221.72
R8420 async_clk_sar.t15 async_clk_sar.t20 221.72
R8421 async_clk_sar.t4 async_clk_sar.t15 221.72
R8422 async_clk_sar.t22 async_clk_sar.t4 221.72
R8423 async_clk_sar.t10 async_clk_sar.t22 221.72
R8424 async_clk_sar.n12 async_clk_sar.t12 153.184
R8425 async_clk_sar.n4 async_clk_sar 89.9738
R8426 async_clk_sar.n5 async_clk_sar.t6 78.7272
R8427 async_clk_sar.n4 async_clk_sar.t10 74.6592
R8428 async_clk_sar async_clk_sar.n2 68.2971
R8429 async_clk_sar.n6 async_clk_sar 40.1672
R8430 async_clk_sar.n3 async_clk_sar.t0 36.1131
R8431 async_clk_sar.n7 async_clk_sar.n5 32.1338
R8432 async_clk_sar.n14 async_clk_sar.n3 29.2039
R8433 async_clk_sar.n0 async_clk_sar.t1 26.5955
R8434 async_clk_sar async_clk_sar.n5 21.4227
R8435 async_clk_sar.n8 async_clk_sar.n4 21.3547
R8436 async_clk_sar.n8 async_clk_sar.n7 17.8279
R8437 async_clk_sar.n10 async_clk_sar.n8 13.4143
R8438 async_clk_sar.n6 async_clk_sar 11.8854
R8439 async_clk_sar.n2 async_clk_sar 11.2721
R8440 async_clk_sar.n1 async_clk_sar 11.2721
R8441 async_clk_sar.n13 async_clk_sar.n11 4.5663
R8442 async_clk_sar.n7 async_clk_sar.n6 3.96214
R8443 async_clk_sar async_clk_sar.n13 3.66629
R8444 async_clk_sar.n3 async_clk_sar 3.32947
R8445 async_clk_sar async_clk_sar.n1 1.7199
R8446 async_clk_sar.n9 async_clk_sar 1.64944
R8447 async_clk_sar.n13 async_clk_sar.n12 1.11962
R8448 async_clk_sar.n9 async_clk_sar 0.124699
R8449 async_clk_sar.n12 async_clk_sar 0.10169
R8450 async_clk_sar.n12 async_clk_sar 0.0391364
R8451 async_clk_sar.n11 async_clk_sar.n10 0.0265016
R8452 async_clk_sar async_clk_sar.n14 0.0225588
R8453 async_clk_sar.n14 async_clk_sar 0.0149231
R8454 async_clk_sar async_clk_sar.n11 0.0118636
R8455 async_clk_sar.n10 async_clk_sar.n9 0.00430609
R8456 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[2].t1 140.387
R8457 async_resetb_delay_ctrl_code[2].n2 async_resetb_delay_ctrl_code[2].t2 140.34
R8458 async_resetb_delay_ctrl_code[2].n1 async_resetb_delay_ctrl_code[2].t3 140.34
R8459 async_resetb_delay_ctrl_code[2].n0 async_resetb_delay_ctrl_code[2].t0 140.34
R8460 async_resetb_delay_ctrl_code[2].n2 async_resetb_delay_ctrl_code[2] 2.83
R8461 async_resetb_delay_ctrl_code[2].n1 async_resetb_delay_ctrl_code[2] 0.285826
R8462 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[2].n0 0.264087
R8463 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[2].n1 0.0466957
R8464 async_resetb_delay_ctrl_code[2].n0 async_resetb_delay_ctrl_code[2] 0.0466957
R8465 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[2].n2 0.0022562
R8466 delay_offset.n11 delay_offset.t0 230.016
R8467 delay_offset.n1 delay_offset.t5 229.964
R8468 delay_offset.n1 delay_offset.t3 158.363
R8469 delay_offset.n10 delay_offset.t2 153.665
R8470 delay_offset.n11 delay_offset 153.601
R8471 delay_offset delay_offset.t4 140.379
R8472 delay_offset delay_offset.t1 140.379
R8473 delay_offset.n10 delay_offset.n9 73.8234
R8474 delay_offset.n12 delay_offset.n11 9.3005
R8475 delay_offset.n2 delay_offset.n1 7.39235
R8476 delay_offset delay_offset.n16 5.89437
R8477 delay_offset.n11 delay_offset.n10 4.91671
R8478 delay_offset.n14 delay_offset.n12 4.9013
R8479 delay_offset.n16 delay_offset 4.80627
R8480 delay_offset.n13 delay_offset 4.22092
R8481 delay_offset.n7 delay_offset 4.22092
R8482 delay_offset.n3 delay_offset 2.48404
R8483 delay_offset.n4 delay_offset.n3 2.47689
R8484 delay_offset delay_offset.n9 2.4005
R8485 delay_offset.n8 delay_offset.n6 1.87694
R8486 delay_offset.n6 delay_offset.n5 1.12626
R8487 delay_offset.n3 delay_offset.n2 1.02104
R8488 delay_offset.n13 delay_offset 1.01229
R8489 delay_offset.n7 delay_offset 1.01229
R8490 delay_offset.n14 delay_offset.n13 0.726043
R8491 delay_offset.n8 delay_offset.n7 0.726043
R8492 delay_offset.n12 delay_offset.n9 0.533833
R8493 delay_offset.n15 delay_offset.n14 0.421696
R8494 delay_offset.n17 delay_offset.n8 0.421696
R8495 delay_offset.n17 delay_offset 0.203802
R8496 delay_offset delay_offset.n15 0.0447308
R8497 delay_offset delay_offset.n17 0.0447308
R8498 delay_offset.n15 delay_offset 0.0195217
R8499 delay_offset.n17 delay_offset 0.0195217
R8500 delay_offset.n4 delay_offset.n0 0.0179598
R8501 delay_offset.n16 delay_offset 0.00626923
R8502 delay_offset.n5 delay_offset.n4 0.00504545
R8503 async_resetb_delay_ctrl_code[3].n0 async_resetb_delay_ctrl_code[3].t1 229.971
R8504 async_resetb_delay_ctrl_code[3].n0 async_resetb_delay_ctrl_code[3].t0 158.35
R8505 async_resetb_delay_ctrl_code[3].n1 async_resetb_delay_ctrl_code[3].n0 8.50845
R8506 async_resetb_delay_ctrl_code[3].n1 async_resetb_delay_ctrl_code[3] 3.95275
R8507 async_resetb_delay_ctrl_code[3].n2 async_resetb_delay_ctrl_code[3].n1 1.73287
R8508 async_resetb_delay_ctrl_code[3].n3 async_resetb_delay_ctrl_code[3] 0.474765
R8509 async_resetb_delay_ctrl_code[3] async_resetb_delay_ctrl_code[3].n3 0.366977
R8510 async_resetb_delay_ctrl_code[3].n2 async_resetb_delay_ctrl_code[3] 0.339042
R8511 async_resetb_delay_ctrl_code[3].n3 async_resetb_delay_ctrl_code[3].n2 0.00334091
R8512 async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[0].t0 140.343
R8513 x2.x10.Y x2.x10.Y.t9 154.847
R8514 x2.x10.Y x2.x10.Y.t2 154.8
R8515 x2.x10.Y x2.x10.Y.t8 154.8
R8516 x2.x10.Y x2.x10.Y.t3 154.8
R8517 x2.x10.Y x2.x10.Y.t6 154.8
R8518 x2.x10.Y x2.x10.Y.t4 154.8
R8519 x2.x10.Y x2.x10.Y.t7 154.8
R8520 x2.x10.Y x2.x10.Y.t5 154.8
R8521 x2.x10.Y.n1 x2.x10.Y 134.254
R8522 x2.x10.Y x2.x10.Y.t1 116.097
R8523 x2.x10.Y.n3 x2.x10.Y.t0 24.6255
R8524 x2.x10.Y.n0 x2.x10.Y 11.6875
R8525 x2.x10.Y.n4 x2.x10.Y.n3 9.3005
R8526 x2.x10.Y x2.x10.Y.n5 8.87659
R8527 x2.x10.Y.n0 x2.x10.Y 7.23528
R8528 x2.x10.Y.n5 x2.x10.Y.n4 5.94566
R8529 x2.x10.Y x2.x10.Y.n0 5.04292
R8530 x2.x10.Y.n3 x2.x10.Y.n2 1.9705
R8531 x2.x10.Y.n4 x2.x10.Y.n1 0.652832
R8532 x2.x5[7].floating.n143 x2.x5[7].floating.t1 68.0345
R8533 x2.x5[7].floating.n155 x2.x5[7].floating.t7 68.0345
R8534 x2.x5[7].floating.n48 x2.x5[7].floating.t0 68.0345
R8535 x2.x5[7].floating.n60 x2.x5[7].floating.t4 68.0345
R8536 x2.x5[7].floating.n78 x2.x5[7].floating.t2 68.0345
R8537 x2.x5[7].floating.n90 x2.x5[7].floating.t5 68.0345
R8538 x2.x5[7].floating.n108 x2.x5[7].floating.t3 68.0345
R8539 x2.x5[7].floating.n122 x2.x5[7].floating.t6 68.0345
R8540 x2.x5[7].floating.n139 x2.x5[7].floating.n5 0.660401
R8541 x2.x5[7].floating.n100 x2.x5[7].floating.n14 0.660401
R8542 x2.x5[7].floating.n85 x2.x5[7].floating.n23 0.660401
R8543 x2.x5[7].floating.n70 x2.x5[7].floating.n32 0.660401
R8544 x2.x5[7].floating.n130 x2.x5[7].floating.n129 0.660401
R8545 x2.x5[7].floating.n46 x2.x5[7].floating.n45 0.320345
R8546 x2.x5[7].floating.n160 x2.x5[7].floating.n159 0.308269
R8547 x2.x5[7].floating.n161 x2.x5[7].floating.n160 0.173084
R8548 x2.x5[7].floating.n45 x2.x5[7].floating.n44 0.162103
R8549 x2.x5[7].floating.n160 x2.x5[7].floating 0.100688
R8550 x2.x5[7].floating.n45 x2.x5[7].floating 0.0755007
R8551 x2.x5[7].floating.n115 x2.x5[7].floating.n5 0.0716912
R8552 x2.x5[7].floating.n5 x2.x5[7].floating.n4 0.0716912
R8553 x2.x5[7].floating.n100 x2.x5[7].floating.n99 0.0716912
R8554 x2.x5[7].floating.n101 x2.x5[7].floating.n100 0.0716912
R8555 x2.x5[7].floating.n70 x2.x5[7].floating.n69 0.0716912
R8556 x2.x5[7].floating.n71 x2.x5[7].floating.n70 0.0716912
R8557 x2.x5[7].floating.n32 x2.x5[7].floating.n31 0.0716912
R8558 x2.x5[7].floating.n14 x2.x5[7].floating.n13 0.0716912
R8559 x2.x5[7].floating.n140 x2.x5[7].floating.n139 0.0716912
R8560 x2.x5[7].floating.n119 x2.x5[7].floating.n118 0.0557941
R8561 x2.x5[7].floating.n118 x2.x5[7].floating.n117 0.0557941
R8562 x2.x5[7].floating.n117 x2.x5[7].floating.n116 0.0557941
R8563 x2.x5[7].floating.n116 x2.x5[7].floating.n115 0.0557941
R8564 x2.x5[7].floating.n4 x2.x5[7].floating.n3 0.0557941
R8565 x2.x5[7].floating.n3 x2.x5[7].floating.n2 0.0557941
R8566 x2.x5[7].floating.n2 x2.x5[7].floating.n1 0.0557941
R8567 x2.x5[7].floating.n1 x2.x5[7].floating.n0 0.0557941
R8568 x2.x5[7].floating.n96 x2.x5[7].floating.n95 0.0557941
R8569 x2.x5[7].floating.n97 x2.x5[7].floating.n96 0.0557941
R8570 x2.x5[7].floating.n98 x2.x5[7].floating.n97 0.0557941
R8571 x2.x5[7].floating.n99 x2.x5[7].floating.n98 0.0557941
R8572 x2.x5[7].floating.n102 x2.x5[7].floating.n101 0.0557941
R8573 x2.x5[7].floating.n103 x2.x5[7].floating.n102 0.0557941
R8574 x2.x5[7].floating.n104 x2.x5[7].floating.n103 0.0557941
R8575 x2.x5[7].floating.n105 x2.x5[7].floating.n104 0.0557941
R8576 x2.x5[7].floating.n66 x2.x5[7].floating.n65 0.0557941
R8577 x2.x5[7].floating.n67 x2.x5[7].floating.n66 0.0557941
R8578 x2.x5[7].floating.n68 x2.x5[7].floating.n67 0.0557941
R8579 x2.x5[7].floating.n69 x2.x5[7].floating.n68 0.0557941
R8580 x2.x5[7].floating.n72 x2.x5[7].floating.n71 0.0557941
R8581 x2.x5[7].floating.n73 x2.x5[7].floating.n72 0.0557941
R8582 x2.x5[7].floating.n74 x2.x5[7].floating.n73 0.0557941
R8583 x2.x5[7].floating.n75 x2.x5[7].floating.n74 0.0557941
R8584 x2.x5[7].floating.n37 x2.x5[7].floating.n36 0.0557941
R8585 x2.x5[7].floating.n36 x2.x5[7].floating.n35 0.0557941
R8586 x2.x5[7].floating.n35 x2.x5[7].floating.n34 0.0557941
R8587 x2.x5[7].floating.n34 x2.x5[7].floating.n33 0.0557941
R8588 x2.x5[7].floating.n30 x2.x5[7].floating.n29 0.0557941
R8589 x2.x5[7].floating.n29 x2.x5[7].floating.n28 0.0557941
R8590 x2.x5[7].floating.n28 x2.x5[7].floating.n27 0.0557941
R8591 x2.x5[7].floating.n19 x2.x5[7].floating.n18 0.0557941
R8592 x2.x5[7].floating.n18 x2.x5[7].floating.n17 0.0557941
R8593 x2.x5[7].floating.n17 x2.x5[7].floating.n16 0.0557941
R8594 x2.x5[7].floating.n16 x2.x5[7].floating.n15 0.0557941
R8595 x2.x5[7].floating.n12 x2.x5[7].floating.n11 0.0557941
R8596 x2.x5[7].floating.n11 x2.x5[7].floating.n10 0.0557941
R8597 x2.x5[7].floating.n10 x2.x5[7].floating.n9 0.0557941
R8598 x2.x5[7].floating.n135 x2.x5[7].floating.n134 0.0557941
R8599 x2.x5[7].floating.n136 x2.x5[7].floating.n135 0.0557941
R8600 x2.x5[7].floating.n137 x2.x5[7].floating.n136 0.0557941
R8601 x2.x5[7].floating.n138 x2.x5[7].floating.n137 0.0557941
R8602 x2.x5[7].floating.n171 x2.x5[7].floating.n170 0.0557941
R8603 x2.x5[7].floating.n170 x2.x5[7].floating.n169 0.0557941
R8604 x2.x5[7].floating.n169 x2.x5[7].floating.n168 0.0557941
R8605 x2.x5[7].floating.n41 x2.x5[7].floating.n40 0.0537206
R8606 x2.x5[7].floating.n23 x2.x5[7].floating.n22 0.0537206
R8607 x2.x5[7].floating.n131 x2.x5[7].floating.n130 0.0537206
R8608 x2.x5[7].floating.n164 x2.x5[7].floating.n163 0.0537206
R8609 x2.x5[7].floating.n42 x2.x5[7].floating.n41 0.0530294
R8610 x2.x5[7].floating.n24 x2.x5[7].floating.n23 0.0530294
R8611 x2.x5[7].floating.n130 x2.x5[7].floating.n6 0.0530294
R8612 x2.x5[7].floating.n165 x2.x5[7].floating.n164 0.0530294
R8613 x2.x5[7].floating.n151 x2.x5[7].floating.n150 0.0529559
R8614 x2.x5[7].floating.n86 x2.x5[7].floating.n85 0.0529559
R8615 x2.x5[7].floating.n56 x2.x5[7].floating.n55 0.0529559
R8616 x2.x5[7].floating.n129 x2.x5[7].floating.n128 0.0529559
R8617 x2.x5[7].floating.n150 x2.x5[7].floating.n149 0.0524559
R8618 x2.x5[7].floating.n129 x2.x5[7].floating.n114 0.0524559
R8619 x2.x5[7].floating.n85 x2.x5[7].floating.n84 0.0524559
R8620 x2.x5[7].floating.n55 x2.x5[7].floating.n54 0.0524559
R8621 x2.x5[7].floating.n27 x2.x5[7].floating.n26 0.0523382
R8622 x2.x5[7].floating.n9 x2.x5[7].floating.n8 0.0523382
R8623 x2.x5[7].floating.n168 x2.x5[7].floating.n167 0.0523382
R8624 x2.x5[7].floating.n38 x2.x5[7].floating.n37 0.0516471
R8625 x2.x5[7].floating.n20 x2.x5[7].floating.n19 0.0516471
R8626 x2.x5[7].floating.n134 x2.x5[7].floating.n133 0.0516471
R8627 x2.x5[7].floating x2.x5[7].floating.n32 0.0495735
R8628 x2.x5[7].floating x2.x5[7].floating.n14 0.0495735
R8629 x2.x5[7].floating.n139 x2.x5[7].floating 0.0495735
R8630 x2.x5[7].floating.n145 x2.x5[7].floating.n142 0.0408846
R8631 x2.x5[7].floating.n50 x2.x5[7].floating.n47 0.0408846
R8632 x2.x5[7].floating.n80 x2.x5[7].floating.n77 0.0408846
R8633 x2.x5[7].floating.n110 x2.x5[7].floating.n107 0.0408846
R8634 x2.x5[7].floating x2.x5[7].floating.n30 0.0336765
R8635 x2.x5[7].floating x2.x5[7].floating.n12 0.0336765
R8636 x2.x5[7].floating x2.x5[7].floating.n171 0.0336765
R8637 x2.x5[7].floating.n106 x2.x5[7].floating.n105 0.0271618
R8638 x2.x5[7].floating.n76 x2.x5[7].floating.n75 0.0271618
R8639 x2.x5[7].floating.n120 x2.x5[7].floating.n119 0.0266618
R8640 x2.x5[7].floating.n95 x2.x5[7].floating.n94 0.0266618
R8641 x2.x5[7].floating.n65 x2.x5[7].floating.n64 0.0266618
R8642 x2.x5[7].floating.n33 x2.x5[7].floating 0.0226176
R8643 x2.x5[7].floating.n31 x2.x5[7].floating 0.0226176
R8644 x2.x5[7].floating.n15 x2.x5[7].floating 0.0226176
R8645 x2.x5[7].floating.n13 x2.x5[7].floating 0.0226176
R8646 x2.x5[7].floating x2.x5[7].floating.n138 0.0226176
R8647 x2.x5[7].floating x2.x5[7].floating.n140 0.0226176
R8648 x2.x5[7].floating.n43 x2.x5[7].floating.n42 0.0191618
R8649 x2.x5[7].floating.n25 x2.x5[7].floating.n24 0.0191618
R8650 x2.x5[7].floating.n7 x2.x5[7].floating.n6 0.0191618
R8651 x2.x5[7].floating.n166 x2.x5[7].floating.n165 0.0191618
R8652 x2.x5[7].floating.n40 x2.x5[7].floating.n39 0.0184706
R8653 x2.x5[7].floating.n22 x2.x5[7].floating.n21 0.0184706
R8654 x2.x5[7].floating.n132 x2.x5[7].floating.n131 0.0184706
R8655 x2.x5[7].floating.n163 x2.x5[7].floating.n162 0.0184706
R8656 x2.x5[7].floating.n159 x2.x5[7].floating.n158 0.014
R8657 x2.x5[7].floating.n149 x2.x5[7].floating.n148 0.014
R8658 x2.x5[7].floating.n114 x2.x5[7].floating.n113 0.014
R8659 x2.x5[7].floating.n94 x2.x5[7].floating.n93 0.014
R8660 x2.x5[7].floating.n84 x2.x5[7].floating.n83 0.014
R8661 x2.x5[7].floating.n64 x2.x5[7].floating.n63 0.014
R8662 x2.x5[7].floating.n54 x2.x5[7].floating.n53 0.014
R8663 x2.x5[7].floating.n125 x2.x5[7].floating.n120 0.014
R8664 x2.x5[7].floating.n152 x2.x5[7].floating.n151 0.0135
R8665 x2.x5[7].floating.n146 x2.x5[7].floating.n141 0.0135
R8666 x2.x5[7].floating.n111 x2.x5[7].floating.n106 0.0135
R8667 x2.x5[7].floating.n87 x2.x5[7].floating.n86 0.0135
R8668 x2.x5[7].floating.n81 x2.x5[7].floating.n76 0.0135
R8669 x2.x5[7].floating.n57 x2.x5[7].floating.n56 0.0135
R8670 x2.x5[7].floating.n51 x2.x5[7].floating.n46 0.0135
R8671 x2.x5[7].floating.n128 x2.x5[7].floating.n127 0.0135
R8672 x2.x5[7].floating.n157 x2.x5[7].floating.n154 0.0101154
R8673 x2.x5[7].floating.n62 x2.x5[7].floating.n59 0.0101154
R8674 x2.x5[7].floating.n92 x2.x5[7].floating.n89 0.0101154
R8675 x2.x5[7].floating.n124 x2.x5[7].floating.n121 0.0101154
R8676 x2.x5[7].floating.n39 x2.x5[7].floating.n38 0.00464706
R8677 x2.x5[7].floating.n21 x2.x5[7].floating.n20 0.00464706
R8678 x2.x5[7].floating.n133 x2.x5[7].floating.n132 0.00464706
R8679 x2.x5[7].floating.n162 x2.x5[7].floating.n161 0.00464706
R8680 x2.x5[7].floating.n44 x2.x5[7].floating.n43 0.00395588
R8681 x2.x5[7].floating.n26 x2.x5[7].floating.n25 0.00395588
R8682 x2.x5[7].floating.n8 x2.x5[7].floating.n7 0.00395588
R8683 x2.x5[7].floating.n167 x2.x5[7].floating.n166 0.00395588
R8684 x2.x5[7].floating.n153 x2.x5[7].floating.n152 0.0035
R8685 x2.x5[7].floating.n147 x2.x5[7].floating.n146 0.0035
R8686 x2.x5[7].floating.n112 x2.x5[7].floating.n111 0.0035
R8687 x2.x5[7].floating.n88 x2.x5[7].floating.n87 0.0035
R8688 x2.x5[7].floating.n82 x2.x5[7].floating.n81 0.0035
R8689 x2.x5[7].floating.n58 x2.x5[7].floating.n57 0.0035
R8690 x2.x5[7].floating.n52 x2.x5[7].floating.n51 0.0035
R8691 x2.x5[7].floating.n127 x2.x5[7].floating.n126 0.0035
R8692 x2.x5[7].floating.n158 x2.x5[7].floating.n153 0.003
R8693 x2.x5[7].floating.n148 x2.x5[7].floating.n147 0.003
R8694 x2.x5[7].floating.n113 x2.x5[7].floating.n112 0.003
R8695 x2.x5[7].floating.n93 x2.x5[7].floating.n88 0.003
R8696 x2.x5[7].floating.n83 x2.x5[7].floating.n82 0.003
R8697 x2.x5[7].floating.n63 x2.x5[7].floating.n58 0.003
R8698 x2.x5[7].floating.n53 x2.x5[7].floating.n52 0.003
R8699 x2.x5[7].floating.n126 x2.x5[7].floating.n125 0.003
R8700 x2.x5[7].floating.n123 x2.x5[7].floating.n122 0.00260608
R8701 x2.x5[7].floating.n156 x2.x5[7].floating.n155 0.00260608
R8702 x2.x5[7].floating.n61 x2.x5[7].floating.n60 0.00260608
R8703 x2.x5[7].floating.n91 x2.x5[7].floating.n90 0.00260608
R8704 x2.x5[7].floating.n144 x2.x5[7].floating.n143 0.00177054
R8705 x2.x5[7].floating.n49 x2.x5[7].floating.n48 0.00177054
R8706 x2.x5[7].floating.n79 x2.x5[7].floating.n78 0.00177054
R8707 x2.x5[7].floating.n109 x2.x5[7].floating.n108 0.00177054
R8708 x2.x5[7].floating.n145 x2.x5[7].floating.n144 0.00174992
R8709 x2.x5[7].floating.n50 x2.x5[7].floating.n49 0.00174992
R8710 x2.x5[7].floating.n80 x2.x5[7].floating.n79 0.00174992
R8711 x2.x5[7].floating.n110 x2.x5[7].floating.n109 0.00174992
R8712 x2.x5[7].floating.n124 x2.x5[7].floating.n123 0.00101477
R8713 x2.x5[7].floating.n157 x2.x5[7].floating.n156 0.00101477
R8714 x2.x5[7].floating.n62 x2.x5[7].floating.n61 0.00101477
R8715 x2.x5[7].floating.n92 x2.x5[7].floating.n91 0.00101477
R8716 x2.x5[7].floating.n158 x2.x5[7].floating.n157 0.00053972
R8717 x2.x5[7].floating.n146 x2.x5[7].floating.n145 0.00053972
R8718 x2.x5[7].floating.n111 x2.x5[7].floating.n110 0.00053972
R8719 x2.x5[7].floating.n93 x2.x5[7].floating.n92 0.00053972
R8720 x2.x5[7].floating.n81 x2.x5[7].floating.n80 0.00053972
R8721 x2.x5[7].floating.n63 x2.x5[7].floating.n62 0.00053972
R8722 x2.x5[7].floating.n51 x2.x5[7].floating.n50 0.00053972
R8723 x2.x5[7].floating.n125 x2.x5[7].floating.n124 0.00053972
R8724 async_setb_delay_ctrl_code[3].n0 async_setb_delay_ctrl_code[3].t1 229.971
R8725 async_setb_delay_ctrl_code[3].n0 async_setb_delay_ctrl_code[3].t0 158.35
R8726 async_setb_delay_ctrl_code[3].n1 async_setb_delay_ctrl_code[3].n0 8.50772
R8727 async_setb_delay_ctrl_code[3].n1 async_setb_delay_ctrl_code[3] 3.95264
R8728 async_setb_delay_ctrl_code[3].n2 async_setb_delay_ctrl_code[3].n1 1.73285
R8729 async_setb_delay_ctrl_code[3].n3 async_setb_delay_ctrl_code[3] 0.474765
R8730 async_setb_delay_ctrl_code[3] async_setb_delay_ctrl_code[3].n3 0.366977
R8731 async_setb_delay_ctrl_code[3].n2 async_setb_delay_ctrl_code[3] 0.339042
R8732 async_setb_delay_ctrl_code[3].n3 async_setb_delay_ctrl_code[3].n2 0.00334091
R8733 async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[1].t1 140.387
R8734 async_setb_delay_ctrl_code[1].n0 async_setb_delay_ctrl_code[1].t0 140.34
R8735 async_setb_delay_ctrl_code[1].n0 async_setb_delay_ctrl_code[1] 0.204648
R8736 async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[1].n0 0.00217851
R8737 async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[0].t0 140.343
C0 vdd x2.x10.Y 2.71f
C1 a_n397_736# x4.x9.output_stack 0.00892f
C2 a_1158_1098# a_n397_1077# 4.72e-20
C3 x4.x2.floating x4.x5[7].floating 0.441f
C4 x2.x6.SW a_n6270_n2738# 0.00707f
C5 x10.A x4.x5[7].floating 0.0208f
C6 a_n6207_137# x4.x7.floating 8.52e-19
C7 a_724_824# a_1094_824# 4.11e-20
C8 x2.x10.Y x9.Y 3.91e-20
C9 a_1094_824# eob 1.43e-20
C10 vdd a_n6295_n1763# 0.00423f
C11 a_n6207_137# async_resetb_delay_ctrl_code[2] 3.74e-19
C12 async_setb_delay_ctrl_code[2] ready 0.00844f
C13 async_clk_sar async_resetb_delay_ctrl_code[0] 2.74e-19
C14 vdd x4.x7.floating 0.0321f
C15 a_2077_824# a_1159_798# 0.0708f
C16 async_setb_delay_ctrl_code[1] x4.x9.output_stack 1.26e-20
C17 a_n6135_n1625# a_n6295_n1763# 0.0388f
C18 async_clk_sar a_n6135_137# 0.0135f
C19 x3.A0 x4.x9.output_stack 4.3e-19
C20 ready a_n6207_n1073# 2.42e-19
C21 a_618_824# a_1363_798# 0.199f
C22 x4.x10.Y x4.x7.floating 0.00345f
C23 vdd a_944_1775# 0.131f
C24 vdd async_resetb_delay_ctrl_code[2] 0.0376f
C25 async_setb_delay_ctrl_code[1] x2.x3[1].floating 0.227f
C26 async_setb_delay_ctrl_code[1] x2.x9.output_stack 0.0745f
C27 a_n6135_n139# x4.x6.SW 7.9e-20
C28 x2.x10.Y a_n397_n2289# 0.00127f
C29 async_setb_delay_ctrl_code[1] a_n6295_n277# 1.69e-20
C30 async_setb_delay_ctrl_code[0] x4.x2.floating 3.73e-20
C31 x3.X a_618_824# 4.42e-20
C32 x4.x10.Y async_resetb_delay_ctrl_code[2] 0.00203f
C33 delay_offset a_n6207_n1763# 0.00168f
C34 a_724_824# a_860_798# 0.0282f
C35 a_n6135_n139# delay_offset 0.00304f
C36 x2.x5[7].floating a_n6182_n2876# 0.00169f
C37 eob a_860_798# 0.00543f
C38 a_944_1775# x9.Y 0.00285f
C39 vdd a_n6270_n2738# 0.106f
C40 async_setb_delay_ctrl_code[1] x2.x6.floating 1.6e-19
C41 a_1577_1106# a_1363_798# 0.0104f
C42 x4.x2.floating a_618_824# 1.71e-19
C43 a_618_824# x10.A 8.37e-19
C44 eob a_1631_1008# 0.0119f
C45 a_n397_1077# a_305_798# 9.86e-19
C46 a_1094_1190# vdd 0.00433f
C47 vdd a_1771_1775# 0.111f
C48 x2.x7.floating x2.x9.output_stack 0.185f
C49 a_1159_798# a_1363_798# 0.117f
C50 a_n6135_413# a_n6135_137# 0.0316f
C51 a_n6295_275# a_n6207_275# 0.00227f
C52 a_1094_1190# x9.Y 3.7e-19
C53 async_setb_delay_ctrl_code[2] a_n6207_n1073# 5.73e-19
C54 x3.X a_1159_798# 0.00305f
C55 a_1771_1775# x9.Y 8.55e-19
C56 delay_offset a_n6270_n3014# 6.38e-19
C57 x2.x2.floating async_resetb_delay_ctrl_code[0] 3.73e-20
C58 x3.A0 a_1086_1582# 0.00164f
C59 a_818_1106# sample_clk 7.44e-22
C60 x2.x7.floating x2.x6.floating 0.202f
C61 a_n6135_n1073# a_n6135_n1349# 0.0316f
C62 a_n6295_n1211# a_n6207_n1211# 0.00227f
C63 async_setb_delay_ctrl_code[1] async_clk_sar 1.7e-19
C64 async_setb_delay_ctrl_code[0] a_n397_n1948# 0.00169f
C65 a_860_798# x4.x5[7].floating 2.17e-19
C66 a_1159_798# x10.A 2.36e-20
C67 a_n397_736# a_1158_1098# 3.77e-20
C68 a_n6295_n277# a_n6295_n935# 0.00472f
C69 async_clk_sar x3.A0 0.12f
C70 x2.x6.SW a_n6270_n3014# 9.98e-20
C71 x4.x9.output_stack x27.Q_N 2.83e-20
C72 delay_offset a_n6207_n797# 9.83e-19
C73 async_resetb_delay_ctrl_code[1] x4.x7.floating 2.24e-20
C74 x2.x3[1].floating x2.x5[7].floating 0.8f
C75 x2.x5[7].floating x2.x9.output_stack 1.19f
C76 vdd a_2200_1841# 0.166f
C77 a_1094_824# a_618_824# 2.87e-21
C78 a_1373_1841# a_1771_1775# 0.00281f
C79 vdd a_n6207_n1763# 1.29e-19
C80 vdd a_n6135_n139# 5.05e-19
C81 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[1] 1.12f
C82 a_n6295_n1763# a_n6207_n1625# 0.00227f
C83 x4.x6.SW x4.x5[7].floating 0.00138f
C84 x2.x7.floating a_n6207_n935# 8.52e-19
C85 x3.A0 a_1158_1098# 0.0026f
C86 ready a_n6135_n1349# 0.0135f
C87 x2.x6.floating x2.x5[7].floating 1.18f
C88 a_n6182_1940# x4.x9.output_stack 1.5e-19
C89 x4.x3[1].floating x4.x2.floating 1.17f
C90 a_n6182_1940# x4.x6.floating 0.0157f
C91 x3.A0 a_1307_1909# 1.14e-19
C92 a_n6182_1940# a_n6182_1664# 0.0316f
C93 x2.x10.Y a_n6182_n2876# 4.2e-19
C94 delay_offset x4.x5[7].floating 0.00308f
C95 x4.x7.floating x4.x4[3].floating 1.18f
C96 a_1298_824# eob 0.00138f
C97 x2.x5[7].floating a_n6182_n3152# 0.00154f
C98 a_n6207_n139# delay_offset 9.85e-19
C99 a_n6207_551# delay_offset 0.00157f
C100 async_resetb_delay_ctrl_code[2] x4.x4[3].floating 0.532f
C101 vdd a_n6270_n3014# 0.0364f
C102 a_618_824# a_860_798# 0.124f
C103 a_2077_824# a_1363_798# 6.99e-20
C104 async_setb_delay_ctrl_code[1] x2.x2.floating 0.0027f
C105 a_n6295_n935# a_n6207_n935# 0.00227f
C106 a_724_824# vdd 0.00629f
C107 a_n397_736# a_305_798# 9.33e-19
C108 vdd a_2134_1909# 4.56e-19
C109 vdd eob 0.965f
C110 a_618_824# a_1631_1008# 0.0633f
C111 async_setb_delay_ctrl_code[0] x4.x6.SW 3.98e-21
C112 a_n6295_275# a_n6295_n1# 0.0316f
C113 async_setb_delay_ctrl_code[0] delay_offset 0.00338f
C114 a_724_824# x9.Y 0.0147f
C115 eob x9.Y 0.0902f
C116 delay_offset a_n6270_n3290# 3.28e-19
C117 x3.A0 a_1913_1582# 0.00141f
C118 a_n397_n1948# x9.A 0.151f
C119 a_944_1775# sample_clk 7.43e-19
C120 a_n6295_n1211# a_n6295_n1487# 0.0316f
C121 x3.A0 a_305_798# 0.0099f
C122 a_860_798# a_1159_798# 0.0334f
C123 async_setb_delay_ctrl_code[0] x2.x6.SW 4.27e-21
C124 async_setb_delay_ctrl_code[0] x2.x4[3].floating 8.48e-20
C125 a_n6270_n2738# a_n6182_n2876# 0.0704f
C126 x2.x6.SW a_n6270_n3290# 5.11e-20
C127 x2.x10.Y x2.x9.output_stack 1.01f
C128 a_1159_798# a_1631_1008# 0.15f
C129 a_1158_1098# x27.Q_N 7.22e-21
C130 async_clk_sar a_n6182_1940# 0.0513f
C131 x2.x3[1].floating x2.x10.Y 0.00302f
C132 delay_offset a_n6135_n1073# 0.00304f
C133 vdd x4.x5[7].floating 44f
C134 vdd a_1086_1909# 6.56e-19
C135 a_1771_1775# a_1913_1909# 0.00783f
C136 a_1771_1775# sample_clk 0.328f
C137 x4.x10.Y x4.x5[7].floating 1.01f
C138 eob a_1373_1841# 0.219f
C139 x4.x9.output_stack x4.x7.floating 0.185f
C140 x2.x6.floating x2.x10.Y 0.0881f
C141 a_n6295_n1763# x2.x9.output_stack 0.0388f
C142 x4.x7.floating x4.x6.floating 0.202f
C143 a_1363_798# x10.A 3.1e-21
C144 x2.x7.floating a_n6295_n1211# 0.00409f
C145 x9.Y x4.x5[7].floating 1.94e-19
C146 x2.x6.SW a_n6135_n1073# 7.9e-20
C147 x2.x4[3].floating a_n6135_n1073# 7.47e-19
C148 a_1086_1909# x9.Y 2.99e-20
C149 ready a_n6207_n1349# 5.05e-19
C150 a_n6270_1526# x4.x6.SW 0.00707f
C151 x2.x2.floating x2.x5[7].floating 0.441f
C152 x4.x9.output_stack async_resetb_delay_ctrl_code[2] 0.335f
C153 eob a_210_798# 6.03e-19
C154 a_n6270_1802# x4.x5[7].floating 2.76e-19
C155 a_n6135_n139# x4.x4[3].floating 7.47e-19
C156 async_resetb_delay_ctrl_code[2] x4.x6.floating 1.72e-19
C157 a_n6295_n277# x4.x7.floating 0.00218f
C158 a_n6207_689# x4.x7.floating 8.52e-19
C159 x2.x10.Y a_n6182_n3152# 1.49e-19
C160 a_n6295_275# x4.x6.SW 8.11e-20
C161 a_n6270_1526# delay_offset 0.00273f
C162 a_724_824# x10.Y 3.78e-20
C163 eob x10.Y 7.72e-19
C164 async_resetb_delay_ctrl_code[2] x2.x9.output_stack 7.64e-21
C165 a_n6295_n277# async_resetb_delay_ctrl_code[2] 0.00555f
C166 a_1298_824# a_618_824# 3.73e-19
C167 a_n6207_689# async_resetb_delay_ctrl_code[2] 1.08e-19
C168 async_setb_delay_ctrl_code[0] vdd 0.00353f
C169 ready delay_offset 0.257f
C170 a_n6295_275# delay_offset 0.0159f
C171 a_n397_736# a_n397_1077# 0.0121f
C172 x4.x2.floating x10.A 0.0196f
C173 vdd a_n6270_n3290# 0.113f
C174 async_setb_delay_ctrl_code[0] x4.x10.Y 2.78e-20
C175 a_n6270_2078# x4.x5[7].floating 2.14e-19
C176 a_n6295_n935# a_n6295_n1211# 0.0316f
C177 vdd a_1403_1582# 0.00116f
C178 async_clk_sar a_n6207_n1# 2.42e-19
C179 a_n6270_n2738# x2.x9.output_stack 0.0702f
C180 sample_clk a_2200_1841# 0.237f
C181 x27.Q_N a_305_798# 0.124f
C182 async_setb_delay_ctrl_code[0] x9.Y 8.99e-21
C183 vdd a_618_824# 0.383f
C184 x2.x4[3].floating ready 6.65e-19
C185 x2.x6.SW ready 0.0928f
C186 a_1499_824# eob 0.00879f
C187 async_setb_delay_ctrl_code[2] a_n6207_n1349# 2.57e-19
C188 vdd a_n6135_n1073# 5.05e-19
C189 a_210_798# x4.x5[7].floating 9.95e-19
C190 x2.x6.floating a_n6270_n2738# 0.00996f
C191 x3.A0 a_n397_1077# 0.0102f
C192 a_618_824# x9.Y 0.0969f
C193 a_944_1775# a_1086_1582# 0.00557f
C194 a_1298_824# a_1159_798# 2.56e-19
C195 a_2077_824# a_1631_1008# 0.0367f
C196 x4.x5[7].floating x10.Y 0.00121f
C197 a_1577_1106# vdd 0.0108f
C198 a_818_1106# a_305_798# 0.00945f
C199 async_clk_sar x4.x7.floating 0.0241f
C200 async_resetb_delay_ctrl_code[1] x4.x5[7].floating 0.00228f
C201 async_setb_delay_ctrl_code[2] delay_offset 0.0282f
C202 a_n6182_n2876# a_n6270_n3014# 0.0704f
C203 async_clk_sar a_944_1775# 0.0812f
C204 async_clk_sar async_resetb_delay_ctrl_code[2] 0.00848f
C205 a_n397_736# async_resetb_delay_ctrl_code[0] 0.00169f
C206 vdd a_1159_798# 0.941f
C207 delay_offset a_n6207_n1073# 0.00105f
C208 x4.x2.floating a_1094_824# 1.94e-20
C209 vdd a_n6270_1526# 0.104f
C210 sample_clk a_2134_1909# 6.34e-19
C211 a_1296_1190# eob 0.00273f
C212 async_setb_delay_ctrl_code[2] x2.x6.SW 9.9e-21
C213 async_setb_delay_ctrl_code[2] x2.x4[3].floating 0.532f
C214 eob sample_clk 0.0556f
C215 a_n6135_n139# x4.x9.output_stack 8.05e-20
C216 a_1373_1841# a_618_824# 2.95e-19
C217 vdd ready 0.342f
C218 a_n6270_1526# x4.x10.Y 0.039f
C219 a_n6135_n139# x4.x6.floating 0.00109f
C220 vdd a_n6295_275# 0.00308f
C221 x2.x2.floating x2.x10.Y 0.00202f
C222 a_860_798# a_1363_798# 0.00187f
C223 x9.Y a_1159_798# 0.0137f
C224 a_n6207_n1763# x2.x9.output_stack 0.00227f
C225 x4.x4[3].floating x4.x5[7].floating 1.55f
C226 x2.x7.floating a_n6207_n1211# 8.52e-19
C227 ready a_n6135_n1625# 0.0135f
C228 a_n6295_275# x4.x10.Y 6.65e-20
C229 x3.X a_860_798# 1.39e-19
C230 async_clk_sar a_1771_1775# 8.97e-20
C231 a_944_1775# a_1158_1098# 7.04e-20
C232 a_n6135_n139# a_n6295_n277# 0.0388f
C233 a_1363_798# a_1631_1008# 0.205f
C234 async_setb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1] 3.47e-20
C235 async_setb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[0] 3.47e-20
C236 a_n6270_1802# a_n6270_1526# 0.0316f
C237 a_618_824# a_210_798# 6.04e-19
C238 x9.A vdd 0.386f
C239 a_n6135_413# x4.x7.floating 0.00959f
C240 x3.X a_1631_1008# 5.15e-20
C241 x4.x3[1].floating vdd 0.0301f
C242 a_618_824# x10.Y 0.0947f
C243 a_n6207_n277# async_resetb_delay_ctrl_code[2] 0.00134f
C244 a_860_798# x10.A 8.46e-20
C245 x4.x2.floating a_860_798# 4.32e-20
C246 x4.x3[1].floating x4.x10.Y 0.00302f
C247 a_n6207_275# delay_offset 0.00125f
C248 x9.A x9.Y 0.077f
C249 a_724_824# x4.x9.output_stack 2.57e-20
C250 a_1094_1190# a_1158_1098# 2.13e-19
C251 x27.Q_N a_n397_1077# 3.71e-19
C252 vdd a_2230_1582# 8.63e-19
C253 a_1771_1775# a_1158_1098# 1.33e-19
C254 a_1373_1841# a_1159_798# 6.83e-20
C255 async_setb_delay_ctrl_code[0] x4.x4[3].floating 7.6e-20
C256 x2.x7.floating async_resetb_delay_ctrl_code[0] 1.9e-20
C257 x2.x10.Y a_n6295_n1211# 4.07e-20
C258 sample_clk a_1086_1909# 1.02e-19
C259 async_setb_delay_ctrl_code[2] vdd 0.0376f
C260 a_1499_824# a_618_824# 0.00943f
C261 a_1159_798# a_210_798# 1.03e-19
C262 x2.x6.floating a_n6270_n3014# 0.00996f
C263 a_818_1106# a_n397_1077# 8.77e-20
C264 x9.A a_n397_n2289# 0.147f
C265 async_clk_sar a_2200_1841# 7.41e-21
C266 a_n397_736# x3.A0 0.00125f
C267 a_1159_798# x10.Y 2.18e-19
C268 a_n6135_n1349# a_n6207_n1349# 0.00227f
C269 async_clk_sar a_n6135_n139# 0.0135f
C270 a_2077_824# vdd 0.257f
C271 a_944_1775# a_305_798# 3.86e-20
C272 async_resetb_delay_ctrl_code[0] a_n6295_n935# 1.94e-19
C273 a_n6295_551# x4.x7.floating 0.00409f
C274 a_n6270_n3014# a_n6182_n3152# 0.0704f
C275 a_1875_824# eob 4.69e-19
C276 a_n6295_551# async_resetb_delay_ctrl_code[2] 3.81e-20
C277 ready async_resetb_delay_ctrl_code[1] 1.7e-19
C278 delay_offset a_n6135_n1349# 0.00347f
C279 a_1094_824# a_860_798# 0.00707f
C280 a_2077_824# x9.Y 2.45e-20
C281 x4.x9.output_stack x4.x5[7].floating 1.19f
C282 x4.x6.floating x4.x5[7].floating 1.18f
C283 a_2200_1841# a_1158_1098# 5.86e-19
C284 x2.x5[7].floating async_resetb_delay_ctrl_code[0] 1.38e-20
C285 a_n6182_1664# x4.x5[7].floating 0.00169f
C286 a_1771_1775# a_1913_1582# 0.00557f
C287 eob a_1086_1582# 0.00746f
C288 a_1499_824# a_1159_798# 6.04e-20
C289 a_1298_824# a_1363_798# 9.75e-19
C290 a_1296_1190# a_618_824# 0.00652f
C291 a_1094_1190# a_305_798# 7.71e-20
C292 sample_clk a_618_824# 0.00227f
C293 x2.x7.floating a_n6295_n1487# 0.00409f
C294 x2.x6.SW a_n6135_n1349# 1.28e-19
C295 x4.x3[1].floating async_resetb_delay_ctrl_code[1] 0.227f
C296 x2.x4[3].floating a_n6135_n1349# 8.29e-19
C297 ready a_n6207_n1625# 0.0013f
C298 async_clk_sar a_2134_1909# 2.27e-20
C299 a_n6295_n277# a_n6207_n139# 0.00227f
C300 async_clk_sar eob 0.0105f
C301 vdd a_1363_798# 0.33f
C302 async_setb_delay_ctrl_code[1] x2.x7.floating 2.24e-20
C303 a_n6207_413# x4.x7.floating 8.52e-19
C304 a_n6295_275# x4.x4[3].floating 1.17e-19
C305 a_n6295_n1# x4.x6.SW 4.74e-20
C306 a_1577_1106# sample_clk 2.8e-19
C307 vdd x3.X 0.281f
C308 async_setb_delay_ctrl_code[0] x4.x9.output_stack 2.59e-20
C309 async_clk_sar a_n6207_n797# 6.27e-21
C310 a_n6207_413# async_resetb_delay_ctrl_code[2] 1.86e-19
C311 async_setb_delay_ctrl_code[0] x4.x6.floating 1.3e-21
C312 a_n6295_n1# delay_offset 0.0151f
C313 x9.Y a_1363_798# 0.176f
C314 async_setb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[1] 6.4e-20
C315 x4.x3[1].floating x4.x4[3].floating 1.19f
C316 async_setb_delay_ctrl_code[0] x2.x3[1].floating 0.0427f
C317 async_setb_delay_ctrl_code[0] x2.x9.output_stack 0.0322f
C318 a_n397_736# x27.Q_N 4.64e-19
C319 a_1296_1190# a_1159_798# 0.00907f
C320 eob a_1158_1098# 0.0353f
C321 sample_clk a_1159_798# 0.33f
C322 vdd x10.A 0.397f
C323 async_setb_delay_ctrl_code[0] a_n6295_n277# 3.28e-20
C324 x3.X x9.Y 6.58e-19
C325 x4.x2.floating vdd 0.0341f
C326 a_1086_1582# x4.x5[7].floating 1.63e-21
C327 ready a_n6182_n2876# 0.00921f
C328 x4.x9.output_stack a_618_824# 1.97e-20
C329 x4.x10.Y x10.A 1.13e-19
C330 async_setb_delay_ctrl_code[1] a_n6295_n935# 6.64e-20
C331 x4.x2.floating x4.x10.Y 0.00202f
C332 a_2077_824# x10.Y 4.26e-21
C333 async_setb_delay_ctrl_code[0] x2.x6.floating 1.49e-19
C334 x9.Y x10.A 0.00132f
C335 async_setb_delay_ctrl_code[2] a_n6207_n1625# 1.39e-19
C336 x4.x2.floating x9.Y 1.03e-19
C337 vdd a_n6135_n1349# 5.05e-19
C338 async_clk_sar x4.x5[7].floating 0.00554f
C339 x2.x6.floating a_n6270_n3290# 0.00578f
C340 async_clk_sar a_1086_1909# 0.00113f
C341 async_setb_delay_ctrl_code[2] x4.x4[3].floating 3.3e-20
C342 async_setb_delay_ctrl_code[1] x2.x5[7].floating 0.00228f
C343 a_n6135_n1073# x2.x9.output_stack 8.05e-20
C344 a_n6135_n1349# a_n6135_n1625# 0.0316f
C345 a_n6295_n1487# a_n6207_n1487# 0.00227f
C346 async_clk_sar a_n6207_n139# 1.8e-19
C347 x3.A0 x27.Q_N 0.00321f
C348 a_1373_1841# a_1363_798# 0.00107f
C349 async_clk_sar a_n6207_551# 0.0013f
C350 x2.x7.floating a_n6295_n935# 0.00218f
C351 a_n6182_n3152# a_n6270_n3290# 0.0704f
C352 x3.X a_1373_1841# 0.216f
C353 x2.x10.Y async_resetb_delay_ctrl_code[0] 2.78e-20
C354 a_n6295_n1# a_n6207_137# 0.00227f
C355 delay_offset a_n6207_n1349# 0.00125f
C356 x2.x6.floating a_n6135_n1073# 0.00109f
C357 a_n6270_1526# x4.x9.output_stack 0.0702f
C358 a_1094_1190# a_n397_1077# 2.38e-20
C359 x2.x7.floating x2.x5[7].floating 0.182f
C360 a_n6270_1526# x4.x6.floating 0.00996f
C361 delay_offset x4.x6.SW 0.19f
C362 sample_clk a_2230_1582# 0.00576f
C363 a_818_1106# x3.A0 4.68e-19
C364 eob a_1913_1582# 6.99e-19
C365 a_1363_798# x10.Y 2.07e-20
C366 a_n6182_1664# a_n6270_1526# 0.0704f
C367 async_setb_delay_ctrl_code[0] async_clk_sar 2.16e-19
C368 a_n397_n1948# vdd 0.235f
C369 a_1094_824# vdd 1.71e-19
C370 a_724_824# a_305_798# 0.0397f
C371 vdd a_n6295_n1# 0.00308f
C372 eob a_305_798# 0.00665f
C373 x2.x7.floating a_n6207_n1487# 8.52e-19
C374 ready x2.x9.output_stack 0.37f
C375 a_n6295_n1# x4.x10.Y 4.07e-20
C376 x4.x2.floating a_210_798# 4.53e-19
C377 x10.A a_210_798# 0.0154f
C378 async_resetb_delay_ctrl_code[0] x4.x7.floating 2.06e-20
C379 a_n397_n1948# x9.Y 0.00338f
C380 async_clk_sar a_618_824# 2.66e-19
C381 a_n6207_551# a_n6135_413# 0.00227f
C382 a_1094_824# x9.Y 0.00148f
C383 a_1298_824# a_860_798# 0.00276f
C384 x4.x3[1].floating x4.x9.output_stack 0.341f
C385 a_n6135_137# x4.x7.floating 0.00959f
C386 x10.A x10.Y 0.0733f
C387 x4.x2.floating x10.Y 5.97e-19
C388 async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[0] 7.32e-19
C389 a_2077_824# sample_clk 0.00445f
C390 a_1875_1190# eob 6.51e-19
C391 x9.A x2.x9.output_stack 0.127f
C392 x2.x6.SW delay_offset 0.19f
C393 async_resetb_delay_ctrl_code[1] x10.A 5.47e-22
C394 a_1499_824# a_1363_798# 0.07f
C395 x2.x4[3].floating delay_offset 0.00498f
C396 x4.x2.floating async_resetb_delay_ctrl_code[1] 0.0027f
C397 x2.x6.floating ready 0.0299f
C398 a_n6207_n935# a_n6135_n1073# 0.00227f
C399 vdd a_860_798# 0.199f
C400 a_n397_n1948# a_n397_n2289# 0.0121f
C401 x2.x10.Y a_n6295_n1487# 6.65e-20
C402 ready a_n6182_n3152# 0.00847f
C403 a_618_824# a_1158_1098# 0.139f
C404 async_setb_delay_ctrl_code[2] x4.x9.output_stack 7.64e-21
C405 vdd a_1631_1008# 0.187f
C406 x4.x5[7].floating a_305_798# 0.00217f
C407 async_setb_delay_ctrl_code[1] x2.x10.Y 7.05e-19
C408 a_860_798# x9.Y 0.175f
C409 async_setb_delay_ctrl_code[2] x2.x3[1].floating 0.00115f
C410 async_setb_delay_ctrl_code[2] x2.x9.output_stack 0.335f
C411 async_setb_delay_ctrl_code[0] x2.x2.floating 0.164f
C412 a_n6207_137# delay_offset 0.00113f
C413 async_clk_sar a_n6270_1526# 0.0469f
C414 async_setb_delay_ctrl_code[2] a_n6295_n277# 1.43e-20
C415 x9.Y a_1631_1008# 0.138f
C416 vdd x4.x6.SW 0.431f
C417 a_n6295_n1487# a_n6295_n1763# 0.0316f
C418 a_818_1106# x27.Q_N 2.02e-20
C419 a_1577_1106# a_1158_1098# 2.46e-19
C420 a_1296_1190# a_1363_798# 9.46e-19
C421 sample_clk a_1363_798# 0.00277f
C422 async_clk_sar ready 0.00254f
C423 async_clk_sar a_n6295_275# 0.0136f
C424 ready a_n6207_n935# 1.8e-19
C425 a_n6295_551# a_n6207_551# 0.00227f
C426 x3.X a_1913_1909# 8.96e-19
C427 x4.x10.Y x4.x6.SW 0.788f
C428 async_setb_delay_ctrl_code[2] x2.x6.floating 1.72e-19
C429 x3.X sample_clk 0.0119f
C430 vdd delay_offset 0.484f
C431 a_1158_1098# a_1159_798# 0.796f
C432 x2.x7.floating x2.x10.Y 0.00345f
C433 delay_offset x4.x10.Y 0.0402f
C434 async_setb_delay_ctrl_code[1] x4.x7.floating 1.76e-20
C435 delay_offset a_n6135_n1625# 0.00561f
C436 a_n6270_1802# x4.x6.SW 9.98e-20
C437 async_setb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[2] 6.4e-20
C438 x2.x6.SW vdd 0.432f
C439 a_944_1775# x3.A0 0.0607f
C440 x2.x4[3].floating vdd 0.0565f
C441 a_1373_1841# a_1631_1008# 5.16e-19
C442 a_n6270_1802# delay_offset 6.38e-19
C443 x2.x6.SW a_n6135_n1625# 2.44e-19
C444 a_618_824# a_305_798# 0.273f
C445 x2.x4[3].floating a_n6135_n1625# 8.29e-19
C446 x2.x7.floating a_n6295_n1763# 0.00409f
C447 a_1094_824# a_1499_824# 2.46e-21
C448 a_2077_824# a_1875_824# 3.67e-19
C449 a_n6207_n277# ready 6.27e-21
C450 a_n6135_137# a_n6135_n139# 0.0316f
C451 x2.x10.Y a_n6295_n935# 2.2e-20
C452 a_n6135_413# a_n6295_275# 0.0388f
C453 a_n6270_2078# x4.x6.SW 5.11e-20
C454 a_860_798# x10.Y 0.00138f
C455 a_n6295_n1# x4.x4[3].floating 1.17e-19
C456 async_setb_delay_ctrl_code[2] async_clk_sar 1.35e-19
C457 async_setb_delay_ctrl_code[2] a_n6207_n935# 9.05e-19
C458 a_1094_1190# x3.A0 2.77e-19
C459 x2.x7.floating async_resetb_delay_ctrl_code[2] 1.63e-20
C460 a_n6270_2078# delay_offset 3.28e-19
C461 a_1771_1775# x3.A0 0.112f
C462 a_1631_1008# x10.Y 2.45e-20
C463 a_n6135_n1073# a_n6295_n1211# 0.0388f
C464 x2.x10.Y x2.x5[7].floating 1.01f
C465 a_1298_824# vdd 0.00255f
C466 x4.x9.output_stack x10.A 0.127f
C467 x4.x2.floating x4.x9.output_stack 0.193f
C468 a_n397_1077# x4.x5[7].floating 0.0129f
C469 x2.x2.floating x9.A 0.0195f
C470 a_1298_824# x9.Y 0.00519f
C471 a_1159_798# a_305_798# 0.0492f
C472 a_1499_824# a_860_798# 0.00316f
C473 x4.x6.SW async_resetb_delay_ctrl_code[1] 7.41e-21
C474 async_resetb_delay_ctrl_code[2] a_n6295_n935# 1.43e-20
C475 a_1499_824# a_1631_1008# 0.0258f
C476 vdd a_n6135_n1625# 5.05e-19
C477 vdd x4.x10.Y 2.71f
C478 delay_offset async_resetb_delay_ctrl_code[1] 0.00331f
C479 vdd x9.Y 0.402f
C480 a_1875_1190# a_1159_798# 0.0018f
C481 a_2077_824# a_1158_1098# 0.163f
C482 a_n6135_n1349# x2.x9.output_stack 1.74e-19
C483 ready a_n6295_n1211# 0.0136f
C484 async_clk_sar a_n6207_275# 5.05e-19
C485 a_n6295_551# a_n6295_275# 0.0316f
C486 vdd a_n6270_1802# 0.035f
C487 x3.A0 a_2200_1841# 0.0396f
C488 x4.x3[1].floating a_305_798# 8.69e-21
C489 a_n6270_1802# x4.x10.Y 2.35e-19
C490 x2.x4[3].floating async_resetb_delay_ctrl_code[1] 7.03e-20
C491 delay_offset a_n6207_n1625# 0.00157f
C492 x2.x6.floating a_n6135_n1349# 0.00167f
C493 a_1296_1190# a_860_798# 0.00412f
C494 x2.x5[7].floating a_n6270_n2738# 2.76e-19
C495 sample_clk a_860_798# 3.22e-20
C496 a_n397_736# a_724_824# 4.86e-19
C497 delay_offset x4.x4[3].floating 0.00498f
C498 async_clk_sar x3.X 0.00553f
C499 vdd a_n397_n2289# 0.256f
C500 async_resetb_delay_ctrl_code[0] x4.x5[7].floating 0.00132f
C501 vdd a_n6270_2078# 0.111f
C502 a_618_824# a_n397_1077# 0.00171f
C503 sample_clk a_1631_1008# 0.00363f
C504 vdd a_1373_1841# 0.173f
C505 a_n6270_2078# x4.x10.Y 1.02e-19
C506 a_n397_n1948# x2.x3[1].floating 3.09e-19
C507 x2.x7.floating a_n6207_n1763# 8.52e-19
C508 a_n397_n1948# x2.x9.output_stack 0.00892f
C509 async_clk_sar x10.A 9.25e-19
C510 x4.x2.floating async_clk_sar 1.96e-21
C511 a_n397_n2289# x9.Y 0.00414f
C512 a_n6295_n1# a_n6295_n277# 0.0316f
C513 a_1158_1098# a_1363_798# 0.153f
C514 a_n6295_275# a_n6207_413# 0.00227f
C515 async_setb_delay_ctrl_code[2] a_n6295_n1211# 1.46e-19
C516 x3.X a_1158_1098# 0.00269f
C517 vdd a_210_798# 0.209f
C518 a_1373_1841# x9.Y 2.64e-20
C519 delay_offset a_n6182_n2876# 3.64e-19
C520 a_n6270_2078# a_n6270_1802# 0.0316f
C521 x3.A0 a_2134_1909# 0.0037f
C522 x3.X a_1307_1909# 0.0057f
C523 eob x3.A0 0.103f
C524 x4.x10.Y a_210_798# 1.19e-20
C525 a_n6295_n1211# a_n6207_n1073# 0.00227f
C526 vdd x10.Y 0.352f
C527 async_setb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[0] 2.95f
C528 x4.x9.output_stack a_860_798# 7.88e-21
C529 vdd async_resetb_delay_ctrl_code[1] 0.0184f
C530 a_1158_1098# x10.A 7.05e-20
C531 x9.Y a_210_798# 0.00119f
C532 a_1159_798# a_n397_1077# 0.00104f
C533 x4.x10.Y x10.Y 3.91e-20
C534 a_1298_824# a_1499_824# 3.34e-19
C535 x4.x10.Y async_resetb_delay_ctrl_code[1] 7.05e-19
C536 x2.x10.Y a_n6295_n1763# 1.69e-19
C537 a_n6207_n1# x4.x7.floating 8.52e-19
C538 x9.Y x10.Y 0.0036f
C539 a_1875_1190# a_2077_824# 8.94e-19
C540 a_n6207_n1# async_resetb_delay_ctrl_code[2] 5.73e-19
C541 a_1499_824# vdd 0.00369f
C542 x4.x6.SW x4.x9.output_stack 0.163f
C543 vdd x4.x4[3].floating 0.0565f
C544 a_n6135_n1625# a_n6207_n1625# 0.00227f
C545 x4.x6.SW x4.x6.floating 0.13f
C546 ready a_n6207_n1211# 3.4e-19
C547 async_clk_sar a_n6295_n1# 0.0136f
C548 x3.A0 x4.x5[7].floating 0.00349f
C549 x4.x10.Y x4.x4[3].floating 0.00668f
C550 delay_offset x4.x9.output_stack 0.256f
C551 x3.A0 a_1086_1909# 0.00118f
C552 a_1499_824# x9.Y 0.0336f
C553 x2.x10.Y a_n6270_n2738# 0.039f
C554 a_n6295_n277# x4.x6.SW 3.1e-20
C555 delay_offset x4.x6.floating 0.0624f
C556 a_n6182_1664# delay_offset 1.97e-19
C557 a_1875_824# a_1631_1008# 0.00812f
C558 delay_offset x2.x9.output_stack 0.256f
C559 x2.x5[7].floating a_n6270_n3014# 2.76e-19
C560 a_n6295_n277# delay_offset 0.0149f
C561 a_n6207_689# delay_offset 0.00168f
C562 async_resetb_delay_ctrl_code[2] x4.x7.floating 0.0177f
C563 vdd a_n6182_n2876# 0.0766f
C564 a_1875_1190# a_1363_798# 6.69e-20
C565 a_n397_736# a_618_824# 3.64e-19
C566 a_n6295_n935# a_n6207_n797# 0.0022f
C567 x4.x2.floating a_305_798# 5.99e-19
C568 eob x27.Q_N 4.98e-19
C569 a_210_798# x10.Y 0.066f
C570 a_1296_1190# vdd 0.0197f
C571 x10.A a_305_798# 4.94e-19
C572 vdd sample_clk 0.93f
C573 async_clk_sar a_860_798# 3.05e-19
C574 x2.x6.floating delay_offset 0.0624f
C575 x2.x6.SW x2.x9.output_stack 0.164f
C576 x2.x4[3].floating x2.x3[1].floating 1.19f
C577 x2.x4[3].floating x2.x9.output_stack 0.636f
C578 ready async_resetb_delay_ctrl_code[0] 2.16e-19
C579 async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[0] 2.53f
C580 a_n6295_275# a_n6135_137# 0.0388f
C581 async_setb_delay_ctrl_code[2] a_n6207_n1211# 3.74e-19
C582 sample_clk x9.Y 5.97e-19
C583 delay_offset a_n6182_n3152# 1.9e-19
C584 x2.x6.SW x2.x6.floating 0.13f
C585 x3.A0 a_1403_1582# 7.81e-19
C586 a_818_1106# eob 3.74e-19
C587 a_n397_n1948# x2.x2.floating 0.0104f
C588 x4.x3[1].floating async_resetb_delay_ctrl_code[0] 0.0427f
C589 a_944_1775# a_1771_1775# 5.22e-19
C590 a_n6295_n1211# a_n6135_n1349# 0.0388f
C591 x3.A0 a_618_824# 8.32e-19
C592 a_860_798# a_1158_1098# 0.137f
C593 async_clk_sar x4.x6.SW 0.0958f
C594 async_setb_delay_ctrl_code[0] x2.x7.floating 2.06e-20
C595 a_n397_736# a_1159_798# 2.71e-20
C596 a_n6207_n1# a_n6135_n139# 0.00227f
C597 a_1158_1098# a_1631_1008# 0.155f
C598 delay_offset a_n6207_n935# 9.85e-19
C599 async_clk_sar delay_offset 0.261f
C600 x27.Q_N x4.x5[7].floating 4.84e-19
C601 vdd x4.x9.output_stack 0.606f
C602 vdd x4.x6.floating 5.78f
C603 async_resetb_delay_ctrl_code[1] x4.x4[3].floating 0.0302f
C604 x4.x10.Y x4.x9.output_stack 1.01f
C605 vdd a_n6182_1664# 0.0715f
C606 a_1577_1106# x3.A0 6.05e-20
C607 async_setb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[0] 6.95e-20
C608 a_1373_1841# sample_clk 0.00307f
C609 x4.x10.Y x4.x6.floating 0.0881f
C610 x2.x3[1].floating vdd 0.0301f
C611 vdd x2.x9.output_stack 0.6f
C612 a_1094_824# a_305_798# 4.2e-20
C613 a_n6182_1664# x4.x10.Y 4.2e-19
C614 vdd a_n6295_n277# 0.00308f
C615 vdd a_n6207_689# 1.29e-19
C616 x4.x9.output_stack x9.Y 1.22e-19
C617 a_n6135_n1625# x2.x9.output_stack 0.032f
C618 a_n6295_n1763# a_n6207_n1763# 0.00227f
C619 a_1363_798# a_n397_1077# 7.84e-21
C620 x2.x7.floating a_n6135_n1073# 0.00925f
C621 a_n6295_n277# x4.x10.Y 2.2e-20
C622 async_setb_delay_ctrl_code[0] a_n6295_n935# 2.48e-19
C623 x3.A0 a_1159_798# 0.00192f
C624 ready a_n6295_n1487# 0.0136f
C625 a_818_1106# x4.x5[7].floating 1.4e-19
C626 x4.x3[1].floating a_n397_736# 3.09e-19
C627 a_n6182_1940# x4.x5[7].floating 0.00154f
C628 x9.Y x2.x9.output_stack 6.94e-19
C629 a_n6270_1802# x4.x6.floating 0.00996f
C630 a_n6270_1802# a_n6182_1664# 0.0704f
C631 x2.x6.floating vdd 5.9f
C632 a_n6135_n139# x4.x7.floating 0.00925f
C633 x2.x10.Y a_n6270_n3014# 2.35e-19
C634 a_n6135_413# x4.x6.SW 2.44e-19
C635 async_setb_delay_ctrl_code[1] ready 3.39e-19
C636 async_setb_delay_ctrl_code[0] x2.x5[7].floating 0.00132f
C637 x2.x6.floating a_n6135_n1625# 0.00278f
C638 a_n6207_n277# delay_offset 9.83e-19
C639 x2.x5[7].floating a_n6270_n3290# 2.14e-19
C640 a_n6135_413# delay_offset 0.00561f
C641 a_n397_1077# x10.A 0.146f
C642 vdd a_n6182_n3152# 0.131f
C643 a_860_798# a_305_798# 0.197f
C644 async_setb_delay_ctrl_code[1] x9.A 5.47e-22
C645 a_n6270_2078# x4.x6.floating 0.00578f
C646 a_n6295_n935# a_n6135_n1073# 0.0388f
C647 async_setb_delay_ctrl_code[1] x4.x3[1].floating 3.44e-20
C648 vdd a_1086_1582# 0.00267f
C649 async_clk_sar a_n6207_137# 3.4e-19
C650 a_n397_n2289# x2.x9.output_stack 0.00887f
C651 a_618_824# x27.Q_N 0.00553f
C652 a_1631_1008# a_305_798# 4.7e-22
C653 a_1875_824# x9.Y 7.76e-21
C654 x2.x7.floating ready 0.0241f
C655 a_n6207_275# a_n6135_137# 0.00227f
C656 async_setb_delay_ctrl_code[2] a_n6295_n1487# 6.81e-20
C657 x4.x9.output_stack a_210_798# 3.94e-20
C658 x9.Y a_1086_1582# 1.74e-19
C659 vdd async_clk_sar 3.21f
C660 a_724_824# a_944_1775# 1.17e-20
C661 async_clk_sar x4.x10.Y 0.11f
C662 x4.x9.output_stack x10.Y 6.58e-19
C663 a_1875_1190# a_1631_1008# 0.00972f
C664 a_1298_824# a_1158_1098# 0.00126f
C665 a_n6207_n1211# a_n6135_n1349# 0.00227f
C666 a_944_1775# eob 0.324f
C667 a_818_1106# a_618_824# 0.00185f
C668 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[1] 1.12f
C669 x4.x9.output_stack async_resetb_delay_ctrl_code[1] 0.0745f
C670 a_n6295_551# x4.x6.SW 0.00179f
C671 async_resetb_delay_ctrl_code[1] x4.x6.floating 1.6e-19
C672 a_n6270_n2738# a_n6270_n3014# 0.0316f
C673 ready a_n6295_n935# 0.0127f
C674 a_1159_798# x27.Q_N 1.07e-19
C675 async_clk_sar a_n6270_1802# 0.0381f
C676 x2.x3[1].floating async_resetb_delay_ctrl_code[1] 3.44e-20
C677 async_resetb_delay_ctrl_code[1] x2.x9.output_stack 1.26e-20
C678 async_resetb_delay_ctrl_code[0] x10.A 4.44e-19
C679 vdd a_1158_1098# 0.38f
C680 x4.x2.floating async_resetb_delay_ctrl_code[0] 0.164f
C681 delay_offset a_n6295_n1211# 0.0151f
C682 a_n6295_n277# async_resetb_delay_ctrl_code[1] 5.54e-20
C683 a_n6295_551# delay_offset 0.0311f
C684 vdd a_1307_1909# 5.08e-19
C685 a_1296_1190# sample_clk 6.91e-21
C686 a_2077_824# x3.A0 1.98e-19
C687 a_1094_1190# eob 5.14e-19
C688 sample_clk a_1913_1909# 4.4e-19
C689 ready x2.x5[7].floating 0.00127f
C690 eob a_1771_1775# 0.0171f
C691 async_setb_delay_ctrl_code[2] x2.x7.floating 0.0177f
C692 x4.x9.output_stack x4.x4[3].floating 0.636f
C693 x9.Y a_1158_1098# 0.313f
C694 vdd a_n6135_413# 5.05e-19
C695 x4.x7.floating x4.x5[7].floating 0.182f
C696 a_n397_736# a_1363_798# 2.96e-20
C697 x2.x4[3].floating a_n6295_n1211# 1.17e-19
C698 x2.x7.floating a_n6207_n1073# 8.52e-19
C699 x2.x6.SW a_n6295_n1211# 4.74e-20
C700 a_818_1106# a_1159_798# 1.25e-19
C701 async_clk_sar a_n6270_2078# 0.0377f
C702 ready a_n6207_n1487# 7.93e-19
C703 async_clk_sar a_1373_1841# 8.61e-20
C704 x9.A x2.x5[7].floating 0.0208f
C705 a_944_1775# x4.x5[7].floating 6.23e-19
C706 async_setb_delay_ctrl_code[0] x2.x10.Y 0.0125f
C707 async_resetb_delay_ctrl_code[2] x4.x5[7].floating 0.00564f
C708 a_n6207_n139# x4.x7.floating 8.52e-19
C709 a_944_1775# a_1086_1909# 0.00783f
C710 a_n6295_n277# x4.x4[3].floating 7.17e-20
C711 x2.x2.floating vdd 0.0334f
C712 x2.x10.Y a_n6270_n3290# 1.02e-19
C713 a_n6207_551# x4.x7.floating 8.52e-19
C714 a_n6207_n139# async_resetb_delay_ctrl_code[2] 9.05e-19
C715 a_860_798# a_n397_1077# 1.21e-19
C716 a_n6207_551# async_resetb_delay_ctrl_code[2] 1.39e-19
C717 async_setb_delay_ctrl_code[2] a_n6295_n935# 0.00555f
C718 a_n6207_413# delay_offset 0.0014f
C719 async_clk_sar a_210_798# 1.47e-20
C720 x4.x2.floating a_n397_736# 0.0104f
C721 a_n397_736# x10.A 0.151f
C722 x2.x2.floating x9.Y 4.13e-19
C723 async_clk_sar x10.Y 1.48e-20
C724 x3.A0 a_1363_798# 2.86e-19
C725 vdd a_1913_1582# 0.00177f
C726 a_1373_1841# a_1158_1098# 3.86e-20
C727 a_1094_1190# x4.x5[7].floating 3.47e-20
C728 a_n6182_n2876# x2.x9.output_stack 0.032f
C729 async_setb_delay_ctrl_code[2] x2.x5[7].floating 0.00564f
C730 async_setb_delay_ctrl_code[0] x4.x7.floating 1.9e-20
C731 async_clk_sar async_resetb_delay_ctrl_code[1] 3.58e-19
C732 x3.X x3.A0 0.199f
C733 eob a_2200_1841# 2.37e-19
C734 vdd a_305_798# 0.615f
C735 a_n6135_137# a_n6295_n1# 0.0388f
C736 async_setb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[2] 6.95e-20
C737 async_setb_delay_ctrl_code[2] a_n6207_n1487# 1.86e-19
C738 x4.x10.Y a_305_798# 3.56e-22
C739 a_1158_1098# a_210_798# 1.73e-20
C740 vdd a_n6295_n1211# 0.00308f
C741 a_n6295_551# vdd 0.00423f
C742 x2.x6.floating a_n6182_n2876# 0.0194f
C743 x3.A0 x10.A 0.00259f
C744 x4.x2.floating x3.A0 3.14e-19
C745 a_944_1775# a_1403_1582# 6.64e-19
C746 x9.Y a_305_798# 0.145f
C747 a_n6295_551# x4.x10.Y 1.69e-19
C748 a_1158_1098# x10.Y 0.00321f
C749 a_n6135_n1349# a_n6295_n1487# 0.0388f
C750 a_1875_1190# vdd 0.0042f
C751 a_944_1775# a_618_824# 2.2e-20
C752 async_clk_sar x4.x4[3].floating 6.65e-19
C753 a_n6182_n2876# a_n6182_n3152# 0.0316f
C754 delay_offset a_n6207_n1211# 0.00113f
C755 ready x2.x10.Y 0.0967f
C756 x4.x9.output_stack x4.x6.floating 0.228f
C757 a_n6182_1664# x4.x9.output_stack 0.032f
C758 a_n397_736# a_1094_824# 4.29e-20
C759 a_n6182_1664# x4.x6.floating 0.0161f
C760 a_1499_824# a_1158_1098# 0.00118f
C761 a_1094_1190# a_618_824# 0.00133f
C762 a_n6207_689# x4.x9.output_stack 0.00227f
C763 x9.A x2.x10.Y 1.13e-19
C764 x2.x3[1].floating x2.x9.output_stack 0.341f
C765 x2.x7.floating a_n6135_n1349# 0.00959f
C766 ready a_n6295_n1763# 0.0217f
C767 async_clk_sar a_1913_1909# 3.56e-20
C768 a_944_1775# a_1159_798# 1.36e-19
C769 async_clk_sar sample_clk 3.03e-19
C770 a_n6135_n139# a_n6207_n139# 0.00227f
C771 x4.x6.SW async_resetb_delay_ctrl_code[0] 4.27e-21
C772 async_setb_delay_ctrl_code[1] a_n397_n1948# 3.4e-20
C773 a_n6295_275# x4.x7.floating 0.00409f
C774 a_n6135_413# x4.x4[3].floating 8.29e-19
C775 a_n6135_137# x4.x6.SW 1.28e-19
C776 a_210_798# a_305_798# 0.0968f
C777 delay_offset async_resetb_delay_ctrl_code[0] 0.0034f
C778 x2.x6.floating x2.x9.output_stack 0.229f
C779 ready async_resetb_delay_ctrl_code[2] 1.35e-19
C780 a_n397_736# a_860_798# 2.1e-19
C781 a_n6295_275# async_resetb_delay_ctrl_code[2] 6.81e-20
C782 x10.Y a_305_798# 0.124f
C783 a_n6135_137# delay_offset 0.00347f
C784 async_setb_delay_ctrl_code[2] x2.x10.Y 0.00203f
C785 a_1296_1190# a_1158_1098# 1.09e-19
C786 x27.Q_N x10.A 1.38e-19
C787 x4.x2.floating x27.Q_N 2.07e-19
C788 sample_clk a_1158_1098# 0.0125f
C789 a_1771_1775# a_1159_798# 3.71e-19
C790 vdd a_n397_1077# 0.26f
C791 a_n6182_n3152# x2.x9.output_stack 1.5e-19
C792 x2.x6.SW async_resetb_delay_ctrl_code[0] 3.98e-21
C793 x2.x4[3].floating async_resetb_delay_ctrl_code[0] 7.6e-20
C794 ready a_n6270_n2738# 0.0175f
C795 eob x4.x5[7].floating 2.39e-19
C796 sample_clk a_1307_1909# 7.17e-20
C797 x4.x3[1].floating async_resetb_delay_ctrl_code[2] 0.00115f
C798 x4.x10.Y a_n397_1077# 0.00127f
C799 async_clk_sar x4.x9.output_stack 0.415f
C800 async_setb_delay_ctrl_code[2] a_n6295_n1763# 3.81e-20
C801 x9.Y a_n397_1077# 8.69e-20
C802 async_clk_sar x4.x6.floating 0.144f
C803 x3.A0 a_860_798# 8.92e-19
C804 async_clk_sar a_n6182_1664# 0.0523f
C805 x2.x6.floating a_n6182_n3152# 0.0191f
C806 async_setb_delay_ctrl_code[2] x4.x7.floating 1.63e-20
C807 a_n6295_n1487# a_n6207_n1349# 0.00227f
C808 x3.A0 a_1631_1008# 1.39e-19
C809 async_clk_sar a_n6295_n277# 0.0127f
C810 async_clk_sar a_n6207_689# 0.00196f
C811 async_setb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[2] 1.86e-19
C812 a_n6295_551# x4.x4[3].floating 1.17e-19
C813 a_n6270_n3014# a_n6270_n3290# 0.0316f
C814 a_n6135_137# a_n6207_137# 0.00227f
C815 delay_offset a_n6295_n1487# 0.0159f
C816 a_2200_1841# a_1159_798# 5.3e-20
C817 a_1086_1909# x4.x5[7].floating 9.13e-22
C818 sample_clk a_1913_1582# 0.00748f
C819 eob a_1403_1582# 0.00575f
C820 a_1771_1775# a_2230_1582# 6.64e-19
C821 vdd async_resetb_delay_ctrl_code[0] 0.00353f
C822 async_setb_delay_ctrl_code[1] delay_offset 0.00333f
C823 a_724_824# a_618_824# 0.0552f
C824 a_n6135_413# x4.x9.output_stack 0.032f
C825 vdd a_n6135_137# 5.05e-19
C826 eob a_618_824# 0.0172f
C827 x4.x10.Y async_resetb_delay_ctrl_code[0] 0.0125f
C828 sample_clk a_305_798# 1.41e-20
C829 a_n6135_413# x4.x6.floating 0.00278f
C830 x2.x4[3].floating a_n6295_n1487# 1.17e-19
C831 x2.x7.floating a_n6207_n1349# 8.52e-19
C832 x2.x6.SW a_n6295_n1487# 8.11e-20
C833 ready a_n6207_n1763# 0.00196f
C834 a_n397_1077# a_210_798# 8.53e-19
C835 a_n6295_n277# a_n6207_n277# 0.0022f
C836 async_setb_delay_ctrl_code[1] x2.x6.SW 7.41e-21
C837 async_setb_delay_ctrl_code[1] x2.x4[3].floating 0.0302f
C838 a_n6207_275# x4.x7.floating 8.52e-19
C839 a_n397_736# a_1298_824# 9.03e-20
C840 a_n397_1077# x10.Y 0.00406f
C841 a_1875_1190# sample_clk 5.07e-19
C842 a_1577_1106# eob 0.00194f
C843 x2.x3[1].floating x2.x2.floating 1.17f
C844 x2.x2.floating x2.x9.output_stack 0.193f
C845 x2.x7.floating delay_offset 0.178f
C846 a_1875_824# a_1158_1098# 0.0019f
C847 a_n6207_275# async_resetb_delay_ctrl_code[2] 2.57e-19
C848 async_setb_delay_ctrl_code[0] x4.x5[7].floating 1.38e-20
C849 a_860_798# x27.Q_N 9.58e-21
C850 eob a_1159_798# 0.0371f
C851 a_n397_736# vdd 0.235f
C852 ready a_n6270_n3014# 0.00866f
C853 x2.x7.floating x2.x6.SW 9.72e-19
C854 x2.x7.floating x2.x4[3].floating 1.18f
C855 a_944_1775# x3.X 0.0612f
C856 a_618_824# x4.x5[7].floating 2.21e-19
C857 x4.x9.output_stack a_305_798# 2.98e-20
C858 async_setb_delay_ctrl_code[2] a_n6207_n1763# 1.08e-19
C859 delay_offset a_n6295_n935# 0.0149f
C860 a_n6295_551# x4.x9.output_stack 0.0388f
C861 a_n397_736# x9.Y 0.00224f
C862 vdd a_n6295_n1487# 0.00308f
C863 async_clk_sar a_1307_1909# 1.2e-19
C864 a_n6295_n1487# a_n6135_n1625# 0.0388f
C865 async_clk_sar a_n6207_n277# 1.34e-19
C866 async_setb_delay_ctrl_code[1] vdd 0.0184f
C867 a_1771_1775# a_1363_798# 5.2e-19
C868 async_clk_sar a_n6135_413# 0.0135f
C869 ready a_n6207_n797# 1.34e-19
C870 a_n6295_551# a_n6207_689# 0.00227f
C871 delay_offset x2.x5[7].floating 0.00308f
C872 vdd x3.A0 1.04f
C873 a_2077_824# a_2200_1841# 3.88e-20
C874 async_resetb_delay_ctrl_code[0] x10.Y 8.99e-21
C875 x2.x4[3].floating a_n6295_n935# 7.17e-20
C876 x3.X a_1771_1775# 0.0804f
C877 x2.x6.SW a_n6295_n935# 3.1e-20
C878 x3.A0 x4.x10.Y 1.39e-19
C879 async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[0] 2.53f
C880 a_n6295_n1# a_n6207_n1# 0.00227f
C881 delay_offset a_n6207_n1487# 0.0014f
C882 x3.A0 x9.Y 8.48e-19
C883 a_1296_1190# a_n397_1077# 1.73e-20
C884 x2.x6.SW x2.x5[7].floating 0.00138f
C885 x2.x4[3].floating x2.x5[7].floating 1.55f
C886 a_n6270_1526# x4.x5[7].floating 2.76e-19
C887 eob a_2230_1582# 1.87e-19
C888 x2.x7.floating vdd 0.0321f
C889 a_n6182_1940# delay_offset 8.71e-20
C890 x2.x7.floating a_n6135_n1625# 0.00959f
C891 async_resetb_delay_ctrl_code[0] x4.x4[3].floating 8.48e-20
C892 a_n397_736# a_210_798# 0.00115f
C893 a_n6135_137# x4.x4[3].floating 8.29e-19
C894 a_n6295_n1# x4.x7.floating 0.00409f
C895 async_clk_sar a_305_798# 5.39e-20
C896 async_setb_delay_ctrl_code[2] a_n6207_n797# 0.00134f
C897 a_n397_736# x10.Y 0.00359f
C898 x4.x3[1].floating x4.x5[7].floating 0.8f
C899 a_2077_824# eob 0.00229f
C900 a_1373_1841# x3.A0 0.0596f
C901 a_n397_736# async_resetb_delay_ctrl_code[1] 3.4e-20
C902 x3.X a_2200_1841# 1.65e-19
C903 a_n6295_n1# async_resetb_delay_ctrl_code[2] 1.46e-19
C904 a_1577_1106# a_618_824# 1.21e-20
C905 a_n6295_551# async_clk_sar 0.0217f
C906 vdd a_n6295_n935# 0.00308f
C907 x4.x9.output_stack a_n397_1077# 0.00887f
C908 async_setb_delay_ctrl_code[0] ready 2.74e-19
C909 vdd x2.x5[7].floating 44f
C910 x3.A0 a_210_798# 0.0792f
C911 ready a_n6270_n3290# 0.00832f
C912 a_618_824# a_1159_798# 0.125f
C913 a_1158_1098# a_305_798# 0.0264f
C914 vdd x27.Q_N 0.0764f
C915 x3.A0 x10.Y 0.175f
C916 x4.x10.Y x27.Q_N 9.42e-21
C917 async_setb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[1] 2.09e-19
C918 async_setb_delay_ctrl_code[0] x9.A 4.05e-19
C919 a_n6207_n1# delay_offset 0.00105f
C920 async_setb_delay_ctrl_code[0] x4.x3[1].floating 3.8e-20
C921 a_944_1775# a_860_798# 1.88e-20
C922 x2.x5[7].floating x9.Y 0.0011f
C923 delay_offset x2.x10.Y 0.0402f
C924 x9.Y x27.Q_N 0.00118f
C925 a_1577_1106# a_1159_798# 0.00276f
C926 a_n6207_n1487# a_n6135_n1625# 0.00227f
C927 a_1875_1190# a_1158_1098# 4.45e-20
C928 ready a_n6135_n1073# 0.0135f
C929 a_818_1106# vdd 0.00622f
C930 async_clk_sar a_n6207_413# 7.93e-19
C931 eob a_1363_798# 0.0222f
C932 a_n6295_551# a_n6135_413# 0.0388f
C933 vdd a_n6182_1940# 0.127f
C934 x3.X a_2134_1909# 2.69e-19
C935 eob x3.X 0.0522f
C936 a_n6182_1940# x4.x10.Y 1.49e-19
C937 x2.x4[3].floating x2.x10.Y 0.00668f
C938 x2.x6.SW x2.x10.Y 0.788f
C939 x4.x6.SW x4.x7.floating 9.72e-19
C940 async_setb_delay_ctrl_code[1] x4.x4[3].floating 7.03e-20
C941 x2.x7.floating async_resetb_delay_ctrl_code[1] 1.76e-20
C942 delay_offset a_n6295_n1763# 0.0311f
C943 async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[0] 4.04e-19
C944 a_1094_1190# a_860_798# 0.00976f
C945 x2.x5[7].floating a_n397_n2289# 0.0132f
C946 a_724_824# x10.A 3.38e-20
C947 x4.x2.floating a_724_824# 3.86e-19
C948 delay_offset x4.x7.floating 0.178f
C949 x4.x9.output_stack async_resetb_delay_ctrl_code[0] 0.0322f
C950 x4.x6.SW async_resetb_delay_ctrl_code[2] 9.9e-21
C951 eob x10.A 1.26e-19
C952 async_resetb_delay_ctrl_code[0] x4.x6.floating 1.49e-19
C953 a_n6135_137# x4.x9.output_stack 1.74e-19
C954 a_n6182_1940# a_n6270_1802# 0.0704f
C955 a_1771_1775# a_1631_1008# 4.17e-20
C956 a_n6135_137# x4.x6.floating 0.00167f
C957 x2.x3[1].floating async_resetb_delay_ctrl_code[0] 3.8e-20
C958 async_resetb_delay_ctrl_code[0] x2.x9.output_stack 2.59e-20
C959 delay_offset async_resetb_delay_ctrl_code[2] 0.0282f
C960 x2.x6.SW a_n6295_n1763# 0.00179f
C961 x2.x4[3].floating a_n6295_n1763# 1.17e-19
C962 x2.x7.floating a_n6207_n1625# 8.52e-19
C963 a_n6295_n277# async_resetb_delay_ctrl_code[0] 4.51e-19
C964 async_clk_sar a_n397_1077# 0.00279f
C965 a_n6295_n1# a_n6135_n139# 0.0388f
C966 a_n6135_413# a_n6207_413# 0.00227f
C967 x27.Q_N a_210_798# 0.178f
C968 async_resetb_delay_ctrl_code[1] a_n6295_n935# 1.41e-20
C969 a_n6270_2078# a_n6182_1940# 0.0704f
C970 delay_offset a_n6270_n2738# 0.00273f
C971 a_1296_1190# x3.A0 5.98e-19
C972 x2.x6.floating async_resetb_delay_ctrl_code[0] 1.3e-21
C973 x3.A0 a_1913_1909# 0.00118f
C974 x2.x4[3].floating async_resetb_delay_ctrl_code[2] 3.3e-20
C975 x3.X a_1086_1909# 6.16e-19
C976 sample_clk x3.A0 0.0622f
C977 x27.Q_N x10.Y 0.0348f
C978 a_2077_824# a_618_824# 3.79e-20
C979 a_n6135_n1073# a_n6207_n1073# 0.00227f
C980 a_n6270_n3290# vss 0.0953f
C981 a_n6182_n3152# vss 0.032f
C982 a_n6270_n3014# vss 0.0815f
C983 a_n6182_n2876# vss 0.0402f
C984 a_n6270_n2738# vss 0.0147f
C985 a_n397_n2289# vss 0.276f
C986 x2.x5[7].floating vss 0.107p
C987 x2.x10.Y vss 2.77f
C988 x2.x6.floating vss 0.357f
C989 x2.x6.SW vss 0.299f
C990 x9.A vss 0.631f
C991 x2.x2.floating vss 6.43f
C992 x2.x3[1].floating vss 10.9f
C993 x2.x4[3].floating vss 21.7f
C994 x2.x7.floating vss 5.9f
C995 a_n397_n1948# vss 0.306f
C996 async_setb_delay_ctrl_code[0] vss 6.82f
C997 async_setb_delay_ctrl_code[1] vss 3.78f
C998 async_setb_delay_ctrl_code[2] vss 2.38f
C999 x2.x9.output_stack vss 1.52f
C1000 a_n6207_n1763# vss 6.32e-19
C1001 a_n6207_n1625# vss 6.69e-19
C1002 a_n6295_n1763# vss 0.118f
C1003 a_n6135_n1625# vss 0.111f
C1004 a_n6207_n1487# vss 7.1e-19
C1005 a_n6207_n1349# vss 7.57e-19
C1006 a_n6295_n1487# vss 0.113f
C1007 a_n6135_n1349# vss 0.114f
C1008 a_n6207_n1211# vss 8.09e-19
C1009 a_n6207_n1073# vss 8.65e-19
C1010 a_n6295_n1211# vss 0.113f
C1011 a_n6135_n1073# vss 0.164f
C1012 a_n6207_n935# vss 9.21e-19
C1013 a_n6207_n797# vss 0.00426f
C1014 a_n6295_n935# vss 0.169f
C1015 ready vss 1.43f
C1016 a_n6207_n277# vss 0.00426f
C1017 a_n6207_n139# vss 9.21e-19
C1018 a_n6295_n277# vss 0.169f
C1019 a_n6135_n139# vss 0.164f
C1020 a_n6207_n1# vss 8.65e-19
C1021 a_n6207_137# vss 8.09e-19
C1022 a_n6295_n1# vss 0.113f
C1023 a_n6135_137# vss 0.114f
C1024 a_n6207_275# vss 7.57e-19
C1025 a_n6207_413# vss 7.1e-19
C1026 a_n6295_275# vss 0.113f
C1027 a_n6135_413# vss 0.111f
C1028 a_n6207_551# vss 6.69e-19
C1029 a_n6207_689# vss 6.32e-19
C1030 a_n6295_551# vss 0.118f
C1031 a_1875_824# vss 0.00317f
C1032 a_1499_824# vss 0.189f
C1033 a_1298_824# vss 0.0132f
C1034 a_1094_824# vss 0.00216f
C1035 a_2077_824# vss 0.114f
C1036 a_1875_1190# vss 0.00179f
C1037 a_1577_1106# vss 7.71e-19
C1038 a_724_824# vss 0.165f
C1039 a_1296_1190# vss 0.00487f
C1040 a_1094_1190# vss 4.93e-19
C1041 a_818_1106# vss 7.73e-19
C1042 a_n397_736# vss 0.294f
C1043 x4.x2.floating vss 6.43f
C1044 x4.x3[1].floating vss 10.9f
C1045 x4.x4[3].floating vss 21.7f
C1046 x4.x7.floating vss 5.9f
C1047 async_resetb_delay_ctrl_code[0] vss 6.82f
C1048 async_resetb_delay_ctrl_code[1] vss 3.78f
C1049 async_resetb_delay_ctrl_code[2] vss 2.38f
C1050 x27.Q_N vss 0.103f
C1051 a_1631_1008# vss 0.285f
C1052 a_1363_798# vss 0.294f
C1053 a_1159_798# vss 0.603f
C1054 a_1158_1098# vss 0.579f
C1055 x9.Y vss 2.5f
C1056 a_860_798# vss 0.256f
C1057 a_618_824# vss 0.393f
C1058 a_305_798# vss 0.464f
C1059 x10.Y vss 0.441f
C1060 x4.x5[7].floating vss 0.107p
C1061 x4.x6.floating vss 0.358f
C1062 a_210_798# vss 0.225f
C1063 x10.A vss 0.598f
C1064 a_n397_1077# vss 0.254f
C1065 a_2230_1582# vss 0.00141f
C1066 a_1913_1582# vss 0.00174f
C1067 a_1403_1582# vss 6.56e-19
C1068 a_1086_1582# vss 6.98e-19
C1069 a_2134_1909# vss 0.0105f
C1070 a_1913_1909# vss 0.00474f
C1071 x4.x9.output_stack vss 1.51f
C1072 x4.x6.SW vss 0.299f
C1073 x4.x10.Y vss 2.76f
C1074 delay_offset vss 3.34f
C1075 a_n6270_1526# vss 0.0147f
C1076 a_1307_1909# vss 0.00815f
C1077 a_1086_1909# vss 0.00388f
C1078 a_n6182_1664# vss 0.0402f
C1079 a_2200_1841# vss 0.485f
C1080 x3.A0 vss 0.967f
C1081 sample_clk vss 1.19f
C1082 a_1771_1775# vss 0.487f
C1083 a_1373_1841# vss 0.39f
C1084 x3.X vss 0.835f
C1085 eob vss 0.738f
C1086 a_944_1775# vss 0.493f
C1087 a_n6270_1802# vss 0.0815f
C1088 a_n6182_1940# vss 0.032f
C1089 a_n6270_2078# vss 0.0953f
C1090 async_clk_sar vss 2.89f
C1091 vdd vss 87.9f
C1092 async_resetb_delay_ctrl_code[0].t0 vss 0.0553f
C1093 async_setb_delay_ctrl_code[1].t1 vss 0.0273f
C1094 async_setb_delay_ctrl_code[1].t0 vss 0.0273f
C1095 async_setb_delay_ctrl_code[1].n0 vss 0.666f
C1096 x2.x5[7].floating.n0 vss -7.99f
C1097 x2.x5[7].floating.n1 vss -28.9f
C1098 x2.x5[7].floating.n2 vss 3.83f
C1099 x2.x5[7].floating.n3 vss -7.07f
C1100 x2.x5[7].floating.n4 vss -28.3f
C1101 x2.x5[7].floating.n5 vss 52.7f
C1102 x2.x5[7].floating.n6 vss 2.47f
C1103 x2.x5[7].floating.n7 vss 0.766f
C1104 x2.x5[7].floating.n8 vss -33f
C1105 x2.x5[7].floating.n9 vss -5.01f
C1106 x2.x5[7].floating.n10 vss 3.83f
C1107 x2.x5[7].floating.n11 vss -28.9f
C1108 x2.x5[7].floating.n12 vss -7.84f
C1109 x2.x5[7].floating.n13 vss 3.23f
C1110 x2.x5[7].floating.n14 vss 52f
C1111 x2.x5[7].floating.n15 vss 2.68f
C1112 x2.x5[7].floating.n16 vss -7.07f
C1113 x2.x5[7].floating.n17 vss -28.9f
C1114 x2.x5[7].floating.n18 vss 3.83f
C1115 x2.x5[7].floating.n19 vss -4.56f
C1116 x2.x5[7].floating.n20 vss -33.5f
C1117 x2.x5[7].floating.n21 vss 0.766f
C1118 x2.x5[7].floating.n22 vss 2.47f
C1119 x2.x5[7].floating.n23 vss 51.5f
C1120 x2.x5[7].floating.n24 vss 2.47f
C1121 x2.x5[7].floating.n25 vss 0.766f
C1122 x2.x5[7].floating.n26 vss -33f
C1123 x2.x5[7].floating.n27 vss -5.01f
C1124 x2.x5[7].floating.n28 vss 3.83f
C1125 x2.x5[7].floating.n29 vss -28.9f
C1126 x2.x5[7].floating.n30 vss -7.84f
C1127 x2.x5[7].floating.n31 vss 3.23f
C1128 x2.x5[7].floating.n32 vss 52f
C1129 x2.x5[7].floating.n33 vss 2.68f
C1130 x2.x5[7].floating.n34 vss -7.07f
C1131 x2.x5[7].floating.n35 vss -28.9f
C1132 x2.x5[7].floating.n36 vss 3.83f
C1133 x2.x5[7].floating.n37 vss -4.56f
C1134 x2.x5[7].floating.n38 vss -33.5f
C1135 x2.x5[7].floating.n39 vss 0.766f
C1136 x2.x5[7].floating.n40 vss 2.47f
C1137 x2.x5[7].floating.n41 vss 51.5f
C1138 x2.x5[7].floating.n42 vss 2.47f
C1139 x2.x5[7].floating.n43 vss 0.766f
C1140 x2.x5[7].floating.n44 vss -41.6f
C1141 x2.x5[7].floating.n45 vss -15.2f
C1142 x2.x5[7].floating.n46 vss -15.2f
C1143 x2.x5[7].floating.n47 vss 1.17f
C1144 x2.x5[7].floating.t0 vss 0.859f
C1145 x2.x5[7].floating.n48 vss 6.5f
C1146 x2.x5[7].floating.n49 vss 1.36f
C1147 x2.x5[7].floating.n50 vss 2.19f
C1148 x2.x5[7].floating.n51 vss 1.06f
C1149 x2.x5[7].floating.n52 vss 0.367f
C1150 x2.x5[7].floating.n53 vss 1.06f
C1151 x2.x5[7].floating.n54 vss 2.79f
C1152 x2.x5[7].floating.n55 vss 51.4f
C1153 x2.x5[7].floating.n56 vss 2.8f
C1154 x2.x5[7].floating.n57 vss 1.06f
C1155 x2.x5[7].floating.n58 vss 0.364f
C1156 x2.x5[7].floating.n59 vss 1.21f
C1157 x2.x5[7].floating.t4 vss 0.859f
C1158 x2.x5[7].floating.n60 vss 6.67f
C1159 x2.x5[7].floating.n61 vss 1.15f
C1160 x2.x5[7].floating.n62 vss 2.17f
C1161 x2.x5[7].floating.n63 vss 1.06f
C1162 x2.x5[7].floating.n64 vss 2.22f
C1163 x2.x5[7].floating.n65 vss -8.01f
C1164 x2.x5[7].floating.n66 vss -28.9f
C1165 x2.x5[7].floating.n67 vss 3.83f
C1166 x2.x5[7].floating.n68 vss -7.07f
C1167 x2.x5[7].floating.n69 vss -28.3f
C1168 x2.x5[7].floating.n70 vss 52.7f
C1169 x2.x5[7].floating.n71 vss -28.3f
C1170 x2.x5[7].floating.n72 vss -7.07f
C1171 x2.x5[7].floating.n73 vss 3.83f
C1172 x2.x5[7].floating.n74 vss -28.9f
C1173 x2.x5[7].floating.n75 vss -7.99f
C1174 x2.x5[7].floating.n76 vss 2.22f
C1175 x2.x5[7].floating.n77 vss 1.17f
C1176 x2.x5[7].floating.t2 vss 0.859f
C1177 x2.x5[7].floating.n78 vss 6.5f
C1178 x2.x5[7].floating.n79 vss 1.36f
C1179 x2.x5[7].floating.n80 vss 2.19f
C1180 x2.x5[7].floating.n81 vss 1.06f
C1181 x2.x5[7].floating.n82 vss 0.367f
C1182 x2.x5[7].floating.n83 vss 1.06f
C1183 x2.x5[7].floating.n84 vss 2.79f
C1184 x2.x5[7].floating.n85 vss 51.4f
C1185 x2.x5[7].floating.n86 vss 2.8f
C1186 x2.x5[7].floating.n87 vss 1.06f
C1187 x2.x5[7].floating.n88 vss 0.364f
C1188 x2.x5[7].floating.n89 vss 1.21f
C1189 x2.x5[7].floating.t5 vss 0.859f
C1190 x2.x5[7].floating.n90 vss 6.67f
C1191 x2.x5[7].floating.n91 vss 1.15f
C1192 x2.x5[7].floating.n92 vss 2.17f
C1193 x2.x5[7].floating.n93 vss 1.06f
C1194 x2.x5[7].floating.n94 vss 2.22f
C1195 x2.x5[7].floating.n95 vss -8.01f
C1196 x2.x5[7].floating.n96 vss -28.9f
C1197 x2.x5[7].floating.n97 vss 3.83f
C1198 x2.x5[7].floating.n98 vss -7.07f
C1199 x2.x5[7].floating.n99 vss -28.3f
C1200 x2.x5[7].floating.n100 vss 52.7f
C1201 x2.x5[7].floating.n101 vss -28.3f
C1202 x2.x5[7].floating.n102 vss -7.07f
C1203 x2.x5[7].floating.n103 vss 3.83f
C1204 x2.x5[7].floating.n104 vss -28.9f
C1205 x2.x5[7].floating.n105 vss -7.99f
C1206 x2.x5[7].floating.n106 vss 2.22f
C1207 x2.x5[7].floating.n107 vss 1.17f
C1208 x2.x5[7].floating.t3 vss 0.859f
C1209 x2.x5[7].floating.n108 vss 6.5f
C1210 x2.x5[7].floating.n109 vss 1.36f
C1211 x2.x5[7].floating.n110 vss 2.19f
C1212 x2.x5[7].floating.n111 vss 1.06f
C1213 x2.x5[7].floating.n112 vss 0.367f
C1214 x2.x5[7].floating.n113 vss 1.06f
C1215 x2.x5[7].floating.n114 vss 2.79f
C1216 x2.x5[7].floating.n115 vss -28.3f
C1217 x2.x5[7].floating.n116 vss -7.07f
C1218 x2.x5[7].floating.n117 vss 3.83f
C1219 x2.x5[7].floating.n118 vss -28.9f
C1220 x2.x5[7].floating.n119 vss -8.01f
C1221 x2.x5[7].floating.n120 vss 2.22f
C1222 x2.x5[7].floating.n121 vss 1.21f
C1223 x2.x5[7].floating.t6 vss 0.859f
C1224 x2.x5[7].floating.n122 vss 6.67f
C1225 x2.x5[7].floating.n123 vss 1.15f
C1226 x2.x5[7].floating.n124 vss 2.17f
C1227 x2.x5[7].floating.n125 vss 1.06f
C1228 x2.x5[7].floating.n126 vss 0.364f
C1229 x2.x5[7].floating.n127 vss 1.06f
C1230 x2.x5[7].floating.n128 vss 2.8f
C1231 x2.x5[7].floating.n129 vss 51.4f
C1232 x2.x5[7].floating.n130 vss 51.5f
C1233 x2.x5[7].floating.n131 vss 2.47f
C1234 x2.x5[7].floating.n132 vss 0.766f
C1235 x2.x5[7].floating.n133 vss -33.5f
C1236 x2.x5[7].floating.n134 vss -4.56f
C1237 x2.x5[7].floating.n135 vss 3.83f
C1238 x2.x5[7].floating.n136 vss -28.9f
C1239 x2.x5[7].floating.n137 vss -7.07f
C1240 x2.x5[7].floating.n138 vss 2.68f
C1241 x2.x5[7].floating.n139 vss 52f
C1242 x2.x5[7].floating.n140 vss 3.23f
C1243 x2.x5[7].floating.n141 vss 2.22f
C1244 x2.x5[7].floating.n142 vss 1.17f
C1245 x2.x5[7].floating.t1 vss 0.859f
C1246 x2.x5[7].floating.n143 vss 6.5f
C1247 x2.x5[7].floating.n144 vss 1.36f
C1248 x2.x5[7].floating.n145 vss 2.19f
C1249 x2.x5[7].floating.n146 vss 1.06f
C1250 x2.x5[7].floating.n147 vss 0.367f
C1251 x2.x5[7].floating.n148 vss 1.06f
C1252 x2.x5[7].floating.n149 vss 2.79f
C1253 x2.x5[7].floating.n150 vss 51.4f
C1254 x2.x5[7].floating.n151 vss 2.8f
C1255 x2.x5[7].floating.n152 vss 1.06f
C1256 x2.x5[7].floating.n153 vss 0.364f
C1257 x2.x5[7].floating.n154 vss 1.21f
C1258 x2.x5[7].floating.t7 vss 0.859f
C1259 x2.x5[7].floating.n155 vss 6.67f
C1260 x2.x5[7].floating.n156 vss 1.15f
C1261 x2.x5[7].floating.n157 vss 2.17f
C1262 x2.x5[7].floating.n158 vss 1.06f
C1263 x2.x5[7].floating.n159 vss -17.4f
C1264 x2.x5[7].floating.n160 vss -17.2f
C1265 x2.x5[7].floating.n161 vss -43.6f
C1266 x2.x5[7].floating.n162 vss 0.766f
C1267 x2.x5[7].floating.n163 vss 2.47f
C1268 x2.x5[7].floating.n164 vss 51.5f
C1269 x2.x5[7].floating.n165 vss 2.47f
C1270 x2.x5[7].floating.n166 vss 0.766f
C1271 x2.x5[7].floating.n167 vss -33f
C1272 x2.x5[7].floating.n168 vss -5.01f
C1273 x2.x5[7].floating.n169 vss 3.83f
C1274 x2.x5[7].floating.n170 vss -28.9f
C1275 x2.x5[7].floating.n171 vss -7.84f
C1276 x2.x10.Y.t1 vss 0.0526f
C1277 x2.x10.Y.n0 vss 0.0169f
C1278 x2.x10.Y.t9 vss 0.0167f
C1279 x2.x10.Y.t5 vss 0.0167f
C1280 x2.x10.Y.t7 vss 0.0167f
C1281 x2.x10.Y.t4 vss 0.0167f
C1282 x2.x10.Y.t6 vss 0.0167f
C1283 x2.x10.Y.t3 vss 0.0167f
C1284 x2.x10.Y.t8 vss 0.0167f
C1285 x2.x10.Y.t2 vss 0.0167f
C1286 x2.x10.Y.n1 vss 0.221f
C1287 x2.x10.Y.n2 vss 0.0366f
C1288 x2.x10.Y.t0 vss 0.0174f
C1289 x2.x10.Y.n3 vss 0.0188f
C1290 x2.x10.Y.n4 vss 0.0189f
C1291 x2.x10.Y.n5 vss 0.00592f
C1292 async_setb_delay_ctrl_code[0].t0 vss 0.0553f
C1293 async_clk_sar.t0 vss 0.0202f
C1294 async_clk_sar.t1 vss 0.0171f
C1295 async_clk_sar.n0 vss 0.0489f
C1296 async_clk_sar.n1 vss 0.0144f
C1297 async_clk_sar.n2 vss 0.0427f
C1298 async_clk_sar.n3 vss 0.833f
C1299 async_clk_sar.t3 vss 0.0162f
C1300 async_clk_sar.t9 vss 0.0263f
C1301 async_clk_sar.t14 vss 0.0263f
C1302 async_clk_sar.t20 vss 0.0263f
C1303 async_clk_sar.t15 vss 0.0263f
C1304 async_clk_sar.t4 vss 0.0263f
C1305 async_clk_sar.t22 vss 0.0263f
C1306 async_clk_sar.t10 vss 0.0179f
C1307 async_clk_sar.n4 vss 0.0292f
C1308 async_clk_sar.t8 vss 0.0162f
C1309 async_clk_sar.t13 vss 0.0263f
C1310 async_clk_sar.t5 vss 0.0263f
C1311 async_clk_sar.t17 vss 0.0263f
C1312 async_clk_sar.t11 vss 0.0263f
C1313 async_clk_sar.t23 vss 0.0263f
C1314 async_clk_sar.t19 vss 0.0263f
C1315 async_clk_sar.t6 vss 0.0178f
C1316 async_clk_sar.n5 vss 0.00542f
C1317 async_clk_sar.n6 vss 0.00813f
C1318 async_clk_sar.n7 vss 0.00794f
C1319 async_clk_sar.n8 vss 0.0187f
C1320 async_clk_sar.n9 vss 1.35f
C1321 async_clk_sar.n10 vss 0.16f
C1322 async_clk_sar.n11 vss 0.00703f
C1323 async_clk_sar.t18 vss 0.0154f
C1324 async_clk_sar.t2 vss 0.0263f
C1325 async_clk_sar.t16 vss 0.0263f
C1326 async_clk_sar.t21 vss 0.0263f
C1327 async_clk_sar.t7 vss 0.0263f
C1328 async_clk_sar.t12 vss 0.0251f
C1329 async_clk_sar.n12 vss 0.056f
C1330 async_clk_sar.n13 vss 0.126f
C1331 async_clk_sar.n14 vss 0.858f
C1332 async_resetb_delay_ctrl_code[1].t0 vss 0.0273f
C1333 async_resetb_delay_ctrl_code[1].t1 vss 0.0273f
C1334 async_resetb_delay_ctrl_code[1].n0 vss 0.666f
C1335 vdd.n0 vss 0.0043f
C1336 vdd.n1 vss 0.0192f
C1337 vdd.n2 vss 0.0111f
C1338 vdd.n3 vss 0.0155f
C1339 vdd.n4 vss 0.00731f
C1340 vdd.n5 vss 0.00368f
C1341 vdd.n6 vss 0.00394f
C1342 vdd.n7 vss -0.174f
C1343 vdd.n8 vss 0.007f
C1344 vdd.n9 vss 0.00311f
C1345 vdd.n10 vss 0.00297f
C1346 vdd.n11 vss 0.00241f
C1347 vdd.n12 vss 0.0141f
C1348 vdd.n13 vss 0.00241f
C1349 vdd.n14 vss 0.00271f
C1350 vdd.n15 vss 0.0115f
C1351 vdd.n16 vss 0.00248f
C1352 vdd.n17 vss 0.178f
C1353 vdd.n18 vss 0.00933f
C1354 vdd.n19 vss 2.83e-19
C1355 vdd.n20 vss 0.00821f
C1356 vdd.n21 vss 0.00368f
C1357 vdd.n22 vss 0.00394f
C1358 vdd.n23 vss 0.00851f
C1359 vdd.n24 vss 0.007f
C1360 vdd.n25 vss 0.00311f
C1361 vdd.n26 vss 0.00297f
C1362 vdd.n27 vss 0.00297f
C1363 vdd.n28 vss 0.00241f
C1364 vdd.n29 vss 0.00248f
C1365 vdd.n30 vss 0.219f
C1366 vdd.n31 vss 0.0115f
C1367 vdd.n32 vss 0.00241f
C1368 vdd.n33 vss 0.00241f
C1369 vdd.n34 vss 4.25e-19
C1370 vdd.n35 vss 0.00594f
C1371 vdd.n36 vss 0.00297f
C1372 vdd.n37 vss 0.00722f
C1373 vdd.n38 vss -0.0674f
C1374 vdd.n39 vss 0.00851f
C1375 vdd.n40 vss 0.00437f
C1376 vdd.n41 vss -0.077f
C1377 vdd.n42 vss 2.92e-19
C1378 vdd.n43 vss 4.25e-19
C1379 vdd.n44 vss 0.00524f
C1380 vdd.n45 vss 0.00311f
C1381 vdd.n46 vss 2.83e-19
C1382 vdd.n47 vss 0.00933f
C1383 vdd.n48 vss 0.0472f
C1384 vdd.n49 vss 0.00248f
C1385 vdd.n50 vss 0.00241f
C1386 vdd.n51 vss 0.00241f
C1387 vdd.n52 vss 0.00594f
C1388 vdd.n53 vss 0.00368f
C1389 vdd.n54 vss 0.00394f
C1390 vdd.n55 vss 0.00423f
C1391 vdd.n56 vss 0.007f
C1392 vdd.n57 vss 0.00851f
C1393 vdd.n58 vss 0.007f
C1394 vdd.n59 vss 0.00311f
C1395 vdd.n60 vss 0.00297f
C1396 vdd.n61 vss 0.00241f
C1397 vdd.n62 vss 0.00821f
C1398 vdd.n63 vss 0.00241f
C1399 vdd.n64 vss 0.0115f
C1400 vdd.n65 vss 0.111f
C1401 vdd.n66 vss 0.0211f
C1402 vdd.n67 vss 0.0282f
C1403 vdd.n68 vss 0.00856f
C1404 vdd.n69 vss 0.00368f
C1405 vdd.n70 vss -0.0674f
C1406 vdd.n71 vss 0.00518f
C1407 vdd.n72 vss 0.00394f
C1408 vdd.n73 vss 0.00297f
C1409 vdd.n74 vss 0.00241f
C1410 vdd.n75 vss 4.25e-19
C1411 vdd.n76 vss 0.00241f
C1412 vdd.n77 vss 0.0161f
C1413 vdd.n78 vss 0.0115f
C1414 vdd.n79 vss 0.00248f
C1415 vdd.n80 vss 0.178f
C1416 vdd.n81 vss 0.00933f
C1417 vdd.n82 vss 2.83e-19
C1418 vdd.n83 vss 0.00821f
C1419 vdd.n84 vss 0.00368f
C1420 vdd.n85 vss 0.00394f
C1421 vdd.n86 vss 0.007f
C1422 vdd.n87 vss 0.0082f
C1423 vdd.n88 vss 0.007f
C1424 vdd.n89 vss 0.00311f
C1425 vdd.n90 vss 0.00297f
C1426 vdd.n91 vss 0.00297f
C1427 vdd.n92 vss 0.00241f
C1428 vdd.n93 vss 0.00248f
C1429 vdd.n94 vss 0.219f
C1430 vdd.n95 vss 0.0115f
C1431 vdd.n96 vss 0.00241f
C1432 vdd.n97 vss 0.00241f
C1433 vdd.n98 vss 4.25e-19
C1434 vdd.n99 vss 0.00594f
C1435 vdd.n100 vss 0.00297f
C1436 vdd.n101 vss 0.00722f
C1437 vdd.n102 vss -0.0674f
C1438 vdd.n103 vss 0.0082f
C1439 vdd.n104 vss 0.00437f
C1440 vdd.n105 vss -0.0772f
C1441 vdd.n106 vss 2.92e-19
C1442 vdd.n107 vss 4.25e-19
C1443 vdd.n108 vss 0.00524f
C1444 vdd.n109 vss 0.00311f
C1445 vdd.n110 vss 2.83e-19
C1446 vdd.n111 vss 0.00933f
C1447 vdd.n112 vss 0.0472f
C1448 vdd.n113 vss 0.00248f
C1449 vdd.n114 vss 0.00241f
C1450 vdd.n115 vss 0.00241f
C1451 vdd.n116 vss 0.00594f
C1452 vdd.n117 vss 0.00368f
C1453 vdd.n118 vss 0.00394f
C1454 vdd.n119 vss 0.00423f
C1455 vdd.n120 vss 0.007f
C1456 vdd.n121 vss 0.0082f
C1457 vdd.n122 vss 0.007f
C1458 vdd.n123 vss 0.00311f
C1459 vdd.n124 vss 0.00297f
C1460 vdd.n125 vss 0.00241f
C1461 vdd.n126 vss 0.00821f
C1462 vdd.n127 vss 0.00241f
C1463 vdd.n128 vss 0.0115f
C1464 vdd.n129 vss 0.111f
C1465 vdd.n130 vss 0.0211f
C1466 vdd.n131 vss 2.83e-19
C1467 vdd.n132 vss 0.00821f
C1468 vdd.n133 vss 0.00368f
C1469 vdd.n134 vss -0.0674f
C1470 vdd.n135 vss 0.0294f
C1471 vdd.n136 vss 0.0255f
C1472 vdd.n137 vss 0.00311f
C1473 vdd.n138 vss 0.00297f
C1474 vdd.n139 vss 0.00297f
C1475 vdd.n140 vss 0.00241f
C1476 vdd.n141 vss 0.00241f
C1477 vdd.n142 vss 0.0234f
C1478 vdd.n143 vss 0.00297f
C1479 vdd.n144 vss 0.00437f
C1480 vdd.n145 vss 0.00821f
C1481 vdd.n146 vss 0.00241f
C1482 vdd.n147 vss 0.00248f
C1483 vdd.n148 vss 0.178f
C1484 vdd.n149 vss 0.00933f
C1485 vdd.n150 vss 0.00241f
C1486 vdd.n151 vss 0.00241f
C1487 vdd.n152 vss 0.00311f
C1488 vdd.n153 vss 0.00368f
C1489 vdd.n154 vss 0.00335f
C1490 vdd.n155 vss 2.92e-19
C1491 vdd.n156 vss 0.00518f
C1492 vdd.n157 vss 2.92e-19
C1493 vdd.n158 vss 0.00297f
C1494 vdd.n159 vss 0.00821f
C1495 vdd.n160 vss 0.00877f
C1496 vdd.n161 vss 0.0115f
C1497 vdd.n162 vss 0.0472f
C1498 vdd.n163 vss 0.00248f
C1499 vdd.n164 vss 0.00241f
C1500 vdd.n165 vss 0.00241f
C1501 vdd.n166 vss 0.00821f
C1502 vdd.n167 vss 4.25e-19
C1503 vdd.n168 vss 0.00877f
C1504 vdd.n169 vss 0.00297f
C1505 vdd.n170 vss 0.00368f
C1506 vdd.n171 vss 0.00335f
C1507 vdd.n172 vss -0.0832f
C1508 vdd.n173 vss 0.00423f
C1509 vdd.n174 vss 0.00502f
C1510 vdd.n175 vss 0.00311f
C1511 vdd.n176 vss 0.00241f
C1512 vdd.n177 vss 0.00241f
C1513 vdd.n178 vss 0.00933f
C1514 vdd.n179 vss 0.219f
C1515 vdd.n180 vss 0.0115f
C1516 vdd.n181 vss 0.00877f
C1517 vdd.n182 vss 0.00821f
C1518 vdd.n183 vss 0.00297f
C1519 vdd.n184 vss 2.92e-19
C1520 vdd.n185 vss 0.00335f
C1521 vdd.n186 vss 0.0082f
C1522 vdd.n187 vss 0.00335f
C1523 vdd.n188 vss 0.00311f
C1524 vdd.n189 vss 0.00241f
C1525 vdd.n190 vss 0.00241f
C1526 vdd.n191 vss 0.00311f
C1527 vdd.n192 vss 0.00248f
C1528 vdd.n193 vss 0.178f
C1529 vdd.n194 vss 0.00933f
C1530 vdd.n195 vss 0.00241f
C1531 vdd.n196 vss 0.00241f
C1532 vdd.n197 vss 0.00821f
C1533 vdd.n198 vss 0.00311f
C1534 vdd.n199 vss 0.00368f
C1535 vdd.n200 vss 0.00335f
C1536 vdd.n201 vss 2.92e-19
C1537 vdd.n202 vss -0.0832f
C1538 vdd.n203 vss 2.92e-19
C1539 vdd.n204 vss 0.00297f
C1540 vdd.n205 vss 0.0265f
C1541 vdd.n206 vss 0.0269f
C1542 vdd.n207 vss 0.0166f
C1543 vdd.n208 vss 0.0472f
C1544 vdd.n209 vss 0.00248f
C1545 vdd.n210 vss 0.00241f
C1546 vdd.n211 vss 0.00311f
C1547 vdd.n212 vss 0.0115f
C1548 vdd.n213 vss 0.178f
C1549 vdd.n214 vss 0.00933f
C1550 vdd.n215 vss 2.83e-19
C1551 vdd.n216 vss 0.00594f
C1552 vdd.n217 vss 0.00722f
C1553 vdd.n218 vss 0.00297f
C1554 vdd.n219 vss 0.007f
C1555 vdd.n220 vss 0.00394f
C1556 vdd.n221 vss 0.00518f
C1557 vdd.n222 vss 0.00394f
C1558 vdd.n223 vss 0.00297f
C1559 vdd.n224 vss 0.00241f
C1560 vdd.n225 vss 0.00311f
C1561 vdd.n226 vss 0.007f
C1562 vdd.n227 vss 0.00518f
C1563 vdd.n228 vss -0.0674f
C1564 vdd.n229 vss 0.00368f
C1565 vdd.n230 vss 0.00821f
C1566 vdd.n231 vss 0.00241f
C1567 vdd.n232 vss 0.00248f
C1568 vdd.n233 vss 0.219f
C1569 vdd.n234 vss 0.0115f
C1570 vdd.n235 vss 0.00241f
C1571 vdd.n236 vss 0.00241f
C1572 vdd.n237 vss 0.00311f
C1573 vdd.n238 vss 0.00297f
C1574 vdd.n239 vss 0.007f
C1575 vdd.n240 vss 0.00518f
C1576 vdd.n241 vss 0.00394f
C1577 vdd.n242 vss 0.00368f
C1578 vdd.n243 vss 0.00821f
C1579 vdd.n244 vss 2.83e-19
C1580 vdd.n245 vss 0.00933f
C1581 vdd.n246 vss 0.0472f
C1582 vdd.n247 vss 0.00248f
C1583 vdd.n248 vss 0.00241f
C1584 vdd.n249 vss 0.00241f
C1585 vdd.n250 vss 0.00594f
C1586 vdd.n251 vss 0.00311f
C1587 vdd.n252 vss 0.00722f
C1588 vdd.n253 vss 0.00297f
C1589 vdd.n254 vss 0.007f
C1590 vdd.n255 vss 0.00518f
C1591 vdd.n256 vss 0.00394f
C1592 vdd.n257 vss 0.00297f
C1593 vdd.n258 vss 0.00241f
C1594 vdd.n259 vss 4.25e-19
C1595 vdd.n260 vss 0.00241f
C1596 vdd.n261 vss 0.0115f
C1597 vdd.n262 vss 0.111f
C1598 vdd.n263 vss 0.0211f
C1599 vdd.n264 vss 2.83e-19
C1600 vdd.n265 vss 0.00821f
C1601 vdd.n266 vss 0.00368f
C1602 vdd.n267 vss -0.0674f
C1603 vdd.n268 vss 0.007f
C1604 vdd.n269 vss 0.0294f
C1605 vdd.n270 vss 0.0255f
C1606 vdd.n271 vss 0.00311f
C1607 vdd.n272 vss 0.00297f
C1608 vdd.n273 vss 0.00297f
C1609 vdd.n274 vss 0.00241f
C1610 vdd.n275 vss 0.00241f
C1611 vdd.n276 vss 0.0234f
C1612 vdd.n277 vss 0.00297f
C1613 vdd.n278 vss 0.00437f
C1614 vdd.n279 vss 0.00821f
C1615 vdd.n280 vss 0.00241f
C1616 vdd.n281 vss 0.00248f
C1617 vdd.n282 vss 0.178f
C1618 vdd.n283 vss 0.00933f
C1619 vdd.n284 vss 0.00241f
C1620 vdd.n285 vss 0.00241f
C1621 vdd.n286 vss 0.00311f
C1622 vdd.n287 vss 0.00368f
C1623 vdd.n288 vss 0.00335f
C1624 vdd.n289 vss 2.92e-19
C1625 vdd.n290 vss 0.00518f
C1626 vdd.n291 vss 2.92e-19
C1627 vdd.n292 vss 0.00297f
C1628 vdd.n293 vss 0.00821f
C1629 vdd.n294 vss 0.00877f
C1630 vdd.n295 vss 0.0115f
C1631 vdd.n296 vss 0.0472f
C1632 vdd.n297 vss 0.00248f
C1633 vdd.n298 vss 0.00241f
C1634 vdd.n299 vss 0.00241f
C1635 vdd.n300 vss 0.00821f
C1636 vdd.n301 vss 4.25e-19
C1637 vdd.n302 vss 0.00877f
C1638 vdd.n303 vss 0.00297f
C1639 vdd.n304 vss 0.00368f
C1640 vdd.n305 vss 0.00335f
C1641 vdd.n306 vss -0.0832f
C1642 vdd.n307 vss 0.00423f
C1643 vdd.n308 vss 0.00502f
C1644 vdd.n309 vss 0.00311f
C1645 vdd.n310 vss 0.00241f
C1646 vdd.n311 vss 0.00241f
C1647 vdd.n312 vss 0.00933f
C1648 vdd.n313 vss 0.219f
C1649 vdd.n314 vss 0.0115f
C1650 vdd.n315 vss 0.00877f
C1651 vdd.n316 vss 0.00821f
C1652 vdd.n317 vss 0.00297f
C1653 vdd.n318 vss 2.92e-19
C1654 vdd.n319 vss 0.00335f
C1655 vdd.n320 vss 0.0082f
C1656 vdd.n321 vss 0.00335f
C1657 vdd.n322 vss 0.00311f
C1658 vdd.n323 vss 0.00241f
C1659 vdd.n324 vss 0.00241f
C1660 vdd.n325 vss 0.00311f
C1661 vdd.n326 vss 0.00248f
C1662 vdd.n327 vss 0.178f
C1663 vdd.n328 vss 0.00933f
C1664 vdd.n329 vss 0.00241f
C1665 vdd.n330 vss 0.00241f
C1666 vdd.n331 vss 0.00821f
C1667 vdd.n332 vss 0.00311f
C1668 vdd.n333 vss 0.00368f
C1669 vdd.n334 vss 0.00335f
C1670 vdd.n335 vss 2.92e-19
C1671 vdd.n336 vss -0.0832f
C1672 vdd.n337 vss 2.92e-19
C1673 vdd.n338 vss 0.00297f
C1674 vdd.n339 vss 0.0265f
C1675 vdd.n340 vss 0.0269f
C1676 vdd.n341 vss 0.0166f
C1677 vdd.n342 vss 0.0472f
C1678 vdd.n343 vss 0.00248f
C1679 vdd.n344 vss 0.00241f
C1680 vdd.n345 vss 0.00311f
C1681 vdd.n346 vss 0.0115f
C1682 vdd.n347 vss 0.178f
C1683 vdd.n348 vss 0.00933f
C1684 vdd.n349 vss 2.83e-19
C1685 vdd.n350 vss 0.00594f
C1686 vdd.n351 vss 0.00722f
C1687 vdd.n352 vss 0.00297f
C1688 vdd.n353 vss 0.007f
C1689 vdd.n354 vss 0.00394f
C1690 vdd.n355 vss 0.00518f
C1691 vdd.n356 vss 0.00394f
C1692 vdd.n357 vss 0.00297f
C1693 vdd.n358 vss 0.00241f
C1694 vdd.n359 vss 0.00311f
C1695 vdd.n360 vss 0.007f
C1696 vdd.n361 vss 0.00518f
C1697 vdd.n362 vss -0.0674f
C1698 vdd.n363 vss 0.00368f
C1699 vdd.n364 vss 0.00821f
C1700 vdd.n365 vss 0.00241f
C1701 vdd.n366 vss 0.00248f
C1702 vdd.n367 vss 0.219f
C1703 vdd.n368 vss 0.0115f
C1704 vdd.n369 vss 0.00241f
C1705 vdd.n370 vss 0.00241f
C1706 vdd.n371 vss 0.00311f
C1707 vdd.n372 vss 0.00297f
C1708 vdd.n373 vss 0.007f
C1709 vdd.n374 vss 0.00518f
C1710 vdd.n375 vss 0.00394f
C1711 vdd.n376 vss 0.00368f
C1712 vdd.n377 vss 0.00821f
C1713 vdd.n378 vss 2.83e-19
C1714 vdd.n379 vss 0.00933f
C1715 vdd.n380 vss 0.0472f
C1716 vdd.n381 vss 0.00248f
C1717 vdd.n382 vss 0.00241f
C1718 vdd.n383 vss 0.00241f
C1719 vdd.n384 vss 0.00594f
C1720 vdd.n385 vss 0.00311f
C1721 vdd.n386 vss 0.00722f
C1722 vdd.n387 vss 0.00297f
C1723 vdd.n388 vss 0.007f
C1724 vdd.n389 vss 0.00518f
C1725 vdd.n390 vss 0.00394f
C1726 vdd.n391 vss 0.00297f
C1727 vdd.n392 vss 0.00241f
C1728 vdd.n393 vss 4.25e-19
C1729 vdd.n394 vss 0.00241f
C1730 vdd.n395 vss 0.0115f
C1731 vdd.n396 vss 0.111f
C1732 vdd.n397 vss 0.0211f
C1733 vdd.n398 vss 2.83e-19
C1734 vdd.n399 vss 0.00821f
C1735 vdd.n400 vss 0.00368f
C1736 vdd.n401 vss -0.0674f
C1737 vdd.n402 vss 0.007f
C1738 vdd.n403 vss 0.0294f
C1739 vdd.n404 vss 0.0255f
C1740 vdd.n405 vss 0.00311f
C1741 vdd.n406 vss 0.00297f
C1742 vdd.n407 vss 0.00297f
C1743 vdd.n408 vss 0.00241f
C1744 vdd.n409 vss 0.00241f
C1745 vdd.n410 vss 0.0234f
C1746 vdd.n411 vss 0.00297f
C1747 vdd.n412 vss 0.00437f
C1748 vdd.n413 vss 0.00821f
C1749 vdd.n414 vss 0.00241f
C1750 vdd.n415 vss 0.00248f
C1751 vdd.n416 vss 0.178f
C1752 vdd.n417 vss 0.00933f
C1753 vdd.n418 vss 0.00241f
C1754 vdd.n419 vss 0.00241f
C1755 vdd.n420 vss 0.00311f
C1756 vdd.n421 vss 0.00368f
C1757 vdd.n422 vss 0.00335f
C1758 vdd.n423 vss 2.92e-19
C1759 vdd.n424 vss 0.00518f
C1760 vdd.n425 vss 2.92e-19
C1761 vdd.n426 vss 0.00297f
C1762 vdd.n427 vss 0.00821f
C1763 vdd.n428 vss 0.00877f
C1764 vdd.n429 vss 0.0115f
C1765 vdd.n430 vss 0.0472f
C1766 vdd.n431 vss 0.00248f
C1767 vdd.n432 vss 0.00241f
C1768 vdd.n433 vss 0.00241f
C1769 vdd.n434 vss 0.00821f
C1770 vdd.n435 vss 4.25e-19
C1771 vdd.n436 vss 0.00877f
C1772 vdd.n437 vss 0.00297f
C1773 vdd.n438 vss 0.00368f
C1774 vdd.n439 vss 0.00335f
C1775 vdd.n440 vss -0.0832f
C1776 vdd.n441 vss 0.00423f
C1777 vdd.n442 vss 0.00502f
C1778 vdd.n443 vss 0.00311f
C1779 vdd.n444 vss 0.00241f
C1780 vdd.n445 vss 0.00241f
C1781 vdd.n446 vss 0.00933f
C1782 vdd.n447 vss 0.219f
C1783 vdd.n448 vss 0.0115f
C1784 vdd.n449 vss 0.00877f
C1785 vdd.n450 vss 0.00821f
C1786 vdd.n451 vss 0.00297f
C1787 vdd.n452 vss 2.92e-19
C1788 vdd.n453 vss 0.00335f
C1789 vdd.n454 vss 0.0082f
C1790 vdd.n455 vss 0.00335f
C1791 vdd.n456 vss 0.00311f
C1792 vdd.n457 vss 0.00241f
C1793 vdd.n458 vss 0.00241f
C1794 vdd.n459 vss 0.00311f
C1795 vdd.n460 vss 0.00248f
C1796 vdd.n461 vss 0.178f
C1797 vdd.n462 vss 0.00933f
C1798 vdd.n463 vss 0.00241f
C1799 vdd.n464 vss 0.00241f
C1800 vdd.n465 vss 0.00821f
C1801 vdd.n466 vss 0.00311f
C1802 vdd.n467 vss 0.00368f
C1803 vdd.n468 vss 0.00335f
C1804 vdd.n469 vss 2.92e-19
C1805 vdd.n470 vss -0.0832f
C1806 vdd.n471 vss 2.92e-19
C1807 vdd.n472 vss 0.00297f
C1808 vdd.n473 vss 0.0265f
C1809 vdd.n474 vss 0.0269f
C1810 vdd.n475 vss 0.0166f
C1811 vdd.n476 vss 0.0472f
C1812 vdd.n477 vss 0.00248f
C1813 vdd.n478 vss 0.00241f
C1814 vdd.n479 vss 0.00311f
C1815 vdd.n480 vss 0.0115f
C1816 vdd.n481 vss 0.178f
C1817 vdd.n482 vss 0.00933f
C1818 vdd.n483 vss 2.83e-19
C1819 vdd.n484 vss 0.00594f
C1820 vdd.n485 vss 0.00722f
C1821 vdd.n486 vss 0.00297f
C1822 vdd.n487 vss 0.007f
C1823 vdd.n488 vss 0.00394f
C1824 vdd.n489 vss 0.00518f
C1825 vdd.n490 vss 0.00394f
C1826 vdd.n491 vss 0.00297f
C1827 vdd.n492 vss 0.00241f
C1828 vdd.n493 vss 0.00311f
C1829 vdd.n494 vss 0.007f
C1830 vdd.n495 vss 0.00518f
C1831 vdd.n496 vss -0.0674f
C1832 vdd.n497 vss 0.00368f
C1833 vdd.n498 vss 0.00821f
C1834 vdd.n499 vss 0.00241f
C1835 vdd.n500 vss 0.00248f
C1836 vdd.n501 vss 0.219f
C1837 vdd.n502 vss 0.0115f
C1838 vdd.n503 vss 0.00241f
C1839 vdd.n504 vss 0.00241f
C1840 vdd.n505 vss 0.00311f
C1841 vdd.n506 vss 0.00297f
C1842 vdd.n507 vss 0.007f
C1843 vdd.n508 vss 0.00518f
C1844 vdd.n509 vss 0.00394f
C1845 vdd.n510 vss 0.00368f
C1846 vdd.n511 vss 0.00821f
C1847 vdd.n512 vss 2.83e-19
C1848 vdd.n513 vss 0.00933f
C1849 vdd.n514 vss 0.0472f
C1850 vdd.n515 vss 0.00248f
C1851 vdd.n516 vss 0.00241f
C1852 vdd.n517 vss 0.00241f
C1853 vdd.n518 vss 0.00594f
C1854 vdd.n519 vss 0.00311f
C1855 vdd.n520 vss 0.00722f
C1856 vdd.n521 vss 0.00297f
C1857 vdd.n522 vss 0.007f
C1858 vdd.n523 vss 0.00518f
C1859 vdd.n524 vss 0.00394f
C1860 vdd.n525 vss 0.00297f
C1861 vdd.n526 vss 0.00241f
C1862 vdd.n527 vss 4.25e-19
C1863 vdd.n528 vss 0.00241f
C1864 vdd.n529 vss 0.0115f
C1865 vdd.n530 vss 0.111f
C1866 vdd.n531 vss 0.0211f
C1867 vdd.n532 vss 2.83e-19
C1868 vdd.n533 vss 0.00821f
C1869 vdd.n534 vss 0.00368f
C1870 vdd.n535 vss -0.0674f
C1871 vdd.n536 vss 0.007f
C1872 vdd.n537 vss 0.0294f
C1873 vdd.n538 vss 0.0255f
C1874 vdd.n539 vss 0.00311f
C1875 vdd.n540 vss 0.00297f
C1876 vdd.n541 vss 0.00297f
C1877 vdd.n542 vss 0.00241f
C1878 vdd.n543 vss 0.00241f
C1879 vdd.n544 vss 0.0234f
C1880 vdd.n545 vss 0.00297f
C1881 vdd.n546 vss 0.00437f
C1882 vdd.n547 vss 0.00821f
C1883 vdd.n548 vss 0.00241f
C1884 vdd.n549 vss 0.00248f
C1885 vdd.n550 vss 0.178f
C1886 vdd.n551 vss 0.00933f
C1887 vdd.n552 vss 0.00241f
C1888 vdd.n553 vss 0.00241f
C1889 vdd.n554 vss 0.00311f
C1890 vdd.n555 vss 0.00368f
C1891 vdd.n556 vss 0.00335f
C1892 vdd.n557 vss 2.92e-19
C1893 vdd.n558 vss 0.00518f
C1894 vdd.n559 vss 2.92e-19
C1895 vdd.n560 vss 0.00297f
C1896 vdd.n561 vss 0.00821f
C1897 vdd.n562 vss 0.00877f
C1898 vdd.n563 vss 0.0115f
C1899 vdd.n564 vss 0.0472f
C1900 vdd.n565 vss 0.00248f
C1901 vdd.n566 vss 0.00241f
C1902 vdd.n567 vss 0.00241f
C1903 vdd.n568 vss 0.00821f
C1904 vdd.n569 vss 4.25e-19
C1905 vdd.n570 vss 0.00877f
C1906 vdd.n571 vss 0.00297f
C1907 vdd.n572 vss 0.00368f
C1908 vdd.n573 vss 0.00335f
C1909 vdd.n574 vss -0.0832f
C1910 vdd.n575 vss 0.00423f
C1911 vdd.n576 vss 0.00502f
C1912 vdd.n577 vss 0.00311f
C1913 vdd.n578 vss 0.00241f
C1914 vdd.n579 vss 0.00241f
C1915 vdd.n580 vss 0.00933f
C1916 vdd.n581 vss 0.219f
C1917 vdd.n582 vss 0.0115f
C1918 vdd.n583 vss 0.00877f
C1919 vdd.n584 vss 0.00821f
C1920 vdd.n585 vss 0.00297f
C1921 vdd.n586 vss 2.92e-19
C1922 vdd.n587 vss 0.00335f
C1923 vdd.n588 vss 0.0082f
C1924 vdd.n589 vss 0.00335f
C1925 vdd.n590 vss 0.00311f
C1926 vdd.n591 vss 0.00241f
C1927 vdd.n592 vss 0.00241f
C1928 vdd.n593 vss 0.00311f
C1929 vdd.n594 vss 0.00248f
C1930 vdd.n595 vss 0.178f
C1931 vdd.n596 vss 0.00933f
C1932 vdd.n597 vss 0.00241f
C1933 vdd.n598 vss 0.00241f
C1934 vdd.n599 vss 0.00821f
C1935 vdd.n600 vss 0.00311f
C1936 vdd.n601 vss 0.00368f
C1937 vdd.n602 vss 0.00335f
C1938 vdd.n603 vss 2.92e-19
C1939 vdd.n604 vss -0.0832f
C1940 vdd.n605 vss 2.92e-19
C1941 vdd.n606 vss 0.00297f
C1942 vdd.n607 vss 0.0349f
C1943 vdd.n608 vss 0.00248f
C1944 vdd.t48 vss 0.514f
C1945 vdd.n609 vss 0.0623f
C1946 vdd.n610 vss 0.00744f
C1947 vdd.n611 vss 0.0179f
C1948 vdd.n612 vss 0.0178f
C1949 vdd.n613 vss 0.00502f
C1950 vdd.n614 vss 0.00394f
C1951 vdd.n615 vss 0.0357f
C1952 vdd.n616 vss 0.0052f
C1953 vdd.n617 vss 0.138f
C1954 vdd.n618 vss 0.0409f
C1955 vdd.n619 vss 0.0178f
C1956 vdd.n620 vss 0.00568f
C1957 vdd.n621 vss 0.00744f
C1958 vdd.n622 vss 0.0728f
C1959 vdd.n623 vss 0.00733f
C1960 vdd.n624 vss 0.0179f
C1961 vdd.n625 vss 0.0409f
C1962 vdd.n626 vss 0.0178f
C1963 vdd.n627 vss 0.00568f
C1964 vdd.n628 vss 0.0179f
C1965 vdd.n629 vss 0.0409f
C1966 vdd.n630 vss 0.0178f
C1967 vdd.n631 vss 0.00568f
C1968 vdd.n632 vss 0.00744f
C1969 vdd.n633 vss 0.00733f
C1970 vdd.n634 vss 0.0728f
C1971 vdd.n635 vss 0.19f
C1972 vdd.n636 vss 0.00744f
C1973 vdd.n637 vss 0.0728f
C1974 vdd.n638 vss 0.00733f
C1975 vdd.n639 vss 0.0179f
C1976 vdd.n640 vss 0.0409f
C1977 vdd.n641 vss 0.0178f
C1978 vdd.n642 vss 0.00568f
C1979 vdd.n643 vss 0.00744f
C1980 vdd.n644 vss 0.0728f
C1981 vdd.n645 vss 0.00733f
C1982 vdd.n646 vss 0.0179f
C1983 vdd.n647 vss 0.041f
C1984 vdd.n648 vss 0.0178f
C1985 vdd.t69 vss 0.00845f
C1986 vdd.n649 vss 0.122f
C1987 vdd.n650 vss 0.0179f
C1988 vdd.n651 vss 0.0173f
C1989 vdd.n652 vss 0.015f
C1990 vdd.n653 vss 0.00704f
C1991 vdd.n654 vss 0.0154f
C1992 vdd.n655 vss 0.00594f
C1993 vdd.t44 vss 0.00594f
C1994 vdd.t43 vss 0.00594f
C1995 vdd.n656 vss 0.0146f
C1996 vdd.n657 vss 0.0432f
C1997 vdd.n658 vss 0.00722f
C1998 vdd.n659 vss 0.0147f
C1999 vdd.n660 vss 0.0901f
C2000 vdd.n661 vss 0.101f
C2001 vdd.n662 vss 0.00973f
C2002 vdd.n663 vss 0.06f
C2003 vdd.n664 vss 0.0463f
C2004 vdd.n665 vss 0.0481f
C2005 vdd.t46 vss 0.0456f
C2006 vdd.n666 vss 0.0586f
C2007 vdd.n667 vss 0.0425f
C2008 vdd.n668 vss 0.0272f
C2009 vdd.t45 vss 0.251f
C2010 vdd.n669 vss 0.394f
C2011 vdd.n670 vss 0.198f
C2012 vdd.n671 vss 0.0253f
C2013 vdd.n672 vss 0.0253f
C2014 vdd.n673 vss 0.0284f
C2015 vdd.n674 vss 0.0424f
C2016 vdd.n675 vss 0.136f
C2017 vdd.n676 vss 0.385f
C2018 vdd.n677 vss 0.105f
C2019 vdd.n678 vss 0.00973f
C2020 vdd.n679 vss 0.0866f
C2021 vdd.n680 vss 0.0866f
C2022 vdd.n681 vss 0.00973f
C2023 vdd.n682 vss 0.0955f
C2024 vdd.n683 vss 0.0955f
C2025 vdd.n684 vss 0.00973f
C2026 vdd.n685 vss 0.0832f
C2027 vdd.n686 vss 0.0832f
C2028 vdd.n687 vss 0.00973f
C2029 vdd.n688 vss 0.0777f
C2030 vdd.n689 vss 0.0409f
C2031 vdd.n690 vss 0.0777f
C2032 vdd.n691 vss 0.00973f
C2033 vdd.n692 vss 0.00568f
C2034 vdd.n693 vss 0.00733f
C2035 vdd.n694 vss 0.0728f
C2036 vdd.n695 vss 0.125f
C2037 vdd.n696 vss 0.118f
C2038 vdd.t47 vss 0.285f
C2039 vdd.t68 vss 0.822f
C2040 vdd.n697 vss 0.0472f
C2041 vdd.n698 vss 0.581f
C2042 vdd.n699 vss 0.0161f
C2043 vdd.n700 vss 0.0374f
C2044 vdd.n701 vss 0.0378f
C2045 vdd.n702 vss 4.25e-19
C2046 vdd.n703 vss 0.00437f
C2047 vdd.n704 vss 0.00714f
C2048 vdd.n705 vss -0.168f
C2049 vdd.n706 vss 0.0082f
C2050 vdd.n707 vss 0.00502f
C2051 vdd.n708 vss 0.00518f
C2052 vdd.n709 vss 0.00836f
C2053 vdd.n710 vss 0.00714f
C2054 vdd.n711 vss 0.00437f
C2055 vdd.n712 vss 4.25e-19
C2056 vdd.n713 vss 0.00297f
C2057 vdd.n714 vss 0.00394f
C2058 vdd.n715 vss 0.00423f
C2059 vdd.n716 vss 0.00524f
C2060 vdd.n717 vss 0.00722f
C2061 vdd.n718 vss 0.00594f
C2062 vdd.n719 vss 0.00297f
C2063 vdd.n720 vss 0.00877f
C2064 vdd.n721 vss 0.00877f
C2065 vdd.n722 vss 0.0115f
C2066 vdd.n723 vss 0.219f
C2067 vdd.n724 vss 0.0472f
C2068 vdd.n725 vss 0.178f
C2069 vdd.n726 vss 0.00933f
C2070 vdd.n727 vss 2.83e-19
C2071 vdd.n728 vss 0.00241f
C2072 vdd.n729 vss 0.00877f
C2073 vdd.n730 vss 0.00297f
C2074 vdd.n731 vss 0.00594f
C2075 vdd.n732 vss 0.00722f
C2076 vdd.n733 vss 0.00368f
C2077 vdd.n734 vss 0.00524f
C2078 vdd.n735 vss -0.189f
C2079 vdd.n736 vss -0.0674f
C2080 vdd.n737 vss 0.00502f
C2081 vdd.n738 vss 0.00518f
C2082 vdd.n739 vss 0.0082f
C2083 vdd.n740 vss 0.00836f
C2084 vdd.n741 vss 0.00714f
C2085 vdd.n742 vss 0.00437f
C2086 vdd.n743 vss 4.25e-19
C2087 vdd.n744 vss 0.00311f
C2088 vdd.n745 vss 2.83e-19
C2089 vdd.n746 vss 0.00241f
C2090 vdd.n747 vss 0.00248f
C2091 vdd.n748 vss 0.0472f
C2092 vdd.n749 vss 0.178f
C2093 vdd.n750 vss 0.219f
C2094 vdd.n751 vss 0.0115f
C2095 vdd.n752 vss 0.00877f
C2096 vdd.n753 vss 0.00877f
C2097 vdd.n754 vss 0.00297f
C2098 vdd.n755 vss 0.00594f
C2099 vdd.n756 vss 0.00722f
C2100 vdd.n757 vss 0.00524f
C2101 vdd.n758 vss 0.00368f
C2102 vdd.n759 vss 0.00297f
C2103 vdd.n760 vss 0.00394f
C2104 vdd.n761 vss 2.92e-19
C2105 vdd.n762 vss 0.00437f
C2106 vdd.n763 vss 0.00714f
C2107 vdd.n764 vss -0.168f
C2108 vdd.n765 vss 0.0082f
C2109 vdd.n766 vss 0.00502f
C2110 vdd.n767 vss 0.00394f
C2111 vdd.n768 vss 0.00423f
C2112 vdd.n769 vss 0.00524f
C2113 vdd.n770 vss 0.00594f
C2114 vdd.n771 vss 0.00722f
C2115 vdd.n772 vss 0.00311f
C2116 vdd.n773 vss 0.00241f
C2117 vdd.n774 vss 0.00311f
C2118 vdd.n775 vss 2.83e-19
C2119 vdd.n776 vss 0.00933f
C2120 vdd.n777 vss 0.178f
C2121 vdd.n778 vss 0.219f
C2122 vdd.n779 vss 0.0472f
C2123 vdd.n780 vss 0.00248f
C2124 vdd.n781 vss 0.00241f
C2125 vdd.n782 vss 2.83e-19
C2126 vdd.n783 vss 0.00311f
C2127 vdd.n784 vss 4.25e-19
C2128 vdd.n785 vss 0.00437f
C2129 vdd.n786 vss 0.00714f
C2130 vdd.n787 vss 0.00836f
C2131 vdd.n788 vss 0.0082f
C2132 vdd.n789 vss 0.0257f
C2133 vdd.n790 vss 0.0296f
C2134 vdd.n791 vss 0.00518f
C2135 vdd.n792 vss 0.00502f
C2136 vdd.n793 vss -0.0674f
C2137 vdd.n794 vss -0.189f
C2138 vdd.n795 vss 0.00524f
C2139 vdd.n796 vss 0.00722f
C2140 vdd.n797 vss 0.00594f
C2141 vdd.n798 vss 0.00297f
C2142 vdd.n799 vss 0.00877f
C2143 vdd.n800 vss 0.00877f
C2144 vdd.n801 vss 0.0115f
C2145 vdd.n802 vss 0.219f
C2146 vdd.n803 vss 0.0472f
C2147 vdd.t49 vss 0.227f
C2148 vdd.n804 vss 0.186f
C2149 vdd.t94 vss 0.421f
C2150 vdd.n805 vss 0.111f
C2151 vdd.n806 vss 0.0211f
C2152 vdd.n807 vss 2.83e-19
C2153 vdd.n808 vss 0.00311f
C2154 vdd.n809 vss 4.25e-19
C2155 vdd.n810 vss 0.00311f
C2156 vdd.n811 vss 0.0256f
C2157 vdd.n812 vss 0.0256f
C2158 vdd.n813 vss 0.0234f
C2159 vdd.n814 vss 0.00297f
C2160 vdd.n815 vss 0.0263f
C2161 vdd.n816 vss 0.0263f
C2162 vdd.n817 vss 0.00241f
C2163 vdd.n818 vss 0.00241f
C2164 vdd.n819 vss 0.00311f
C2165 vdd.n820 vss 4.25e-19
C2166 vdd.n821 vss 0.00423f
C2167 vdd.n822 vss 2.92e-19
C2168 vdd.n823 vss 0.00502f
C2169 vdd.n824 vss 0.00518f
C2170 vdd.n825 vss 0.00423f
C2171 vdd.n826 vss 2.92e-19
C2172 vdd.n827 vss 0.00502f
C2173 vdd.n828 vss 0.0082f
C2174 vdd.n829 vss 0.00836f
C2175 vdd.n830 vss 0.0035f
C2176 vdd.n831 vss -0.189f
C2177 vdd.n832 vss 0.00524f
C2178 vdd.n833 vss 0.00311f
C2179 vdd.n834 vss 0.00722f
C2180 vdd.n835 vss 0.00594f
C2181 vdd.n836 vss 0.00297f
C2182 vdd.n837 vss 0.00877f
C2183 vdd.n838 vss 0.00877f
C2184 vdd.n839 vss 0.00241f
C2185 vdd.n840 vss 0.00248f
C2186 vdd.n841 vss 0.0472f
C2187 vdd.n842 vss 0.219f
C2188 vdd.n843 vss 0.178f
C2189 vdd.n844 vss 0.00933f
C2190 vdd.n845 vss 2.83e-19
C2191 vdd.n846 vss 0.00311f
C2192 vdd.n847 vss 0.00821f
C2193 vdd.n848 vss 0.00368f
C2194 vdd.n849 vss 0.00524f
C2195 vdd.n850 vss 0.00437f
C2196 vdd.n851 vss 0.0035f
C2197 vdd.n852 vss 0.00836f
C2198 vdd.n853 vss -0.175f
C2199 vdd.n854 vss -0.0772f
C2200 vdd.n855 vss 2.92e-19
C2201 vdd.n856 vss 0.00423f
C2202 vdd.n857 vss 4.25e-19
C2203 vdd.n858 vss 0.00311f
C2204 vdd.n859 vss 0.00241f
C2205 vdd.n860 vss 0.00297f
C2206 vdd.n861 vss 0.00877f
C2207 vdd.n862 vss 0.00877f
C2208 vdd.n863 vss 0.0115f
C2209 vdd.n864 vss 0.219f
C2210 vdd.n865 vss 0.178f
C2211 vdd.n866 vss 0.0472f
C2212 vdd.n867 vss 0.00248f
C2213 vdd.n868 vss 0.00241f
C2214 vdd.n869 vss 0.00877f
C2215 vdd.n870 vss 0.00877f
C2216 vdd.n871 vss 0.00297f
C2217 vdd.n872 vss 0.00594f
C2218 vdd.n873 vss 0.00722f
C2219 vdd.n874 vss 0.00524f
C2220 vdd.n875 vss 0.00437f
C2221 vdd.n876 vss 0.0035f
C2222 vdd.n877 vss 0.00836f
C2223 vdd.n878 vss 0.0082f
C2224 vdd.n879 vss 0.00502f
C2225 vdd.n880 vss 2.92e-19
C2226 vdd.n881 vss 0.00423f
C2227 vdd.n882 vss 4.25e-19
C2228 vdd.n883 vss 0.00311f
C2229 vdd.n884 vss 2.83e-19
C2230 vdd.n885 vss 0.00933f
C2231 vdd.n886 vss 0.178f
C2232 vdd.n887 vss 0.0472f
C2233 vdd.n888 vss 0.219f
C2234 vdd.n889 vss 0.0115f
C2235 vdd.n890 vss 0.00877f
C2236 vdd.n891 vss 0.00241f
C2237 vdd.n892 vss 0.00877f
C2238 vdd.n893 vss 0.00297f
C2239 vdd.n894 vss 0.00594f
C2240 vdd.n895 vss 0.00722f
C2241 vdd.n896 vss 0.00524f
C2242 vdd.n897 vss -0.189f
C2243 vdd.n898 vss 0.0035f
C2244 vdd.n899 vss 0.00836f
C2245 vdd.n900 vss 0.0082f
C2246 vdd.n901 vss 0.00502f
C2247 vdd.n902 vss 2.92e-19
C2248 vdd.n903 vss 0.00423f
C2249 vdd.n904 vss 4.25e-19
C2250 vdd.n905 vss 0.00311f
C2251 vdd.n906 vss 0.00821f
C2252 vdd.n907 vss 0.00368f
C2253 vdd.n908 vss 0.00524f
C2254 vdd.n909 vss 0.00437f
C2255 vdd.n910 vss 0.0035f
C2256 vdd.n911 vss 0.00836f
C2257 vdd.n912 vss -0.175f
C2258 vdd.n913 vss 0.00437f
C2259 vdd.n914 vss 0.0265f
C2260 vdd.n915 vss 0.00368f
C2261 vdd.n916 vss 0.0225f
C2262 vdd.n917 vss 0.00368f
C2263 vdd.n918 vss 0.0225f
C2264 vdd.n919 vss 0.00423f
C2265 vdd.n920 vss 0.00394f
C2266 vdd.n921 vss 0.00502f
C2267 vdd.n922 vss 0.00518f
C2268 vdd.n923 vss 0.0216f
C2269 vdd.n924 vss 0.0217f
C2270 vdd.n925 vss 0.0221f
C2271 vdd.n926 vss 0.00518f
C2272 vdd.n927 vss -0.0772f
C2273 vdd.n928 vss 2.92e-19
C2274 vdd.n929 vss 0.00423f
C2275 vdd.n930 vss 4.25e-19
C2276 vdd.n931 vss 0.00311f
C2277 vdd.n932 vss 0.00241f
C2278 vdd.n933 vss 0.00297f
C2279 vdd.n934 vss 0.00877f
C2280 vdd.n935 vss 0.00877f
C2281 vdd.n936 vss 0.00241f
C2282 vdd.n937 vss 0.00248f
C2283 vdd.n938 vss 0.0472f
C2284 vdd.n939 vss 0.219f
C2285 vdd.n940 vss 0.178f
C2286 vdd.n941 vss 0.00933f
C2287 vdd.n942 vss 2.83e-19
C2288 vdd.n943 vss 0.00241f
C2289 vdd.n944 vss 0.0269f
C2290 vdd.n945 vss 0.0166f
C2291 vdd.n946 vss 0.369f
C2292 vdd.n947 vss 0.203f
C2293 vdd.n948 vss 0.0472f
C2294 vdd.n949 vss 0.00248f
C2295 vdd.n950 vss 0.00241f
C2296 vdd.n951 vss 2.83e-19
C2297 vdd.n952 vss 0.00311f
C2298 vdd.n953 vss 4.25e-19
C2299 vdd.n954 vss 0.00437f
C2300 vdd.n955 vss 0.00714f
C2301 vdd.n956 vss -0.168f
C2302 vdd.n957 vss 0.0082f
C2303 vdd.n958 vss 0.00502f
C2304 vdd.n959 vss 0.00518f
C2305 vdd.n960 vss 0.00836f
C2306 vdd.n961 vss 0.00714f
C2307 vdd.n962 vss 0.00437f
C2308 vdd.n963 vss 4.25e-19
C2309 vdd.n964 vss 0.00297f
C2310 vdd.n965 vss 0.00394f
C2311 vdd.n966 vss 0.00423f
C2312 vdd.n967 vss 0.00524f
C2313 vdd.n968 vss 0.00722f
C2314 vdd.n969 vss 0.00594f
C2315 vdd.n970 vss 0.00297f
C2316 vdd.n971 vss 0.00877f
C2317 vdd.n972 vss 0.00877f
C2318 vdd.n973 vss 0.0115f
C2319 vdd.n974 vss 0.219f
C2320 vdd.n975 vss 0.0472f
C2321 vdd.n976 vss 0.178f
C2322 vdd.n977 vss 0.00933f
C2323 vdd.n978 vss 2.83e-19
C2324 vdd.n979 vss 0.00241f
C2325 vdd.n980 vss 0.00877f
C2326 vdd.n981 vss 0.00297f
C2327 vdd.n982 vss 0.00594f
C2328 vdd.n983 vss 0.00722f
C2329 vdd.n984 vss 0.00368f
C2330 vdd.n985 vss 0.00524f
C2331 vdd.n986 vss -0.189f
C2332 vdd.n987 vss -0.0674f
C2333 vdd.n988 vss 0.00502f
C2334 vdd.n989 vss 0.00518f
C2335 vdd.n990 vss 0.0082f
C2336 vdd.n991 vss 0.00836f
C2337 vdd.n992 vss 0.00714f
C2338 vdd.n993 vss 0.00437f
C2339 vdd.n994 vss 4.25e-19
C2340 vdd.n995 vss 0.00311f
C2341 vdd.n996 vss 2.83e-19
C2342 vdd.n997 vss 0.00241f
C2343 vdd.n998 vss 0.00248f
C2344 vdd.n999 vss 0.0472f
C2345 vdd.n1000 vss 0.178f
C2346 vdd.n1001 vss 0.219f
C2347 vdd.n1002 vss 0.0115f
C2348 vdd.n1003 vss 0.00877f
C2349 vdd.n1004 vss 0.00877f
C2350 vdd.n1005 vss 0.00297f
C2351 vdd.n1006 vss 0.00594f
C2352 vdd.n1007 vss 0.00722f
C2353 vdd.n1008 vss 0.00524f
C2354 vdd.n1009 vss 0.00368f
C2355 vdd.n1010 vss 0.00297f
C2356 vdd.n1011 vss 0.00394f
C2357 vdd.n1012 vss 2.92e-19
C2358 vdd.n1013 vss 0.00437f
C2359 vdd.n1014 vss 0.00714f
C2360 vdd.n1015 vss -0.168f
C2361 vdd.n1016 vss 0.0082f
C2362 vdd.n1017 vss 0.00502f
C2363 vdd.n1018 vss 0.00394f
C2364 vdd.n1019 vss 0.00423f
C2365 vdd.n1020 vss 0.00524f
C2366 vdd.n1021 vss 0.00594f
C2367 vdd.n1022 vss 0.00722f
C2368 vdd.n1023 vss 0.00311f
C2369 vdd.n1024 vss 0.00241f
C2370 vdd.n1025 vss 0.00311f
C2371 vdd.n1026 vss 2.83e-19
C2372 vdd.n1027 vss 0.00933f
C2373 vdd.n1028 vss 0.178f
C2374 vdd.n1029 vss 0.219f
C2375 vdd.n1030 vss 0.0472f
C2376 vdd.n1031 vss 0.00248f
C2377 vdd.n1032 vss 0.00241f
C2378 vdd.n1033 vss 2.83e-19
C2379 vdd.n1034 vss 0.00311f
C2380 vdd.n1035 vss 4.25e-19
C2381 vdd.n1036 vss 0.00437f
C2382 vdd.n1037 vss 0.00714f
C2383 vdd.n1038 vss 0.00836f
C2384 vdd.n1039 vss 0.0082f
C2385 vdd.n1040 vss 0.0257f
C2386 vdd.n1041 vss 0.0296f
C2387 vdd.n1042 vss 0.00518f
C2388 vdd.n1043 vss 0.00502f
C2389 vdd.n1044 vss -0.0674f
C2390 vdd.n1045 vss -0.189f
C2391 vdd.n1046 vss 0.00524f
C2392 vdd.n1047 vss 0.00722f
C2393 vdd.n1048 vss 0.00594f
C2394 vdd.n1049 vss 0.00297f
C2395 vdd.n1050 vss 0.00877f
C2396 vdd.n1051 vss 0.00877f
C2397 vdd.n1052 vss 0.0115f
C2398 vdd.n1053 vss 0.219f
C2399 vdd.n1054 vss 0.0472f
C2400 vdd.t40 vss 0.227f
C2401 vdd.n1055 vss 0.186f
C2402 vdd.t78 vss 0.421f
C2403 vdd.n1056 vss 0.111f
C2404 vdd.n1057 vss 0.0211f
C2405 vdd.n1058 vss 2.83e-19
C2406 vdd.n1059 vss 0.00311f
C2407 vdd.n1060 vss 4.25e-19
C2408 vdd.n1061 vss 0.00311f
C2409 vdd.n1062 vss 0.0256f
C2410 vdd.n1063 vss 0.0256f
C2411 vdd.n1064 vss 0.0234f
C2412 vdd.n1065 vss 0.00297f
C2413 vdd.n1066 vss 0.0263f
C2414 vdd.n1067 vss 0.0263f
C2415 vdd.n1068 vss 0.00241f
C2416 vdd.n1069 vss 0.00241f
C2417 vdd.n1070 vss 0.00311f
C2418 vdd.n1071 vss 4.25e-19
C2419 vdd.n1072 vss 0.00423f
C2420 vdd.n1073 vss 2.92e-19
C2421 vdd.n1074 vss 0.00502f
C2422 vdd.n1075 vss 0.00518f
C2423 vdd.n1076 vss 0.00423f
C2424 vdd.n1077 vss 2.92e-19
C2425 vdd.n1078 vss 0.00502f
C2426 vdd.n1079 vss 0.0082f
C2427 vdd.n1080 vss 0.00836f
C2428 vdd.n1081 vss 0.0035f
C2429 vdd.n1082 vss -0.189f
C2430 vdd.n1083 vss 0.00524f
C2431 vdd.n1084 vss 0.00311f
C2432 vdd.n1085 vss 0.00722f
C2433 vdd.n1086 vss 0.00594f
C2434 vdd.n1087 vss 0.00297f
C2435 vdd.n1088 vss 0.00877f
C2436 vdd.n1089 vss 0.00877f
C2437 vdd.n1090 vss 0.00241f
C2438 vdd.n1091 vss 0.00248f
C2439 vdd.n1092 vss 0.0472f
C2440 vdd.n1093 vss 0.219f
C2441 vdd.n1094 vss 0.178f
C2442 vdd.n1095 vss 0.00933f
C2443 vdd.n1096 vss 2.83e-19
C2444 vdd.n1097 vss 0.00311f
C2445 vdd.n1098 vss 0.00821f
C2446 vdd.n1099 vss 0.00368f
C2447 vdd.n1100 vss 0.00524f
C2448 vdd.n1101 vss 0.00437f
C2449 vdd.n1102 vss 0.0035f
C2450 vdd.n1103 vss 0.00836f
C2451 vdd.n1104 vss -0.175f
C2452 vdd.n1105 vss -0.0772f
C2453 vdd.n1106 vss 2.92e-19
C2454 vdd.n1107 vss 0.00423f
C2455 vdd.n1108 vss 4.25e-19
C2456 vdd.n1109 vss 0.00311f
C2457 vdd.n1110 vss 0.00241f
C2458 vdd.n1111 vss 0.00297f
C2459 vdd.n1112 vss 0.00877f
C2460 vdd.n1113 vss 0.00877f
C2461 vdd.n1114 vss 0.0115f
C2462 vdd.n1115 vss 0.219f
C2463 vdd.n1116 vss 0.178f
C2464 vdd.n1117 vss 0.0472f
C2465 vdd.n1118 vss 0.00248f
C2466 vdd.n1119 vss 0.00241f
C2467 vdd.n1120 vss 0.00877f
C2468 vdd.n1121 vss 0.00877f
C2469 vdd.n1122 vss 0.00297f
C2470 vdd.n1123 vss 0.00594f
C2471 vdd.n1124 vss 0.00722f
C2472 vdd.n1125 vss 0.00524f
C2473 vdd.n1126 vss 0.00437f
C2474 vdd.n1127 vss 0.0035f
C2475 vdd.n1128 vss 0.00836f
C2476 vdd.n1129 vss 0.0082f
C2477 vdd.n1130 vss 0.00502f
C2478 vdd.n1131 vss 2.92e-19
C2479 vdd.n1132 vss 0.00423f
C2480 vdd.n1133 vss 4.25e-19
C2481 vdd.n1134 vss 0.00311f
C2482 vdd.n1135 vss 2.83e-19
C2483 vdd.n1136 vss 0.00933f
C2484 vdd.n1137 vss 0.178f
C2485 vdd.n1138 vss 0.0472f
C2486 vdd.n1139 vss 0.219f
C2487 vdd.n1140 vss 0.0115f
C2488 vdd.n1141 vss 0.00877f
C2489 vdd.n1142 vss 0.00241f
C2490 vdd.n1143 vss 0.00877f
C2491 vdd.n1144 vss 0.00297f
C2492 vdd.n1145 vss 0.00594f
C2493 vdd.n1146 vss 0.00722f
C2494 vdd.n1147 vss 0.00524f
C2495 vdd.n1148 vss -0.189f
C2496 vdd.n1149 vss 0.0035f
C2497 vdd.n1150 vss 0.00836f
C2498 vdd.n1151 vss 0.0082f
C2499 vdd.n1152 vss 0.00502f
C2500 vdd.n1153 vss 2.92e-19
C2501 vdd.n1154 vss 0.00423f
C2502 vdd.n1155 vss 4.25e-19
C2503 vdd.n1156 vss 0.00311f
C2504 vdd.n1157 vss 0.00821f
C2505 vdd.n1158 vss 0.00368f
C2506 vdd.n1159 vss 0.00524f
C2507 vdd.n1160 vss 0.00437f
C2508 vdd.n1161 vss 0.0035f
C2509 vdd.n1162 vss 0.00836f
C2510 vdd.n1163 vss -0.175f
C2511 vdd.n1164 vss 0.00437f
C2512 vdd.n1165 vss 0.0265f
C2513 vdd.n1166 vss 0.00368f
C2514 vdd.n1167 vss 0.0225f
C2515 vdd.n1168 vss 0.00368f
C2516 vdd.n1169 vss 0.0225f
C2517 vdd.n1170 vss 0.00423f
C2518 vdd.n1171 vss 0.00394f
C2519 vdd.n1172 vss 0.00502f
C2520 vdd.n1173 vss 0.00518f
C2521 vdd.n1174 vss 0.0216f
C2522 vdd.n1175 vss 0.0217f
C2523 vdd.n1176 vss 0.0221f
C2524 vdd.n1177 vss 0.00518f
C2525 vdd.n1178 vss -0.0772f
C2526 vdd.n1179 vss 2.92e-19
C2527 vdd.n1180 vss 0.00423f
C2528 vdd.n1181 vss 4.25e-19
C2529 vdd.n1182 vss 0.00311f
C2530 vdd.n1183 vss 0.00241f
C2531 vdd.n1184 vss 0.00297f
C2532 vdd.n1185 vss 0.00877f
C2533 vdd.n1186 vss 0.00877f
C2534 vdd.n1187 vss 0.00241f
C2535 vdd.n1188 vss 0.00248f
C2536 vdd.n1189 vss 0.0472f
C2537 vdd.n1190 vss 0.219f
C2538 vdd.n1191 vss 0.178f
C2539 vdd.n1192 vss 0.00933f
C2540 vdd.n1193 vss 2.83e-19
C2541 vdd.n1194 vss 0.00241f
C2542 vdd.n1195 vss 0.0269f
C2543 vdd.n1196 vss 0.0166f
C2544 vdd.n1197 vss 0.369f
C2545 vdd.n1198 vss 0.203f
C2546 vdd.n1199 vss 0.0472f
C2547 vdd.n1200 vss 0.00248f
C2548 vdd.n1201 vss 0.00241f
C2549 vdd.n1202 vss 2.83e-19
C2550 vdd.n1203 vss 0.00311f
C2551 vdd.n1204 vss 4.25e-19
C2552 vdd.n1205 vss 0.00437f
C2553 vdd.n1206 vss 0.00714f
C2554 vdd.n1207 vss -0.168f
C2555 vdd.n1208 vss 0.0082f
C2556 vdd.n1209 vss 0.00502f
C2557 vdd.n1210 vss 0.00518f
C2558 vdd.n1211 vss 0.00836f
C2559 vdd.n1212 vss 0.00714f
C2560 vdd.n1213 vss 0.00437f
C2561 vdd.n1214 vss 4.25e-19
C2562 vdd.n1215 vss 0.00297f
C2563 vdd.n1216 vss 0.00394f
C2564 vdd.n1217 vss 0.00423f
C2565 vdd.n1218 vss 0.00524f
C2566 vdd.n1219 vss 0.00722f
C2567 vdd.n1220 vss 0.00594f
C2568 vdd.n1221 vss 0.00297f
C2569 vdd.n1222 vss 0.00877f
C2570 vdd.n1223 vss 0.00877f
C2571 vdd.n1224 vss 0.0115f
C2572 vdd.n1225 vss 0.219f
C2573 vdd.n1226 vss 0.0472f
C2574 vdd.n1227 vss 0.178f
C2575 vdd.n1228 vss 0.00933f
C2576 vdd.n1229 vss 2.83e-19
C2577 vdd.n1230 vss 0.00241f
C2578 vdd.n1231 vss 0.00877f
C2579 vdd.n1232 vss 0.00297f
C2580 vdd.n1233 vss 0.00594f
C2581 vdd.n1234 vss 0.00722f
C2582 vdd.n1235 vss 0.00368f
C2583 vdd.n1236 vss 0.00524f
C2584 vdd.n1237 vss -0.189f
C2585 vdd.n1238 vss -0.0674f
C2586 vdd.n1239 vss 0.00502f
C2587 vdd.n1240 vss 0.00518f
C2588 vdd.n1241 vss 0.0082f
C2589 vdd.n1242 vss 0.00836f
C2590 vdd.n1243 vss 0.00714f
C2591 vdd.n1244 vss 0.00437f
C2592 vdd.n1245 vss 4.25e-19
C2593 vdd.n1246 vss 0.00311f
C2594 vdd.n1247 vss 2.83e-19
C2595 vdd.n1248 vss 0.00241f
C2596 vdd.n1249 vss 0.00248f
C2597 vdd.n1250 vss 0.0472f
C2598 vdd.n1251 vss 0.178f
C2599 vdd.n1252 vss 0.219f
C2600 vdd.n1253 vss 0.0115f
C2601 vdd.n1254 vss 0.00877f
C2602 vdd.n1255 vss 0.00877f
C2603 vdd.n1256 vss 0.00297f
C2604 vdd.n1257 vss 0.00594f
C2605 vdd.n1258 vss 0.00722f
C2606 vdd.n1259 vss 0.00524f
C2607 vdd.n1260 vss 0.00368f
C2608 vdd.n1261 vss 0.00297f
C2609 vdd.n1262 vss 0.00394f
C2610 vdd.n1263 vss 2.92e-19
C2611 vdd.n1264 vss 0.00437f
C2612 vdd.n1265 vss 0.00714f
C2613 vdd.n1266 vss -0.168f
C2614 vdd.n1267 vss 0.0082f
C2615 vdd.n1268 vss 0.00502f
C2616 vdd.n1269 vss 0.00394f
C2617 vdd.n1270 vss 0.00423f
C2618 vdd.n1271 vss 0.00524f
C2619 vdd.n1272 vss 0.00594f
C2620 vdd.n1273 vss 0.00722f
C2621 vdd.n1274 vss 0.00311f
C2622 vdd.n1275 vss 0.00241f
C2623 vdd.n1276 vss 0.00311f
C2624 vdd.n1277 vss 2.83e-19
C2625 vdd.n1278 vss 0.00933f
C2626 vdd.n1279 vss 0.178f
C2627 vdd.n1280 vss 0.219f
C2628 vdd.n1281 vss 0.0472f
C2629 vdd.n1282 vss 0.00248f
C2630 vdd.n1283 vss 0.00241f
C2631 vdd.n1284 vss 2.83e-19
C2632 vdd.n1285 vss 0.00311f
C2633 vdd.n1286 vss 4.25e-19
C2634 vdd.n1287 vss 0.00437f
C2635 vdd.n1288 vss 0.00714f
C2636 vdd.n1289 vss 0.00836f
C2637 vdd.n1290 vss 0.0082f
C2638 vdd.n1291 vss 0.0257f
C2639 vdd.n1292 vss 0.0296f
C2640 vdd.n1293 vss 0.00518f
C2641 vdd.n1294 vss 0.00502f
C2642 vdd.n1295 vss -0.0674f
C2643 vdd.n1296 vss -0.189f
C2644 vdd.n1297 vss 0.00524f
C2645 vdd.n1298 vss 0.00722f
C2646 vdd.n1299 vss 0.00594f
C2647 vdd.n1300 vss 0.00297f
C2648 vdd.n1301 vss 0.00877f
C2649 vdd.n1302 vss 0.00877f
C2650 vdd.n1303 vss 0.0115f
C2651 vdd.n1304 vss 0.219f
C2652 vdd.n1305 vss 0.0472f
C2653 vdd.t88 vss 0.227f
C2654 vdd.n1306 vss 0.186f
C2655 vdd.t42 vss 0.421f
C2656 vdd.n1307 vss 0.111f
C2657 vdd.n1308 vss 0.0211f
C2658 vdd.n1309 vss 2.83e-19
C2659 vdd.n1310 vss 0.00311f
C2660 vdd.n1311 vss 4.25e-19
C2661 vdd.n1312 vss 0.00311f
C2662 vdd.n1313 vss 0.0256f
C2663 vdd.n1314 vss 0.0256f
C2664 vdd.n1315 vss 0.0234f
C2665 vdd.n1316 vss 0.00297f
C2666 vdd.n1317 vss 0.0263f
C2667 vdd.n1318 vss 0.0263f
C2668 vdd.n1319 vss 0.00241f
C2669 vdd.n1320 vss 0.00241f
C2670 vdd.n1321 vss 0.00311f
C2671 vdd.n1322 vss 4.25e-19
C2672 vdd.n1323 vss 0.00423f
C2673 vdd.n1324 vss 2.92e-19
C2674 vdd.n1325 vss 0.00502f
C2675 vdd.n1326 vss 0.00518f
C2676 vdd.n1327 vss 0.00423f
C2677 vdd.n1328 vss 2.92e-19
C2678 vdd.n1329 vss 0.00502f
C2679 vdd.n1330 vss 0.0082f
C2680 vdd.n1331 vss 0.00836f
C2681 vdd.n1332 vss 0.0035f
C2682 vdd.n1333 vss -0.189f
C2683 vdd.n1334 vss 0.00524f
C2684 vdd.n1335 vss 0.00311f
C2685 vdd.n1336 vss 0.00722f
C2686 vdd.n1337 vss 0.00594f
C2687 vdd.n1338 vss 0.00297f
C2688 vdd.n1339 vss 0.00877f
C2689 vdd.n1340 vss 0.00877f
C2690 vdd.n1341 vss 0.00241f
C2691 vdd.n1342 vss 0.00248f
C2692 vdd.n1343 vss 0.0472f
C2693 vdd.n1344 vss 0.219f
C2694 vdd.n1345 vss 0.178f
C2695 vdd.n1346 vss 0.00933f
C2696 vdd.n1347 vss 2.83e-19
C2697 vdd.n1348 vss 0.00311f
C2698 vdd.n1349 vss 0.00821f
C2699 vdd.n1350 vss 0.00368f
C2700 vdd.n1351 vss 0.00524f
C2701 vdd.n1352 vss 0.00437f
C2702 vdd.n1353 vss 0.0035f
C2703 vdd.n1354 vss 0.00836f
C2704 vdd.n1355 vss -0.175f
C2705 vdd.n1356 vss -0.0772f
C2706 vdd.n1357 vss 2.92e-19
C2707 vdd.n1358 vss 0.00423f
C2708 vdd.n1359 vss 4.25e-19
C2709 vdd.n1360 vss 0.00311f
C2710 vdd.n1361 vss 0.00241f
C2711 vdd.n1362 vss 0.00297f
C2712 vdd.n1363 vss 0.00877f
C2713 vdd.n1364 vss 0.00877f
C2714 vdd.n1365 vss 0.0115f
C2715 vdd.n1366 vss 0.219f
C2716 vdd.n1367 vss 0.178f
C2717 vdd.n1368 vss 0.0472f
C2718 vdd.n1369 vss 0.00248f
C2719 vdd.n1370 vss 0.00241f
C2720 vdd.n1371 vss 0.00877f
C2721 vdd.n1372 vss 0.00877f
C2722 vdd.n1373 vss 0.00297f
C2723 vdd.n1374 vss 0.00594f
C2724 vdd.n1375 vss 0.00722f
C2725 vdd.n1376 vss 0.00524f
C2726 vdd.n1377 vss 0.00437f
C2727 vdd.n1378 vss 0.0035f
C2728 vdd.n1379 vss 0.00836f
C2729 vdd.n1380 vss 0.0082f
C2730 vdd.n1381 vss 0.00502f
C2731 vdd.n1382 vss 2.92e-19
C2732 vdd.n1383 vss 0.00423f
C2733 vdd.n1384 vss 4.25e-19
C2734 vdd.n1385 vss 0.00311f
C2735 vdd.n1386 vss 2.83e-19
C2736 vdd.n1387 vss 0.00933f
C2737 vdd.n1388 vss 0.178f
C2738 vdd.n1389 vss 0.0472f
C2739 vdd.n1390 vss 0.219f
C2740 vdd.n1391 vss 0.0115f
C2741 vdd.n1392 vss 0.00877f
C2742 vdd.n1393 vss 0.00241f
C2743 vdd.n1394 vss 0.00877f
C2744 vdd.n1395 vss 0.00297f
C2745 vdd.n1396 vss 0.00594f
C2746 vdd.n1397 vss 0.00722f
C2747 vdd.n1398 vss 0.00524f
C2748 vdd.n1399 vss -0.189f
C2749 vdd.n1400 vss 0.0035f
C2750 vdd.n1401 vss 0.00836f
C2751 vdd.n1402 vss 0.0082f
C2752 vdd.n1403 vss 0.00502f
C2753 vdd.n1404 vss 2.92e-19
C2754 vdd.n1405 vss 0.00423f
C2755 vdd.n1406 vss 4.25e-19
C2756 vdd.n1407 vss 0.00311f
C2757 vdd.n1408 vss 0.00821f
C2758 vdd.n1409 vss 0.00368f
C2759 vdd.n1410 vss 0.00524f
C2760 vdd.n1411 vss 0.00437f
C2761 vdd.n1412 vss 0.0035f
C2762 vdd.n1413 vss 0.00836f
C2763 vdd.n1414 vss -0.175f
C2764 vdd.n1415 vss 0.00437f
C2765 vdd.n1416 vss 0.0265f
C2766 vdd.n1417 vss 0.00368f
C2767 vdd.n1418 vss 0.0225f
C2768 vdd.n1419 vss 0.00368f
C2769 vdd.n1420 vss 0.0225f
C2770 vdd.n1421 vss 0.00423f
C2771 vdd.n1422 vss 0.00394f
C2772 vdd.n1423 vss 0.00502f
C2773 vdd.n1424 vss 0.00518f
C2774 vdd.n1425 vss 0.0216f
C2775 vdd.n1426 vss 0.0217f
C2776 vdd.n1427 vss 0.0221f
C2777 vdd.n1428 vss 0.00518f
C2778 vdd.n1429 vss -0.0772f
C2779 vdd.n1430 vss 2.92e-19
C2780 vdd.n1431 vss 0.00423f
C2781 vdd.n1432 vss 4.25e-19
C2782 vdd.n1433 vss 0.00311f
C2783 vdd.n1434 vss 0.00241f
C2784 vdd.n1435 vss 0.00297f
C2785 vdd.n1436 vss 0.00877f
C2786 vdd.n1437 vss 0.00877f
C2787 vdd.n1438 vss 0.00241f
C2788 vdd.n1439 vss 0.00248f
C2789 vdd.n1440 vss 0.0472f
C2790 vdd.n1441 vss 0.219f
C2791 vdd.n1442 vss 0.178f
C2792 vdd.n1443 vss 0.00933f
C2793 vdd.n1444 vss 2.83e-19
C2794 vdd.n1445 vss 0.00241f
C2795 vdd.n1446 vss 0.0269f
C2796 vdd.n1447 vss 0.0166f
C2797 vdd.n1448 vss 0.369f
C2798 vdd.n1449 vss 0.203f
C2799 vdd.n1450 vss 0.0472f
C2800 vdd.n1451 vss 0.00248f
C2801 vdd.n1452 vss 0.00241f
C2802 vdd.n1453 vss 2.83e-19
C2803 vdd.n1454 vss 0.00311f
C2804 vdd.n1455 vss 4.25e-19
C2805 vdd.n1456 vss 0.00437f
C2806 vdd.n1457 vss 0.00714f
C2807 vdd.n1458 vss -0.168f
C2808 vdd.n1459 vss 0.0082f
C2809 vdd.n1460 vss 0.00502f
C2810 vdd.n1461 vss 0.00518f
C2811 vdd.n1462 vss 0.00836f
C2812 vdd.n1463 vss 0.00714f
C2813 vdd.n1464 vss 0.00437f
C2814 vdd.n1465 vss 4.25e-19
C2815 vdd.n1466 vss 0.00297f
C2816 vdd.n1467 vss 0.00394f
C2817 vdd.n1468 vss 0.00423f
C2818 vdd.n1469 vss 0.00524f
C2819 vdd.n1470 vss 0.00722f
C2820 vdd.n1471 vss 0.00594f
C2821 vdd.n1472 vss 0.00297f
C2822 vdd.n1473 vss 0.00877f
C2823 vdd.n1474 vss 0.00877f
C2824 vdd.n1475 vss 0.0115f
C2825 vdd.n1476 vss 0.219f
C2826 vdd.n1477 vss 0.0472f
C2827 vdd.n1478 vss 0.178f
C2828 vdd.n1479 vss 0.00933f
C2829 vdd.n1480 vss 2.83e-19
C2830 vdd.n1481 vss 0.00241f
C2831 vdd.n1482 vss 0.00877f
C2832 vdd.n1483 vss 0.00297f
C2833 vdd.n1484 vss 0.00594f
C2834 vdd.n1485 vss 0.00722f
C2835 vdd.n1486 vss 0.00368f
C2836 vdd.n1487 vss 0.00524f
C2837 vdd.n1488 vss -0.189f
C2838 vdd.n1489 vss -0.0674f
C2839 vdd.n1490 vss 0.00502f
C2840 vdd.n1491 vss 0.00518f
C2841 vdd.n1492 vss 0.0082f
C2842 vdd.n1493 vss 0.00836f
C2843 vdd.n1494 vss 0.00714f
C2844 vdd.n1495 vss 0.00437f
C2845 vdd.n1496 vss 4.25e-19
C2846 vdd.n1497 vss 0.00311f
C2847 vdd.n1498 vss 2.83e-19
C2848 vdd.n1499 vss 0.00241f
C2849 vdd.n1500 vss 0.00248f
C2850 vdd.n1501 vss 0.0472f
C2851 vdd.n1502 vss 0.178f
C2852 vdd.n1503 vss 0.219f
C2853 vdd.n1504 vss 0.0115f
C2854 vdd.n1505 vss 0.00877f
C2855 vdd.n1506 vss 0.00877f
C2856 vdd.n1507 vss 0.00297f
C2857 vdd.n1508 vss 0.00594f
C2858 vdd.n1509 vss 0.00722f
C2859 vdd.n1510 vss 0.00524f
C2860 vdd.n1511 vss 0.00368f
C2861 vdd.n1512 vss 0.00297f
C2862 vdd.n1513 vss 0.00394f
C2863 vdd.n1514 vss 2.92e-19
C2864 vdd.n1515 vss 0.00437f
C2865 vdd.n1516 vss 0.00714f
C2866 vdd.n1517 vss -0.168f
C2867 vdd.n1518 vss 0.0082f
C2868 vdd.n1519 vss 0.00502f
C2869 vdd.n1520 vss 0.00394f
C2870 vdd.n1521 vss 0.00423f
C2871 vdd.n1522 vss 0.00524f
C2872 vdd.n1523 vss 0.00594f
C2873 vdd.n1524 vss 0.00722f
C2874 vdd.n1525 vss 0.00311f
C2875 vdd.n1526 vss 0.00241f
C2876 vdd.n1527 vss 0.00311f
C2877 vdd.n1528 vss 2.83e-19
C2878 vdd.n1529 vss 0.00933f
C2879 vdd.n1530 vss 0.178f
C2880 vdd.n1531 vss 0.219f
C2881 vdd.n1532 vss 0.0472f
C2882 vdd.n1533 vss 0.00248f
C2883 vdd.n1534 vss 0.00241f
C2884 vdd.n1535 vss 2.83e-19
C2885 vdd.n1536 vss 0.00311f
C2886 vdd.n1537 vss 4.25e-19
C2887 vdd.n1538 vss 0.00437f
C2888 vdd.n1539 vss 0.00714f
C2889 vdd.n1540 vss 0.00836f
C2890 vdd.n1541 vss 0.0082f
C2891 vdd.n1542 vss 0.0257f
C2892 vdd.n1543 vss 0.0296f
C2893 vdd.n1544 vss 0.00518f
C2894 vdd.n1545 vss 0.00502f
C2895 vdd.n1546 vss -0.0674f
C2896 vdd.n1547 vss -0.189f
C2897 vdd.n1548 vss 0.00524f
C2898 vdd.n1549 vss 0.00722f
C2899 vdd.n1550 vss 0.00594f
C2900 vdd.n1551 vss 0.00297f
C2901 vdd.n1552 vss 0.00877f
C2902 vdd.n1553 vss 0.00877f
C2903 vdd.n1554 vss 0.0115f
C2904 vdd.n1555 vss 0.219f
C2905 vdd.n1556 vss 0.0472f
C2906 vdd.t63 vss 0.227f
C2907 vdd.n1557 vss 0.186f
C2908 vdd.t73 vss 0.421f
C2909 vdd.n1558 vss 0.111f
C2910 vdd.n1559 vss 0.0211f
C2911 vdd.n1560 vss 2.83e-19
C2912 vdd.n1561 vss 0.00311f
C2913 vdd.n1562 vss 4.25e-19
C2914 vdd.n1563 vss 0.00311f
C2915 vdd.n1564 vss 0.0256f
C2916 vdd.n1565 vss 0.0256f
C2917 vdd.n1566 vss 0.0234f
C2918 vdd.n1567 vss 0.00297f
C2919 vdd.n1568 vss 0.0263f
C2920 vdd.n1569 vss 0.0263f
C2921 vdd.n1570 vss 0.00241f
C2922 vdd.n1571 vss 0.00241f
C2923 vdd.n1572 vss 0.00311f
C2924 vdd.n1573 vss 4.25e-19
C2925 vdd.n1574 vss 0.00423f
C2926 vdd.n1575 vss 2.92e-19
C2927 vdd.n1576 vss 0.00502f
C2928 vdd.n1577 vss 0.00518f
C2929 vdd.n1578 vss 0.00836f
C2930 vdd.n1579 vss 0.0035f
C2931 vdd.n1580 vss -0.189f
C2932 vdd.n1581 vss 0.00524f
C2933 vdd.n1582 vss 0.00722f
C2934 vdd.n1583 vss 0.00594f
C2935 vdd.n1584 vss 0.00297f
C2936 vdd.n1585 vss 0.00877f
C2937 vdd.n1586 vss 0.00877f
C2938 vdd.n1587 vss 0.00241f
C2939 vdd.n1588 vss 0.00248f
C2940 vdd.n1589 vss 0.0472f
C2941 vdd.n1590 vss 0.219f
C2942 vdd.n1591 vss 0.178f
C2943 vdd.n1592 vss 0.00933f
C2944 vdd.n1593 vss 2.83e-19
C2945 vdd.n1594 vss 0.00311f
C2946 vdd.n1595 vss 4.25e-19
C2947 vdd.n1596 vss 0.00423f
C2948 vdd.n1597 vss 2.92e-19
C2949 vdd.n1598 vss 0.00502f
C2950 vdd.n1599 vss 0.00518f
C2951 vdd.n1600 vss -0.175f
C2952 vdd.n1601 vss 0.00836f
C2953 vdd.n1602 vss 0.0035f
C2954 vdd.n1603 vss 0.00437f
C2955 vdd.n1604 vss 0.00524f
C2956 vdd.n1605 vss 0.00722f
C2957 vdd.n1606 vss 0.00311f
C2958 vdd.n1607 vss 0.00241f
C2959 vdd.n1608 vss 0.00297f
C2960 vdd.n1609 vss 0.00877f
C2961 vdd.n1610 vss 0.00877f
C2962 vdd.n1611 vss 0.0115f
C2963 vdd.n1612 vss 0.219f
C2964 vdd.n1613 vss 0.178f
C2965 vdd.n1614 vss 0.0472f
C2966 vdd.n1615 vss 0.00248f
C2967 vdd.n1616 vss 0.00241f
C2968 vdd.n1617 vss 0.00877f
C2969 vdd.n1618 vss 0.00877f
C2970 vdd.n1619 vss 0.00297f
C2971 vdd.n1620 vss 0.00311f
C2972 vdd.n1621 vss 0.00722f
C2973 vdd.n1622 vss 0.00594f
C2974 vdd.n1623 vss 0.00821f
C2975 vdd.n1624 vss 0.00368f
C2976 vdd.n1625 vss 0.00297f
C2977 vdd.n1626 vss 0.00394f
C2978 vdd.n1627 vss 0.00518f
C2979 vdd.n1628 vss 0.00836f
C2980 vdd.n1629 vss 0.0035f
C2981 vdd.n1630 vss 0.007f
C2982 vdd.n1631 vss 0.00423f
C2983 vdd.n1632 vss 2.92e-19
C2984 vdd.n1633 vss 0.00502f
C2985 vdd.n1634 vss 0.00518f
C2986 vdd.n1635 vss 0.00836f
C2987 vdd.n1636 vss 0.0035f
C2988 vdd.n1637 vss -0.189f
C2989 vdd.n1638 vss 0.00524f
C2990 vdd.n1639 vss 0.00368f
C2991 vdd.n1640 vss 0.00821f
C2992 vdd.n1641 vss 0.00311f
C2993 vdd.n1642 vss 2.83e-19
C2994 vdd.n1643 vss 0.00933f
C2995 vdd.n1644 vss 0.178f
C2996 vdd.n1645 vss 0.0472f
C2997 vdd.n1646 vss 0.219f
C2998 vdd.n1647 vss 0.0115f
C2999 vdd.n1648 vss 0.00877f
C3000 vdd.n1649 vss 0.00877f
C3001 vdd.n1650 vss 0.00241f
C3002 vdd.n1651 vss 0.00241f
C3003 vdd.n1652 vss 0.00311f
C3004 vdd.n1653 vss 4.25e-19
C3005 vdd.n1654 vss 0.00423f
C3006 vdd.n1655 vss 2.92e-19
C3007 vdd.n1656 vss 0.00502f
C3008 vdd.n1657 vss 0.00518f
C3009 vdd.n1658 vss 0.00423f
C3010 vdd.n1659 vss 2.92e-19
C3011 vdd.n1660 vss -0.0772f
C3012 vdd.n1661 vss -0.175f
C3013 vdd.n1662 vss 0.00836f
C3014 vdd.n1663 vss 0.0035f
C3015 vdd.n1664 vss 0.00437f
C3016 vdd.n1665 vss 0.00524f
C3017 vdd.n1666 vss 0.00311f
C3018 vdd.n1667 vss 0.00722f
C3019 vdd.n1668 vss 0.00594f
C3020 vdd.n1669 vss 0.00297f
C3021 vdd.n1670 vss 0.00877f
C3022 vdd.n1671 vss 0.00877f
C3023 vdd.n1672 vss 0.00241f
C3024 vdd.n1673 vss 0.00248f
C3025 vdd.n1674 vss 0.0472f
C3026 vdd.n1675 vss 0.219f
C3027 vdd.t81 vss 0.611f
C3028 vdd.n1676 vss 0.37f
C3029 vdd.n1677 vss 0.0472f
C3030 vdd.n1678 vss 0.178f
C3031 vdd.n1679 vss 0.00933f
C3032 vdd.n1680 vss 0.0374f
C3033 vdd.n1681 vss 0.0378f
C3034 vdd.n1682 vss 0.0349f
C3035 vdd.n1683 vss 0.0357f
C3036 vdd.n1684 vss 0.0221f
C3037 vdd.n1685 vss 0.0349f
C3038 vdd.n1686 vss 0.0516f
C3039 vdd.n1687 vss 0.00297f
C3040 vdd.n1688 vss 0.0388f
C3041 vdd.n1689 vss 0.0393f
C3042 vdd.n1690 vss 2.92e-19
C3043 vdd.n1691 vss 0.00521f
C3044 vdd.n1692 vss 0.00538f
C3045 vdd.n1693 vss 0.00868f
C3046 vdd.n1694 vss 0.0035f
C3047 vdd.n1695 vss -0.189f
C3048 vdd.n1696 vss 0.00524f
C3049 vdd.n1697 vss 0.00722f
C3050 vdd.n1698 vss 0.00594f
C3051 vdd.n1699 vss 0.00297f
C3052 vdd.n1700 vss 0.00877f
C3053 vdd.n1701 vss 0.00877f
C3054 vdd.n1702 vss 0.00241f
C3055 vdd.n1703 vss 0.00248f
C3056 vdd.n1704 vss 0.0472f
C3057 vdd.n1705 vss 0.219f
C3058 vdd.n1706 vss 0.178f
C3059 vdd.n1707 vss 0.00933f
C3060 vdd.n1708 vss 2.83e-19
C3061 vdd.n1709 vss 0.00311f
C3062 vdd.n1710 vss 4.25e-19
C3063 vdd.n1711 vss 0.00423f
C3064 vdd.n1712 vss 2.92e-19
C3065 vdd.n1713 vss 0.00521f
C3066 vdd.n1714 vss 0.00538f
C3067 vdd.n1715 vss -0.174f
C3068 vdd.n1716 vss 0.00868f
C3069 vdd.n1717 vss 0.0035f
C3070 vdd.n1718 vss 0.00437f
C3071 vdd.n1719 vss 0.00524f
C3072 vdd.n1720 vss 0.00722f
C3073 vdd.n1721 vss 0.00311f
C3074 vdd.n1722 vss 0.00241f
C3075 vdd.n1723 vss 0.00297f
C3076 vdd.n1724 vss 0.00877f
C3077 vdd.n1725 vss 0.00877f
C3078 vdd.n1726 vss 0.0115f
C3079 vdd.n1727 vss 0.219f
C3080 vdd.n1728 vss 0.178f
C3081 vdd.n1729 vss 0.0472f
C3082 vdd.n1730 vss 0.00248f
C3083 vdd.n1731 vss 0.00241f
C3084 vdd.n1732 vss 0.00877f
C3085 vdd.n1733 vss 0.00877f
C3086 vdd.n1734 vss 0.00297f
C3087 vdd.n1735 vss -0.00382f
C3088 vdd.n1736 vss -0.132f
C3089 vdd.n1737 vss 0.00594f
C3090 vdd.n1738 vss 0.00821f
C3091 vdd.n1739 vss 0.00368f
C3092 vdd.n1740 vss 0.00297f
C3093 vdd.n1741 vss 0.00394f
C3094 vdd.n1742 vss 0.00538f
C3095 vdd.n1743 vss 0.00868f
C3096 vdd.n1744 vss 0.0035f
C3097 vdd.n1745 vss 0.007f
C3098 vdd.n1746 vss 0.00423f
C3099 vdd.n1747 vss 2.92e-19
C3100 vdd.n1748 vss 0.00521f
C3101 vdd.n1749 vss 0.00538f
C3102 vdd.n1750 vss 0.00868f
C3103 vdd.n1751 vss 0.0035f
C3104 vdd.n1752 vss -0.189f
C3105 vdd.n1753 vss 0.00524f
C3106 vdd.n1754 vss 0.00368f
C3107 vdd.n1755 vss 0.00821f
C3108 vdd.n1756 vss 0.00311f
C3109 vdd.n1757 vss 2.83e-19
C3110 vdd.n1758 vss 0.00933f
C3111 vdd.n1759 vss 0.178f
C3112 vdd.n1760 vss 0.0472f
C3113 vdd.n1761 vss 0.219f
C3114 vdd.n1762 vss 0.0115f
C3115 vdd.n1763 vss 0.00877f
C3116 vdd.n1764 vss 0.00877f
C3117 vdd.n1765 vss 0.00241f
C3118 vdd.n1766 vss 0.00241f
C3119 vdd.n1767 vss 0.00311f
C3120 vdd.n1768 vss 4.25e-19
C3121 vdd.n1769 vss 0.00423f
C3122 vdd.n1770 vss 2.92e-19
C3123 vdd.n1771 vss 0.00521f
C3124 vdd.n1772 vss 0.00538f
C3125 vdd.n1773 vss 0.00868f
C3126 vdd.n1774 vss 0.0035f
C3127 vdd.n1775 vss 0.00437f
C3128 vdd.n1776 vss 0.00524f
C3129 vdd.n1777 vss 0.00722f
C3130 vdd.n1778 vss 0.00594f
C3131 vdd.n1779 vss 0.00297f
C3132 vdd.n1780 vss 0.00877f
C3133 vdd.n1781 vss 0.00877f
C3134 vdd.n1782 vss 0.00241f
C3135 vdd.n1783 vss 0.00248f
C3136 vdd.n1784 vss 0.0472f
C3137 vdd.n1785 vss 0.219f
C3138 vdd.t90 vss 0.0456f
C3139 vdd.n1786 vss 0.0502f
C3140 vdd.n1787 vss 0.0154f
C3141 vdd.t65 vss 0.0456f
C3142 vdd.n1788 vss 0.0834f
C3143 vdd.n1789 vss 0.0181f
C3144 vdd.n1790 vss 0.00714f
C3145 vdd.n1791 vss 0.0498f
C3146 vdd.n1792 vss 0.0201f
C3147 vdd.n1793 vss 0.00618f
C3148 vdd.n1794 vss 0.0153f
C3149 vdd.n1795 vss 0.0208f
C3150 vdd.n1796 vss 0.00991f
C3151 vdd.n1797 vss 0.0167f
C3152 vdd.n1798 vss 0.0367f
C3153 vdd.n1799 vss 0.0143f
C3154 vdd.n1800 vss 0.0118f
C3155 vdd.n1801 vss 7.3e-19
C3156 vdd.n1802 vss 0.0177f
C3157 vdd.n1803 vss 0.0189f
C3158 vdd.n1804 vss 0.00886f
C3159 vdd.n1805 vss 0.0191f
C3160 vdd.n1806 vss 0.00782f
C3161 vdd.n1807 vss 0.00365f
C3162 vdd.n1808 vss 0.00397f
C3163 vdd.n1809 vss 0.0543f
C3164 vdd.n1810 vss 0.0246f
C3165 vdd.n1811 vss 0.0119f
C3166 vdd.n1812 vss 0.0177f
C3167 vdd.n1813 vss 7.3e-19
C3168 vdd.n1814 vss 0.0234f
C3169 vdd.n1815 vss 0.0179f
C3170 vdd.n1816 vss 0.00618f
C3171 vdd.n1817 vss 0.0111f
C3172 vdd.n1818 vss 0.00602f
C3173 vdd.n1819 vss 0.00413f
C3174 vdd.n1820 vss 0.00432f
C3175 vdd.n1821 vss 0.00165f
C3176 vdd.n1822 vss 0.0098f
C3177 vdd.n1823 vss 0.00968f
C3178 vdd.n1824 vss 0.00229f
C3179 vdd.n1825 vss 0.0112f
C3180 vdd.n1826 vss 0.00146f
C3181 vdd.t89 vss 0.112f
C3182 vdd.t64 vss 0.0921f
C3183 vdd.n1827 vss 0.0677f
C3184 vdd.n1828 vss 0.0134f
C3185 vdd.n1829 vss 0.0818f
C3186 vdd.n1830 vss 0.0125f
C3187 vdd.n1831 vss 0.00121f
C3188 vdd.n1832 vss 0.00229f
C3189 vdd.n1833 vss 0.0035f
C3190 vdd.n1834 vss 0.0035f
C3191 vdd.n1835 vss 0.0165f
C3192 vdd.n1836 vss 0.0245f
C3193 vdd.n1837 vss 0.00954f
C3194 vdd.n1838 vss 0.00714f
C3195 vdd.n1839 vss 0.0281f
C3196 vdd.n1840 vss 0.0567f
C3197 vdd.t51 vss 0.673f
C3198 vdd.n1841 vss 0.374f
C3199 vdd.t52 vss 0.00523f
C3200 vdd.n1842 vss 0.0323f
C3201 vdd.n1843 vss 0.0513f
C3202 vdd.n1844 vss 0.0573f
C3203 vdd.n1845 vss 0.00802f
C3204 vdd.n1846 vss 0.0166f
C3205 vdd.n1847 vss 0.0916f
C3206 vdd.n1848 vss 0.0472f
C3207 vdd.n1849 vss 0.178f
C3208 vdd.n1850 vss 0.00933f
C3209 vdd.n1851 vss 2.83e-19
C3210 vdd.n1852 vss 0.00311f
C3211 vdd.n1853 vss 4.25e-19
C3212 vdd.n1854 vss 0.00423f
C3213 vdd.n1855 vss 2.92e-19
C3214 vdd.n1856 vss -0.077f
C3215 vdd.n1857 vss 0.00538f
C3216 vdd.n1858 vss 0.0116f
C3217 vdd.n1859 vss 0.0238f
C3218 vdd.n1860 vss 0.00573f
C3219 vdd.n1861 vss 0.00687f
C3220 vdd.n1862 vss 0.00437f
C3221 vdd.n1863 vss 0.00698f
C3222 vdd.n1864 vss 0.0109f
C3223 vdd.n1865 vss 0.00553f
C3224 vdd.n1866 vss 0.00996f
C3225 vdd.n1867 vss 9.51e-19
C3226 vdd.n1868 vss 0.00664f
C3227 vdd.n1869 vss 0.825f
C3228 vdd.n1870 vss 0.0119f
C3229 vdd.n1871 vss 0.0192f
C3230 vdd.n1872 vss 0.0111f
C3231 vdd.n1873 vss 0.0155f
C3232 vdd.n1874 vss 0.00731f
C3233 vdd.n1875 vss 0.00368f
C3234 vdd.n1876 vss 0.00394f
C3235 vdd.n1877 vss -0.174f
C3236 vdd.n1878 vss 0.007f
C3237 vdd.n1879 vss 0.00311f
C3238 vdd.n1880 vss 0.00297f
C3239 vdd.n1881 vss 0.00241f
C3240 vdd.n1882 vss 0.0141f
C3241 vdd.n1883 vss 0.00241f
C3242 vdd.n1884 vss 0.00271f
C3243 vdd.n1885 vss 0.00248f
C3244 vdd.n1886 vss 0.413f
C3245 vdd.n1887 vss 0.00248f
C3246 vdd.n1888 vss 0.00241f
C3247 vdd.n1889 vss 0.00821f
C3248 vdd.n1890 vss 0.00368f
C3249 vdd.n1891 vss 0.00394f
C3250 vdd.n1892 vss 0.00851f
C3251 vdd.n1893 vss 0.007f
C3252 vdd.n1894 vss 0.00311f
C3253 vdd.n1895 vss 0.00297f
C3254 vdd.n1896 vss 0.00241f
C3255 vdd.n1897 vss 0.00241f
C3256 vdd.n1898 vss 0.00248f
C3257 vdd.n1899 vss 0.00241f
C3258 vdd.n1900 vss 0.00821f
C3259 vdd.n1901 vss 0.00368f
C3260 vdd.n1902 vss -0.0674f
C3261 vdd.n1903 vss 0.00851f
C3262 vdd.n1904 vss 0.007f
C3263 vdd.n1905 vss 0.00311f
C3264 vdd.n1906 vss 0.00297f
C3265 vdd.n1907 vss 0.00241f
C3266 vdd.n1908 vss 0.00241f
C3267 vdd.n1909 vss 0.00248f
C3268 vdd.n1910 vss 0.00241f
C3269 vdd.n1911 vss 0.00821f
C3270 vdd.n1912 vss 0.00368f
C3271 vdd.n1913 vss 0.00394f
C3272 vdd.n1914 vss -0.174f
C3273 vdd.n1915 vss 0.007f
C3274 vdd.n1916 vss 0.00311f
C3275 vdd.n1917 vss 0.00297f
C3276 vdd.n1918 vss 0.00241f
C3277 vdd.n1919 vss 0.00241f
C3278 vdd.n1920 vss 0.00248f
C3279 vdd.n1921 vss 0.00241f
C3280 vdd.n1922 vss 0.00821f
C3281 vdd.n1923 vss 0.00368f
C3282 vdd.n1924 vss 0.00394f
C3283 vdd.n1925 vss 0.00851f
C3284 vdd.n1926 vss 0.007f
C3285 vdd.n1927 vss 0.00311f
C3286 vdd.n1928 vss 0.00297f
C3287 vdd.n1929 vss 0.00241f
C3288 vdd.n1930 vss 0.00241f
C3289 vdd.n1932 vss 0.00241f
C3290 vdd.n1933 vss 0.00856f
C3291 vdd.n1934 vss 0.00368f
C3292 vdd.n1935 vss -0.0674f
C3293 vdd.n1936 vss 0.00518f
C3294 vdd.n1937 vss 0.00394f
C3295 vdd.n1938 vss 0.00297f
C3296 vdd.n1939 vss 0.00241f
C3297 vdd.n1940 vss 4.25e-19
C3298 vdd.n1941 vss 0.00241f
C3299 vdd.n1942 vss 2.28f
C3300 vdd.n1943 vss 0.00248f
C3301 vdd.n1944 vss 0.00241f
C3302 vdd.n1945 vss 0.00821f
C3303 vdd.n1946 vss 0.00368f
C3304 vdd.n1947 vss 0.00394f
C3305 vdd.n1948 vss 0.007f
C3306 vdd.n1949 vss 0.0082f
C3307 vdd.n1950 vss 0.007f
C3308 vdd.n1951 vss 0.00311f
C3309 vdd.n1952 vss 0.00297f
C3310 vdd.n1953 vss 0.00241f
C3311 vdd.n1954 vss 0.00241f
C3312 vdd.n1955 vss 0.00877f
C3313 vdd.n1956 vss 0.00933f
C3314 vdd.n1957 vss 0.00241f
C3315 vdd.n1958 vss 0.00241f
C3316 vdd.n1959 vss 4.25e-19
C3317 vdd.n1960 vss 0.00877f
C3318 vdd.n1961 vss 0.00297f
C3319 vdd.n1962 vss 0.00594f
C3320 vdd.n1963 vss 0.00297f
C3321 vdd.n1964 vss 0.00722f
C3322 vdd.n1965 vss -0.0674f
C3323 vdd.n1966 vss 0.0082f
C3324 vdd.n1967 vss 0.00437f
C3325 vdd.n1968 vss -0.0772f
C3326 vdd.n1969 vss 2.92e-19
C3327 vdd.n1970 vss 4.25e-19
C3328 vdd.n1971 vss 0.00524f
C3329 vdd.n1972 vss 0.00311f
C3330 vdd.n1973 vss 0.00241f
C3331 vdd.n1974 vss 0.0115f
C3332 vdd.n1975 vss 0.00877f
C3333 vdd.n1976 vss 0.00297f
C3334 vdd.n1977 vss 0.00524f
C3335 vdd.n1978 vss 0.00311f
C3336 vdd.n1979 vss 4.25e-19
C3337 vdd.n1980 vss 2.92e-19
C3338 vdd.n1981 vss 0.00437f
C3339 vdd.n1982 vss 0.00836f
C3340 vdd.n1983 vss -0.0674f
C3341 vdd.n1984 vss 0.00368f
C3342 vdd.n1985 vss 0.00311f
C3343 vdd.n1986 vss 0.00821f
C3344 vdd.n1987 vss 0.00241f
C3345 vdd.n1988 vss 0.00877f
C3346 vdd.n1989 vss 0.00877f
C3347 vdd.n1990 vss 0.00241f
C3348 vdd.n1991 vss 0.00241f
C3349 vdd.n1992 vss 0.00241f
C3350 vdd.n1993 vss 0.00241f
C3351 vdd.n1994 vss 0.00311f
C3352 vdd.n1995 vss 0.00297f
C3353 vdd.n1996 vss 0.0255f
C3354 vdd.n1997 vss 0.00518f
C3355 vdd.n1998 vss 2.92e-19
C3356 vdd.n1999 vss 0.00297f
C3357 vdd.n2000 vss 0.00311f
C3358 vdd.n2001 vss 0.00821f
C3359 vdd.n2002 vss 0.00241f
C3360 vdd.n2003 vss 0.00241f
C3361 vdd.n2004 vss 0.0263f
C3362 vdd.n2005 vss 0.00297f
C3363 vdd.n2006 vss 0.0234f
C3364 vdd.n2007 vss 0.0256f
C3365 vdd.n2008 vss 0.0256f
C3366 vdd.n2009 vss 0.0234f
C3367 vdd.n2010 vss 0.00297f
C3368 vdd.n2011 vss 0.0263f
C3369 vdd.n2012 vss 0.00241f
C3370 vdd.n2014 vss 0.00241f
C3371 vdd.n2015 vss 0.00241f
C3372 vdd.n2016 vss 0.00311f
C3373 vdd.n2017 vss 0.00368f
C3374 vdd.n2018 vss 0.00335f
C3375 vdd.n2019 vss 0.00518f
C3376 vdd.n2020 vss 2.92e-19
C3377 vdd.n2021 vss 0.00297f
C3378 vdd.n2022 vss 0.00821f
C3379 vdd.n2023 vss 0.00241f
C3380 vdd.n2024 vss 0.00933f
C3381 vdd.n2025 vss 0.00241f
C3382 vdd.n2026 vss 0.00241f
C3383 vdd.n2027 vss 0.00311f
C3384 vdd.n2028 vss 0.00368f
C3385 vdd.n2029 vss 0.00335f
C3386 vdd.n2030 vss -0.0832f
C3387 vdd.n2031 vss 2.92e-19
C3388 vdd.n2032 vss 0.00297f
C3389 vdd.n2033 vss 0.00821f
C3390 vdd.n2034 vss 0.00877f
C3391 vdd.n2035 vss 0.00248f
C3392 vdd.n2036 vss 0.00241f
C3393 vdd.n2037 vss 0.00241f
C3394 vdd.n2038 vss 0.00821f
C3395 vdd.n2039 vss 4.25e-19
C3396 vdd.n2040 vss 0.00877f
C3397 vdd.n2041 vss 0.00297f
C3398 vdd.n2042 vss 0.00368f
C3399 vdd.n2043 vss 0.00335f
C3400 vdd.n2044 vss 0.00518f
C3401 vdd.n2045 vss -0.189f
C3402 vdd.n2046 vss 0.00502f
C3403 vdd.n2047 vss 0.00311f
C3404 vdd.n2048 vss 0.00241f
C3405 vdd.n2049 vss 0.00241f
C3406 vdd.n2050 vss 0.00248f
C3407 vdd.n2051 vss 0.00241f
C3408 vdd.n2052 vss 0.00821f
C3409 vdd.n2053 vss 0.00297f
C3410 vdd.n2054 vss 2.92e-19
C3411 vdd.n2055 vss 0.00335f
C3412 vdd.n2056 vss 0.0082f
C3413 vdd.n2057 vss 0.00335f
C3414 vdd.n2058 vss 0.00311f
C3415 vdd.n2059 vss 0.00241f
C3416 vdd.n2060 vss 0.00241f
C3417 vdd.n2061 vss 0.00248f
C3418 vdd.n2062 vss 0.00241f
C3419 vdd.n2063 vss 0.0265f
C3420 vdd.n2064 vss 0.00297f
C3421 vdd.n2065 vss 2.92e-19
C3422 vdd.n2066 vss 0.00518f
C3423 vdd.n2067 vss 0.0216f
C3424 vdd.n2068 vss 0.00368f
C3425 vdd.n2069 vss 0.00394f
C3426 vdd.n2070 vss -0.175f
C3427 vdd.n2071 vss 0.007f
C3428 vdd.n2072 vss 0.00311f
C3429 vdd.n2073 vss 0.00297f
C3430 vdd.n2074 vss 0.00241f
C3431 vdd.n2075 vss 0.0265f
C3432 vdd.n2076 vss 0.00241f
C3433 vdd.n2077 vss 0.00241f
C3434 vdd.n2078 vss 0.00248f
C3435 vdd.n2079 vss 0.00241f
C3436 vdd.n2080 vss 0.00821f
C3437 vdd.n2081 vss 0.00368f
C3438 vdd.n2082 vss 0.00394f
C3439 vdd.n2083 vss 0.0082f
C3440 vdd.n2084 vss 0.007f
C3441 vdd.n2085 vss 0.00311f
C3442 vdd.n2086 vss 0.00297f
C3443 vdd.n2087 vss 0.00241f
C3444 vdd.n2088 vss 0.00241f
C3445 vdd.n2089 vss 0.00877f
C3446 vdd.n2090 vss 0.00933f
C3447 vdd.n2091 vss 0.00241f
C3448 vdd.n2092 vss 0.00241f
C3449 vdd.n2093 vss 4.25e-19
C3450 vdd.n2094 vss 0.00877f
C3451 vdd.n2095 vss 0.00297f
C3452 vdd.n2096 vss 0.00594f
C3453 vdd.n2097 vss 0.00297f
C3454 vdd.n2098 vss 0.00722f
C3455 vdd.n2099 vss -0.0674f
C3456 vdd.n2100 vss 0.0082f
C3457 vdd.n2101 vss 0.00437f
C3458 vdd.n2102 vss -0.0772f
C3459 vdd.n2103 vss 2.92e-19
C3460 vdd.n2104 vss 4.25e-19
C3461 vdd.n2105 vss 0.00524f
C3462 vdd.n2106 vss 0.00311f
C3463 vdd.n2107 vss 0.00241f
C3464 vdd.n2108 vss 0.0115f
C3465 vdd.n2109 vss 0.00877f
C3466 vdd.n2110 vss 0.00297f
C3467 vdd.n2111 vss 0.00524f
C3468 vdd.n2112 vss 0.00311f
C3469 vdd.n2113 vss 4.25e-19
C3470 vdd.n2114 vss 2.92e-19
C3471 vdd.n2115 vss 0.00437f
C3472 vdd.n2116 vss 0.00836f
C3473 vdd.n2117 vss -0.0674f
C3474 vdd.n2118 vss 0.00368f
C3475 vdd.n2119 vss 0.00311f
C3476 vdd.n2120 vss 0.00821f
C3477 vdd.n2121 vss 0.00241f
C3478 vdd.n2122 vss 0.00877f
C3479 vdd.n2123 vss 0.00877f
C3480 vdd.n2124 vss 0.00241f
C3481 vdd.n2125 vss 0.00241f
C3482 vdd.n2126 vss 0.00241f
C3483 vdd.n2127 vss 0.00241f
C3484 vdd.n2128 vss 0.00311f
C3485 vdd.n2129 vss 0.00297f
C3486 vdd.n2130 vss 0.0255f
C3487 vdd.n2131 vss 0.00518f
C3488 vdd.n2132 vss 2.92e-19
C3489 vdd.n2133 vss 0.00297f
C3490 vdd.n2134 vss 0.00311f
C3491 vdd.n2135 vss 0.00821f
C3492 vdd.n2136 vss 0.00241f
C3493 vdd.n2137 vss 0.00241f
C3494 vdd.n2138 vss 0.0263f
C3495 vdd.n2139 vss 0.00297f
C3496 vdd.n2140 vss 0.0234f
C3497 vdd.n2141 vss 0.0256f
C3498 vdd.n2142 vss 0.0256f
C3499 vdd.n2143 vss 0.0234f
C3500 vdd.n2144 vss 0.00297f
C3501 vdd.n2145 vss 0.0263f
C3502 vdd.n2146 vss 0.00241f
C3503 vdd.n2148 vss 0.00241f
C3504 vdd.n2149 vss 0.00241f
C3505 vdd.n2150 vss 0.00311f
C3506 vdd.n2151 vss 0.00368f
C3507 vdd.n2152 vss 0.00335f
C3508 vdd.n2153 vss 0.00518f
C3509 vdd.n2154 vss 2.92e-19
C3510 vdd.n2155 vss 0.00297f
C3511 vdd.n2156 vss 0.00821f
C3512 vdd.n2157 vss 0.00241f
C3513 vdd.n2158 vss 0.00933f
C3514 vdd.n2159 vss 0.00241f
C3515 vdd.n2160 vss 0.00241f
C3516 vdd.n2161 vss 0.00311f
C3517 vdd.n2162 vss 0.00368f
C3518 vdd.n2163 vss 0.00335f
C3519 vdd.n2164 vss -0.0832f
C3520 vdd.n2165 vss 2.92e-19
C3521 vdd.n2166 vss 0.00297f
C3522 vdd.n2167 vss 0.00821f
C3523 vdd.n2168 vss 0.00877f
C3524 vdd.n2169 vss 0.00248f
C3525 vdd.n2170 vss 0.00241f
C3526 vdd.n2171 vss 0.00241f
C3527 vdd.n2172 vss 0.00821f
C3528 vdd.n2173 vss 4.25e-19
C3529 vdd.n2174 vss 0.00877f
C3530 vdd.n2175 vss 0.00297f
C3531 vdd.n2176 vss 0.00368f
C3532 vdd.n2177 vss 0.00335f
C3533 vdd.n2178 vss 0.00518f
C3534 vdd.n2179 vss -0.189f
C3535 vdd.n2180 vss 0.00502f
C3536 vdd.n2181 vss 0.00311f
C3537 vdd.n2182 vss 0.00241f
C3538 vdd.n2183 vss 0.00241f
C3539 vdd.n2184 vss 0.00248f
C3540 vdd.n2185 vss 0.00241f
C3541 vdd.n2186 vss 0.00821f
C3542 vdd.n2187 vss 0.00297f
C3543 vdd.n2188 vss 2.92e-19
C3544 vdd.n2189 vss 0.00335f
C3545 vdd.n2190 vss 0.0082f
C3546 vdd.n2191 vss 0.00335f
C3547 vdd.n2192 vss 0.00311f
C3548 vdd.n2193 vss 0.00241f
C3549 vdd.n2194 vss 0.00241f
C3550 vdd.n2195 vss 0.00248f
C3551 vdd.n2196 vss 0.00241f
C3552 vdd.n2197 vss 0.0265f
C3553 vdd.n2198 vss 0.00297f
C3554 vdd.n2199 vss 2.92e-19
C3555 vdd.n2200 vss 0.00518f
C3556 vdd.n2201 vss 0.0216f
C3557 vdd.n2202 vss 0.00368f
C3558 vdd.n2203 vss 0.00394f
C3559 vdd.n2204 vss -0.175f
C3560 vdd.n2205 vss 0.007f
C3561 vdd.n2206 vss 0.00311f
C3562 vdd.n2207 vss 0.00297f
C3563 vdd.n2208 vss 0.00241f
C3564 vdd.n2209 vss 0.0265f
C3565 vdd.n2210 vss 0.00241f
C3566 vdd.n2211 vss 0.00241f
C3567 vdd.n2212 vss 0.00248f
C3568 vdd.n2213 vss 0.00241f
C3569 vdd.n2214 vss 0.00821f
C3570 vdd.n2215 vss 0.00368f
C3571 vdd.n2216 vss 0.00394f
C3572 vdd.n2217 vss 0.0082f
C3573 vdd.n2218 vss 0.007f
C3574 vdd.n2219 vss 0.00311f
C3575 vdd.n2220 vss 0.00297f
C3576 vdd.n2221 vss 0.00241f
C3577 vdd.n2222 vss 0.00241f
C3578 vdd.n2223 vss 0.00877f
C3579 vdd.n2224 vss 0.00933f
C3580 vdd.n2225 vss 0.00241f
C3581 vdd.n2226 vss 0.00241f
C3582 vdd.n2227 vss 4.25e-19
C3583 vdd.n2228 vss 0.00877f
C3584 vdd.n2229 vss 0.00297f
C3585 vdd.n2230 vss 0.00594f
C3586 vdd.n2231 vss 0.00297f
C3587 vdd.n2232 vss 0.00722f
C3588 vdd.n2233 vss -0.0674f
C3589 vdd.n2234 vss 0.0082f
C3590 vdd.n2235 vss 0.00437f
C3591 vdd.n2236 vss -0.0772f
C3592 vdd.n2237 vss 2.92e-19
C3593 vdd.n2238 vss 4.25e-19
C3594 vdd.n2239 vss 0.00524f
C3595 vdd.n2240 vss 0.00311f
C3596 vdd.n2241 vss 0.00241f
C3597 vdd.n2242 vss 0.0115f
C3598 vdd.n2243 vss 0.00877f
C3599 vdd.n2244 vss 0.00297f
C3600 vdd.n2245 vss 0.00524f
C3601 vdd.n2246 vss 0.00311f
C3602 vdd.n2247 vss 4.25e-19
C3603 vdd.n2248 vss 2.92e-19
C3604 vdd.n2249 vss 0.00437f
C3605 vdd.n2250 vss 0.00836f
C3606 vdd.n2251 vss -0.0674f
C3607 vdd.n2252 vss 0.00368f
C3608 vdd.n2253 vss 0.00311f
C3609 vdd.n2254 vss 0.00821f
C3610 vdd.n2255 vss 0.00241f
C3611 vdd.n2256 vss 0.00877f
C3612 vdd.n2257 vss 0.00877f
C3613 vdd.n2258 vss 0.00241f
C3614 vdd.n2259 vss 0.00241f
C3615 vdd.n2260 vss 0.00241f
C3616 vdd.n2261 vss 0.00241f
C3617 vdd.n2262 vss 0.00311f
C3618 vdd.n2263 vss 0.00297f
C3619 vdd.n2264 vss 0.0255f
C3620 vdd.n2265 vss 0.00518f
C3621 vdd.n2266 vss 2.92e-19
C3622 vdd.n2267 vss 0.00297f
C3623 vdd.n2268 vss 0.00311f
C3624 vdd.n2269 vss 0.00821f
C3625 vdd.n2270 vss 0.00241f
C3626 vdd.n2271 vss 0.00241f
C3627 vdd.n2272 vss 0.0263f
C3628 vdd.n2273 vss 0.00297f
C3629 vdd.n2274 vss 0.0234f
C3630 vdd.n2275 vss 0.0256f
C3631 vdd.n2276 vss 0.0256f
C3632 vdd.n2277 vss 0.0234f
C3633 vdd.n2278 vss 0.00297f
C3634 vdd.n2279 vss 0.0263f
C3635 vdd.n2280 vss 0.00241f
C3636 vdd.n2282 vss 0.00241f
C3637 vdd.n2283 vss 0.00241f
C3638 vdd.n2284 vss 0.00311f
C3639 vdd.n2285 vss 0.00368f
C3640 vdd.n2286 vss 0.00335f
C3641 vdd.n2287 vss 0.00518f
C3642 vdd.n2288 vss 2.92e-19
C3643 vdd.n2289 vss 0.00297f
C3644 vdd.n2290 vss 0.00821f
C3645 vdd.n2291 vss 0.00241f
C3646 vdd.n2292 vss 0.00933f
C3647 vdd.n2293 vss 0.00241f
C3648 vdd.n2294 vss 0.00241f
C3649 vdd.n2295 vss 0.00311f
C3650 vdd.n2296 vss 0.00368f
C3651 vdd.n2297 vss 0.00335f
C3652 vdd.n2298 vss -0.0832f
C3653 vdd.n2299 vss 2.92e-19
C3654 vdd.n2300 vss 0.00297f
C3655 vdd.n2301 vss 0.00821f
C3656 vdd.n2302 vss 0.00877f
C3657 vdd.n2303 vss 0.00248f
C3658 vdd.n2304 vss 0.00241f
C3659 vdd.n2305 vss 0.00241f
C3660 vdd.n2306 vss 0.00821f
C3661 vdd.n2307 vss 4.25e-19
C3662 vdd.n2308 vss 0.00877f
C3663 vdd.n2309 vss 0.00297f
C3664 vdd.n2310 vss 0.00368f
C3665 vdd.n2311 vss 0.00335f
C3666 vdd.n2312 vss 0.00518f
C3667 vdd.n2313 vss -0.189f
C3668 vdd.n2314 vss 0.00502f
C3669 vdd.n2315 vss 0.00311f
C3670 vdd.n2316 vss 0.00241f
C3671 vdd.n2317 vss 0.00241f
C3672 vdd.n2318 vss 0.00248f
C3673 vdd.n2319 vss 0.00241f
C3674 vdd.n2320 vss 0.00821f
C3675 vdd.n2321 vss 0.00297f
C3676 vdd.n2322 vss 2.92e-19
C3677 vdd.n2323 vss 0.00335f
C3678 vdd.n2324 vss 0.0082f
C3679 vdd.n2325 vss 0.00335f
C3680 vdd.n2326 vss 0.00311f
C3681 vdd.n2327 vss 0.00241f
C3682 vdd.n2328 vss 0.00241f
C3683 vdd.n2329 vss 0.00248f
C3684 vdd.n2330 vss 0.00241f
C3685 vdd.n2331 vss 0.0265f
C3686 vdd.n2332 vss 0.00297f
C3687 vdd.n2333 vss 2.92e-19
C3688 vdd.n2334 vss 0.00518f
C3689 vdd.n2335 vss 0.0216f
C3690 vdd.n2336 vss 0.00368f
C3691 vdd.n2337 vss 0.00394f
C3692 vdd.n2338 vss -0.175f
C3693 vdd.n2339 vss 0.007f
C3694 vdd.n2340 vss 0.00311f
C3695 vdd.n2341 vss 0.00297f
C3696 vdd.n2342 vss 0.00241f
C3697 vdd.n2343 vss 0.0265f
C3698 vdd.n2344 vss 0.00241f
C3699 vdd.n2345 vss 0.00241f
C3700 vdd.n2346 vss 0.00248f
C3701 vdd.n2347 vss 0.00241f
C3702 vdd.n2348 vss 0.00821f
C3703 vdd.n2349 vss 0.00368f
C3704 vdd.n2350 vss 0.00394f
C3705 vdd.n2351 vss 0.0082f
C3706 vdd.n2352 vss 0.007f
C3707 vdd.n2353 vss 0.00311f
C3708 vdd.n2354 vss 0.00297f
C3709 vdd.n2355 vss 0.00241f
C3710 vdd.n2356 vss 0.00241f
C3711 vdd.n2357 vss 0.00877f
C3712 vdd.n2358 vss 0.00933f
C3713 vdd.n2359 vss 0.00241f
C3714 vdd.n2360 vss 0.00241f
C3715 vdd.n2361 vss 4.25e-19
C3716 vdd.n2362 vss 0.00877f
C3717 vdd.n2363 vss 0.00297f
C3718 vdd.n2364 vss 0.00594f
C3719 vdd.n2365 vss 0.00297f
C3720 vdd.n2366 vss 0.00722f
C3721 vdd.n2367 vss -0.0674f
C3722 vdd.n2368 vss 0.0082f
C3723 vdd.n2369 vss 0.00437f
C3724 vdd.n2370 vss -0.0772f
C3725 vdd.n2371 vss 2.92e-19
C3726 vdd.n2372 vss 4.25e-19
C3727 vdd.n2373 vss 0.00524f
C3728 vdd.n2374 vss 0.00311f
C3729 vdd.n2375 vss 0.00241f
C3730 vdd.n2376 vss 0.0115f
C3731 vdd.n2377 vss 0.00877f
C3732 vdd.n2378 vss 0.00297f
C3733 vdd.n2379 vss 0.00524f
C3734 vdd.n2380 vss 0.00311f
C3735 vdd.n2381 vss 4.25e-19
C3736 vdd.n2382 vss 2.92e-19
C3737 vdd.n2383 vss 0.00437f
C3738 vdd.n2384 vss 0.00836f
C3739 vdd.n2385 vss -0.0674f
C3740 vdd.n2386 vss 0.00368f
C3741 vdd.n2387 vss 0.00311f
C3742 vdd.n2388 vss 0.00821f
C3743 vdd.n2389 vss 0.00241f
C3744 vdd.n2390 vss 0.00877f
C3745 vdd.n2391 vss 0.00877f
C3746 vdd.n2392 vss 0.00241f
C3747 vdd.n2393 vss 0.00241f
C3748 vdd.n2394 vss 0.00241f
C3749 vdd.n2395 vss 0.00241f
C3750 vdd.n2396 vss 0.00311f
C3751 vdd.n2397 vss 0.00297f
C3752 vdd.n2398 vss 0.0255f
C3753 vdd.n2399 vss 0.00518f
C3754 vdd.n2400 vss 2.92e-19
C3755 vdd.n2401 vss 0.00297f
C3756 vdd.n2402 vss 0.00311f
C3757 vdd.n2403 vss 0.00821f
C3758 vdd.n2404 vss 0.00241f
C3759 vdd.n2405 vss 0.00241f
C3760 vdd.n2406 vss 0.0263f
C3761 vdd.n2407 vss 0.00297f
C3762 vdd.n2408 vss 0.0234f
C3763 vdd.n2409 vss 0.0256f
C3764 vdd.n2410 vss 0.0256f
C3765 vdd.n2411 vss 0.0234f
C3766 vdd.n2412 vss 0.00297f
C3767 vdd.n2413 vss 0.0263f
C3768 vdd.n2414 vss 0.00241f
C3769 vdd.n2416 vss 0.00241f
C3770 vdd.n2417 vss 0.00241f
C3771 vdd.n2418 vss 0.00311f
C3772 vdd.n2419 vss 0.00368f
C3773 vdd.n2420 vss 0.00335f
C3774 vdd.n2421 vss 0.00518f
C3775 vdd.n2422 vss 2.92e-19
C3776 vdd.n2423 vss 0.00297f
C3777 vdd.n2424 vss 0.00821f
C3778 vdd.n2425 vss 0.00241f
C3779 vdd.n2426 vss 0.00933f
C3780 vdd.n2427 vss 0.00241f
C3781 vdd.n2428 vss 0.00241f
C3782 vdd.n2429 vss 0.00311f
C3783 vdd.n2430 vss 0.00368f
C3784 vdd.n2431 vss 0.00335f
C3785 vdd.n2432 vss -0.0832f
C3786 vdd.n2433 vss 2.92e-19
C3787 vdd.n2434 vss 0.00297f
C3788 vdd.n2435 vss 0.00821f
C3789 vdd.n2436 vss 0.00877f
C3790 vdd.n2437 vss 0.00248f
C3791 vdd.n2438 vss 0.00241f
C3792 vdd.n2439 vss 0.00241f
C3793 vdd.n2440 vss 0.00821f
C3794 vdd.n2441 vss 4.25e-19
C3795 vdd.n2442 vss 0.00877f
C3796 vdd.n2443 vss 0.00297f
C3797 vdd.n2444 vss 0.00368f
C3798 vdd.n2445 vss 0.00335f
C3799 vdd.n2446 vss 0.00518f
C3800 vdd.n2447 vss -0.189f
C3801 vdd.n2448 vss 0.00502f
C3802 vdd.n2449 vss 0.00311f
C3803 vdd.n2450 vss 0.00241f
C3804 vdd.n2451 vss 0.00241f
C3805 vdd.n2453 vss 0.00241f
C3806 vdd.n2454 vss 0.00821f
C3807 vdd.n2455 vss 0.00297f
C3808 vdd.n2456 vss 2.92e-19
C3809 vdd.n2457 vss 0.00335f
C3810 vdd.n2458 vss 0.0082f
C3811 vdd.n2459 vss 0.00335f
C3812 vdd.n2460 vss 0.00311f
C3813 vdd.n2461 vss 0.00241f
C3814 vdd.n2462 vss 0.00241f
C3815 vdd.n2463 vss 0.0349f
C3816 vdd.n2464 vss 0.00297f
C3817 vdd.n2465 vss 2.92e-19
C3818 vdd.n2466 vss 0.072f
C3819 vdd.n2467 vss 0.0396f
C3820 vdd.n2468 vss 0.0178f
C3821 vdd.n2469 vss 0.0839f
C3822 vdd.n2470 vss 0.00568f
C3823 vdd.t87 vss 2.02f
C3824 vdd.n2471 vss 0.00744f
C3825 vdd.n2472 vss 0.0179f
C3826 vdd.n2473 vss 0.0178f
C3827 vdd.n2474 vss 0.0396f
C3828 vdd.n2475 vss 0.0178f
C3829 vdd.n2476 vss 0.00568f
C3830 vdd.n2477 vss 0.0179f
C3831 vdd.n2478 vss 0.15f
C3832 vdd.n2479 vss 0.0178f
C3833 vdd.n2480 vss 0.00568f
C3834 vdd.t0 vss 0.226f
C3835 vdd.n2481 vss 0.0155f
C3836 vdd.n2482 vss 0.00912f
C3837 vdd.t1 vss 0.00523f
C3838 vdd.n2483 vss 0.0323f
C3839 vdd.n2484 vss 0.0519f
C3840 vdd.n2485 vss 0.0567f
C3841 vdd.n2486 vss 0.00744f
C3842 vdd.n2487 vss 0.00733f
C3843 vdd.n2488 vss 0.0728f
C3844 vdd.n2489 vss 1.81f
C3845 vdd.n2490 vss 0.275f
C3846 vdd.t61 vss 1.49f
C3847 vdd.n2491 vss 0.422f
C3848 vdd.n2492 vss 0.00744f
C3849 vdd.n2493 vss 0.0728f
C3850 vdd.n2494 vss 0.00733f
C3851 vdd.n2495 vss 0.0179f
C3852 vdd.n2496 vss 0.00988f
C3853 vdd.n2497 vss 0.0618f
C3854 vdd.n2498 vss 0.0887f
C3855 vdd.n2499 vss 0.00973f
C3856 vdd.n2500 vss 0.0806f
C3857 vdd.n2501 vss 0.0396f
C3858 vdd.n2502 vss 0.0806f
C3859 vdd.n2503 vss 0.00973f
C3860 vdd.n2504 vss 0.00568f
C3861 vdd.n2505 vss 0.00733f
C3862 vdd.n2506 vss 0.0728f
C3863 vdd.n2507 vss 1.86f
C3864 vdd.t10 vss 2.26f
C3865 vdd.n2508 vss 0.0397f
C3866 vdd.n2509 vss 0.00744f
C3867 vdd.n2510 vss 0.0179f
C3868 vdd.n2511 vss 0.0178f
C3869 vdd.n2512 vss 0.0368f
C3870 vdd.n2513 vss 0.00973f
C3871 vdd.n2514 vss 0.00503f
C3872 vdd.n2515 vss 0.0309f
C3873 vdd.n2516 vss 0.0594f
C3874 vdd.n2517 vss 0.0298f
C3875 vdd.t35 vss 0.0456f
C3876 vdd.n2518 vss 0.0771f
C3877 vdd.n2519 vss 0.0381f
C3878 vdd.n2520 vss 0.0188f
C3879 vdd.n2521 vss 0.00752f
C3880 vdd.n2522 vss 0.0275f
C3881 vdd.n2523 vss 0.0287f
C3882 vdd.t30 vss 0.0322f
C3883 vdd.n2524 vss 0.0457f
C3884 vdd.n2525 vss 0.0408f
C3885 vdd.n2526 vss 0.0531f
C3886 vdd.n2527 vss 0.0351f
C3887 vdd.t25 vss 0.0113f
C3888 vdd.t13 vss -0.00623f
C3889 vdd.n2528 vss 0.0441f
C3890 vdd.n2529 vss 0.0348f
C3891 vdd.n2530 vss 0.0538f
C3892 vdd.n2531 vss 0.0232f
C3893 vdd.n2532 vss 0.0312f
C3894 vdd.n2533 vss 0.0281f
C3895 vdd.t24 vss 0.466f
C3896 vdd.t12 vss 0.0903f
C3897 vdd.t29 vss 0.0376f
C3898 vdd.t14 vss 0.376f
C3899 vdd.n2534 vss 0.37f
C3900 vdd.n2535 vss 0.00376f
C3901 vdd.n2536 vss 0.024f
C3902 vdd.t15 vss 0.0104f
C3903 vdd.t50 vss -0.00332f
C3904 vdd.n2537 vss 0.048f
C3905 vdd.n2538 vss 0.049f
C3906 vdd.n2539 vss 0.0202f
C3907 vdd.n2540 vss 0.0168f
C3908 vdd.n2541 vss 0.142f
C3909 vdd.n2542 vss 0.142f
C3910 vdd.n2543 vss 0.0368f
C3911 vdd.n2544 vss 0.00949f
C3912 vdd.n2545 vss 0.0368f
C3913 vdd.n2546 vss 0.00949f
C3914 vdd.n2547 vss 0.0168f
C3915 vdd.n2548 vss 0.0535f
C3916 vdd.t72 vss 0.00949f
C3917 vdd.t5 vss 0.00309f
C3918 vdd.n2549 vss 0.0486f
C3919 vdd.n2550 vss 0.0672f
C3920 vdd.n2551 vss 0.0276f
C3921 vdd.t26 vss 0.141f
C3922 vdd.n2552 vss 0.0284f
C3923 vdd.n2553 vss 0.0408f
C3924 vdd.n2554 vss 0.035f
C3925 vdd.n2555 vss 0.0535f
C3926 vdd.n2556 vss 0.00268f
C3927 vdd.n2557 vss 0.0476f
C3928 vdd.n2558 vss 0.0168f
C3929 vdd.n2559 vss 0.215f
C3930 vdd.n2560 vss 0.215f
C3931 vdd.n2561 vss 0.0535f
C3932 vdd.n2562 vss 0.0408f
C3933 vdd.n2563 vss 0.00313f
C3934 vdd.n2564 vss 0.0279f
C3935 vdd.n2565 vss 0.0284f
C3936 vdd.t85 vss 0.0303f
C3937 vdd.n2566 vss 0.0261f
C3938 vdd.t7 vss 0.00666f
C3939 vdd.t86 vss 0.00702f
C3940 vdd.n2567 vss 0.0143f
C3941 vdd.n2568 vss 0.0637f
C3942 vdd.n2569 vss 0.0321f
C3943 vdd.n2570 vss 0.0379f
C3944 vdd.n2571 vss 0.0417f
C3945 vdd.n2572 vss 0.0505f
C3946 vdd.t18 vss 0.144f
C3947 vdd.n2573 vss 0.0272f
C3948 vdd.t60 vss 0.00522f
C3949 vdd.t3 vss 0.00666f
C3950 vdd.n2574 vss 0.0137f
C3951 vdd.n2575 vss 0.0616f
C3952 vdd.n2576 vss 0.0379f
C3953 vdd.t58 vss 0.0171f
C3954 vdd.n2577 vss 0.0899f
C3955 vdd.n2578 vss 0.0421f
C3956 vdd.t39 vss 0.00741f
C3957 vdd.t19 vss 0.00741f
C3958 vdd.n2579 vss 0.0157f
C3959 vdd.t59 vss 0.0735f
C3960 vdd.n2580 vss 0.0735f
C3961 vdd.t38 vss 0.109f
C3962 vdd.n2581 vss 0.0272f
C3963 vdd.n2582 vss 0.0269f
C3964 vdd.n2583 vss 0.00806f
C3965 vdd.n2584 vss 0.0323f
C3966 vdd.n2585 vss 0.0301f
C3967 vdd.n2586 vss 0.0748f
C3968 vdd.n2587 vss 0.0215f
C3969 vdd.n2588 vss 0.0748f
C3970 vdd.n2589 vss 0.0379f
C3971 vdd.n2590 vss 0.012f
C3972 vdd.t96 vss 0.0108f
C3973 vdd.n2591 vss 0.0316f
C3974 vdd.t56 vss 0.0285f
C3975 vdd.n2592 vss 0.0566f
C3976 vdd.n2593 vss 0.0379f
C3977 vdd.n2594 vss 0.0379f
C3978 vdd.n2595 vss 0.0379f
C3979 vdd.n2596 vss 0.0379f
C3980 vdd.n2597 vss 0.0435f
C3981 vdd.n2598 vss 0.0412f
C3982 vdd.n2599 vss 0.0632f
C3983 vdd.n2600 vss 0.0379f
C3984 vdd.n2601 vss 0.0379f
C3985 vdd.n2602 vss 0.0379f
C3986 vdd.n2603 vss 0.0618f
C3987 vdd.n2604 vss 0.0494f
C3988 vdd.n2605 vss 0.0927f
C3989 vdd.t2 vss 0.125f
C3990 vdd.t31 vss 0.208f
C3991 vdd.t57 vss 0.241f
C3992 vdd.t75 vss 0.216f
C3993 vdd.n2606 vss 0.101f
C3994 vdd.t91 vss 0.0671f
C3995 vdd.t20 vss 0.123f
C3996 vdd.t92 vss 0.104f
C3997 vdd.n2607 vss 0.113f
C3998 vdd.t6 vss 0.102f
C3999 vdd.t36 vss 0.102f
C4000 vdd.n2608 vss 0.131f
C4001 vdd.n2609 vss 0.0282f
C4002 vdd.n2610 vss 0.0408f
C4003 vdd.n2611 vss 0.0408f
C4004 vdd.t37 vss 0.00949f
C4005 vdd.t93 vss 0.00309f
C4006 vdd.n2612 vss 0.0486f
C4007 vdd.n2613 vss 0.0399f
C4008 vdd.n2614 vss 0.00134f
C4009 vdd.n2615 vss 0.0321f
C4010 vdd.n2616 vss 0.395f
C4011 vdd.n2617 vss 0.0256f
C4012 vdd.n2618 vss 0.0435f
C4013 vdd.n2619 vss 0.0278f
C4014 vdd.n2620 vss 0.0272f
C4015 vdd.n2621 vss 0.161f
C4016 vdd.n2622 vss 0.166f
C4017 vdd.t82 vss 0.142f
C4018 vdd.n2623 vss 0.0367f
C4019 vdd.t74 vss 0.152f
C4020 vdd.t21 vss 0.144f
C4021 vdd.n2624 vss 0.15f
C4022 vdd.n2625 vss 0.0284f
C4023 vdd.n2626 vss 0.0408f
C4024 vdd.n2627 vss 0.0408f
C4025 vdd.n2628 vss 0.039f
C4026 vdd.n2629 vss 0.0535f
C4027 vdd.n2630 vss 0.0535f
C4028 vdd.t77 vss 0.00522f
C4029 vdd.t23 vss 0.00666f
C4030 vdd.n2631 vss 0.0137f
C4031 vdd.t28 vss 0.0119f
C4032 vdd.t9 vss 0.0267f
C4033 vdd.n2632 vss 0.0414f
C4034 vdd.n2633 vss 0.0197f
C4035 vdd.n2634 vss 0.058f
C4036 vdd.n2635 vss 0.041f
C4037 vdd.n2636 vss 0.0206f
C4038 vdd.n2637 vss 0.00134f
C4039 vdd.n2638 vss 0.0535f
C4040 vdd.n2639 vss 0.0535f
C4041 vdd.n2640 vss 0.0535f
C4042 vdd.n2641 vss 8.92e-19
C4043 vdd.n2642 vss 0.0408f
C4044 vdd.n2643 vss 0.0272f
C4045 vdd.n2644 vss 0.161f
C4046 vdd.t41 vss 0.0799f
C4047 vdd.t8 vss 0.115f
C4048 vdd.t22 vss 0.0687f
C4049 vdd.n2645 vss 0.153f
C4050 vdd.t76 vss 0.15f
C4051 vdd.t27 vss 0.0128f
C4052 vdd.n2646 vss 0.134f
C4053 vdd.n2647 vss 0.0278f
C4054 vdd.n2648 vss 0.0408f
C4055 vdd.n2649 vss 0.0385f
C4056 vdd.n2650 vss 0.00179f
C4057 vdd.n2651 vss 0.0116f
C4058 vdd.n2652 vss 0.0487f
C4059 vdd.n2653 vss 0.608f
C4060 vdd.n2654 vss 0.0368f
C4061 vdd.n2655 vss 0.00949f
C4062 vdd.n2656 vss 0.0181f
C4063 vdd.n2657 vss 0.0201f
C4064 vdd.n2658 vss 0.0529f
C4065 vdd.n2659 vss 0.00639f
C4066 vdd.n2660 vss 0.0535f
C4067 vdd.n2661 vss 0.0412f
C4068 vdd.n2662 vss 0.0412f
C4069 vdd.n2663 vss 0.00179f
C4070 vdd.n2664 vss 0.0535f
C4071 vdd.n2665 vss 0.0535f
C4072 vdd.t17 vss 0.00702f
C4073 vdd.t84 vss 0.00702f
C4074 vdd.n2666 vss 0.0145f
C4075 vdd.n2667 vss 0.0651f
C4076 vdd.n2668 vss 8.92e-19
C4077 vdd.n2669 vss 0.00672f
C4078 vdd.n2670 vss 0.0535f
C4079 vdd.n2671 vss 0.0535f
C4080 vdd.n2672 vss 0.0535f
C4081 vdd.n2673 vss 0.0399f
C4082 vdd.n2674 vss 0.027f
C4083 vdd.n2675 vss 0.152f
C4084 vdd.t16 vss 0.0431f
C4085 vdd.t71 vss 0.117f
C4086 vdd.n2676 vss 0.16f
C4087 vdd.t83 vss 0.0703f
C4088 vdd.t4 vss 0.0463f
C4089 vdd.n2677 vss 1.49f
C4090 vdd.t95 vss 0.134f
C4091 vdd.n2678 vss 0.107f
C4092 vdd.n2679 vss 0.0267f
C4093 vdd.n2680 vss 0.0408f
C4094 vdd.n2681 vss 0.0192f
C4095 vdd.n2682 vss 0.0253f
C4096 vdd.n2683 vss 0.0375f
C4097 vdd.n2684 vss 0.00174f
C4098 vdd.n2685 vss 0.00871f
C4099 vdd.n2686 vss 0.0201f
C4100 vdd.n2687 vss 0.0181f
C4101 vdd.n2688 vss 0.182f
C4102 vdd.n2689 vss 0.182f
C4103 vdd.n2690 vss 0.0168f
C4104 vdd.n2691 vss 0.0201f
C4105 vdd.n2692 vss 0.0181f
C4106 vdd.n2693 vss 0.148f
C4107 vdd.n2694 vss 0.148f
C4108 vdd.n2695 vss 0.0368f
C4109 vdd.n2696 vss 0.00949f
C4110 vdd.n2697 vss 0.0181f
C4111 vdd.n2698 vss 0.0201f
C4112 vdd.n2699 vss 0.0351f
C4113 vdd.n2700 vss 0.0275f
C4114 vdd.n2701 vss 0.0515f
C4115 vdd.n2702 vss 0.0527f
C4116 vdd.n2703 vss 0.0331f
C4117 vdd.n2704 vss 0.0242f
C4118 vdd.n2705 vss 0.0392f
C4119 vdd.n2707 vss 0.0327f
C4120 vdd.n2708 vss 0.0258f
C4121 vdd.n2709 vss 0.0211f
C4122 vdd.n2710 vss 0.0702f
C4123 vdd.n2711 vss 0.05f
C4124 vdd.n2712 vss 0.00443f
C4125 vdd.n2713 vss 0.0445f
C4126 vdd.n2714 vss 0.0408f
C4127 vdd.n2715 vss 0.0553f
C4128 vdd.n2716 vss 0.0702f
C4129 vdd.n2717 vss 0.0395f
C4130 vdd.n2718 vss 0.0142f
C4131 vdd.n2719 vss 0.0279f
C4132 vdd.n2720 vss 0.0094f
C4133 vdd.n2721 vss 0.0528f
C4134 vdd.n2722 vss 0.0138f
C4135 vdd.n2723 vss 0.0343f
C4136 vdd.n2724 vss 0.0492f
C4137 vdd.n2725 vss 0.0351f
C4138 vdd.n2726 vss 0.0201f
C4139 vdd.n2727 vss 0.00502f
C4140 vdd.n2728 vss 0.0963f
C4141 vdd.n2729 vss 0.0977f
C4142 vdd.n2730 vss 0.0173f
C4143 vdd.n2731 vss 0.0154f
C4144 vdd.n2732 vss 0.00704f
C4145 vdd.n2733 vss 0.0151f
C4146 vdd.n2734 vss 0.00594f
C4147 vdd.t33 vss 0.00594f
C4148 vdd.t34 vss 0.00594f
C4149 vdd.n2735 vss 0.0146f
C4150 vdd.n2736 vss 0.0432f
C4151 vdd.n2737 vss 0.00722f
C4152 vdd.n2738 vss 0.0147f
C4153 vdd.n2739 vss 0.0844f
C4154 vdd.n2740 vss 0.182f
C4155 vdd.n2741 vss 0.0178f
C4156 vdd.n2742 vss 0.0377f
C4157 vdd.t80 vss 0.0079f
C4158 vdd.n2743 vss 0.102f
C4159 vdd.n2744 vss 0.0179f
C4160 vdd.n2745 vss 0.00973f
C4161 vdd.n2746 vss 0.122f
C4162 vdd.n2747 vss 0.14f
C4163 vdd.n2748 vss 0.0396f
C4164 vdd.n2749 vss 0.0839f
C4165 vdd.n2750 vss 0.00973f
C4166 vdd.n2751 vss 0.00568f
C4167 vdd.n2752 vss 0.00733f
C4168 vdd.n2753 vss 0.0728f
C4169 vdd.t62 vss 0.384f
C4170 vdd.t11 vss 0.826f
C4171 vdd.n2754 vss 0.0145f
C4172 vdd.t32 vss 2f
C4173 vdd.t79 vss 5.97f
C4174 vdd.t55 vss 4.58f
C4175 vdd.n2755 vss 0.0281f
C4176 vdd.n2756 vss 0.0134f
C4177 vdd.n2757 vss 0.00146f
C4178 vdd.n2758 vss 0.00229f
C4179 vdd.n2759 vss 0.00229f
C4180 vdd.n2760 vss 0.0035f
C4181 vdd.n2761 vss 0.00782f
C4182 vdd.n2762 vss 0.00397f
C4183 vdd.n2763 vss 0.00602f
C4184 vdd.n2764 vss 0.0179f
C4185 vdd.n2765 vss 0.0245f
C4186 vdd.t54 vss 0.0456f
C4187 vdd.n2766 vss 0.0245f
C4188 vdd.n2767 vss 0.0543f
C4189 vdd.n2768 vss 0.0234f
C4190 vdd.n2769 vss 7.3e-19
C4191 vdd.n2770 vss 0.0177f
C4192 vdd.n2771 vss 0.0154f
C4193 vdd.n2772 vss 0.0502f
C4194 vdd.n2773 vss 0.00714f
C4195 vdd.n2774 vss 0.00954f
C4196 vdd.n2775 vss 0.0098f
C4197 vdd.n2776 vss 0.0035f
C4198 vdd.n2777 vss 0.0165f
C4199 vdd.n2778 vss 0.00365f
C4200 vdd.n2779 vss 0.00618f
C4201 vdd.n2780 vss 0.00991f
C4202 vdd.n2781 vss 0.00618f
C4203 vdd.n2782 vss 7.3e-19
C4204 vdd.n2783 vss 0.0167f
C4205 vdd.n2784 vss 0.0153f
C4206 vdd.n2785 vss 0.0208f
C4207 vdd.n2786 vss 0.0367f
C4208 vdd.n2787 vss 0.0191f
C4209 vdd.t67 vss 0.0456f
C4210 vdd.n2788 vss 0.00886f
C4211 vdd.n2789 vss 0.00968f
C4212 vdd.n2790 vss 0.0112f
C4213 vdd.n2791 vss 0.0677f
C4214 vdd.t66 vss 0.0921f
C4215 vdd.n2792 vss 0.0834f
C4216 vdd.n2793 vss 0.0181f
C4217 vdd.n2794 vss 0.00714f
C4218 vdd.n2795 vss 0.0498f
C4219 vdd.n2796 vss 0.0201f
C4220 vdd.n2797 vss 0.0189f
C4221 vdd.n2798 vss 0.0177f
C4222 vdd.n2799 vss 0.0143f
C4223 vdd.n2800 vss 0.0118f
C4224 vdd.n2801 vss 0.0043f
C4225 vdd.n2802 vss 0.0111f
C4226 vdd.n2803 vss 0.00413f
C4227 vdd.n2804 vss 0.00432f
C4228 vdd.n2805 vss 0.00165f
C4229 vdd.n2806 vss 0.00121f
C4230 vdd.n2807 vss 0.0125f
C4231 vdd.n2808 vss 0.0818f
C4232 vdd.t53 vss 0.112f
C4233 vdd.n2809 vss 0.0567f
C4234 vdd.n2810 vss 0.819f
C4235 vdd.n2811 vss 0.355f
C4236 vdd.n2812 vss 1.24f
C4237 vdd.t70 vss 2.06f
C4238 vdd.n2813 vss 1.86f
C4239 vdd.n2814 vss 0.00744f
C4240 vdd.n2815 vss 0.0728f
C4241 vdd.n2816 vss 0.00733f
C4242 vdd.n2817 vss 0.0179f
C4243 vdd.n2818 vss 0.00973f
C4244 vdd.n2819 vss 0.0403f
C4245 vdd.n2820 vss 0.106f
C4246 vdd.n2821 vss 0.0052f
C4247 vdd.n2822 vss 0.0357f
C4248 vdd.n2823 vss 0.00394f
C4249 vdd.n2824 vss 0.00502f
C4250 vdd.n2825 vss -0.0832f
C4251 vdd.n2826 vss -0.168f
C4252 vdd.n2827 vss 0.00714f
C4253 vdd.n2828 vss 0.00437f
C4254 vdd.n2829 vss 4.25e-19
C4255 vdd.n2830 vss 0.0378f
C4256 vdd.n2831 vss 0.0462f
C4257 vdd.n2832 vss 0.0181f
C4258 vdd.n2833 vss 0.00248f
C4259 vdd.n2834 vss 0.0115f
C4260 vdd.n2835 vss 0.00877f
C4261 vdd.n2836 vss 0.00877f
C4262 vdd.n2837 vss 0.00297f
C4263 vdd.n2838 vss 0.00594f
C4264 vdd.n2839 vss 0.00722f
C4265 vdd.n2840 vss 0.00368f
C4266 vdd.n2841 vss 0.00524f
C4267 vdd.n2842 vss 0.00423f
C4268 vdd.n2843 vss 0.00394f
C4269 vdd.n2844 vss 0.00502f
C4270 vdd.n2845 vss 0.00518f
C4271 vdd.n2846 vss 0.0082f
C4272 vdd.n2847 vss 0.00836f
C4273 vdd.n2848 vss 0.00714f
C4274 vdd.n2849 vss 0.00437f
C4275 vdd.n2850 vss 4.25e-19
C4276 vdd.n2851 vss 0.00311f
C4277 vdd.n2852 vss 2.83e-19
C4278 vdd.n2853 vss 0.00933f
C4279 vdd.n2855 vss 0.0115f
C4280 vdd.n2856 vss 0.00877f
C4281 vdd.n2857 vss 0.00877f
C4282 vdd.n2858 vss 0.00297f
C4283 vdd.n2859 vss 0.00594f
C4284 vdd.n2860 vss 0.00722f
C4285 vdd.n2861 vss 0.00524f
C4286 vdd.n2862 vss 0.00368f
C4287 vdd.n2863 vss 0.00297f
C4288 vdd.n2864 vss -0.0674f
C4289 vdd.n2865 vss 2.92e-19
C4290 vdd.n2866 vss 0.00437f
C4291 vdd.n2867 vss 0.00714f
C4292 vdd.n2868 vss 0.00836f
C4293 vdd.n2869 vss 0.0082f
C4294 vdd.n2870 vss 0.00502f
C4295 vdd.n2871 vss 0.00394f
C4296 vdd.n2872 vss 0.00423f
C4297 vdd.n2873 vss 0.00524f
C4298 vdd.n2874 vss 0.00594f
C4299 vdd.n2875 vss 0.00722f
C4300 vdd.n2876 vss 0.00311f
C4301 vdd.n2877 vss 0.00241f
C4302 vdd.n2878 vss 0.00311f
C4303 vdd.n2879 vss 2.83e-19
C4304 vdd.n2880 vss 0.00933f
C4305 vdd.n2881 vss 0.0115f
C4306 vdd.n2883 vss 0.00248f
C4307 vdd.n2884 vss 0.00241f
C4308 vdd.n2885 vss 2.83e-19
C4309 vdd.n2886 vss 0.00311f
C4310 vdd.n2887 vss 4.25e-19
C4311 vdd.n2888 vss 0.00437f
C4312 vdd.n2889 vss 0.00714f
C4313 vdd.n2890 vss -0.168f
C4314 vdd.n2891 vss 0.0082f
C4315 vdd.n2892 vss 0.00502f
C4316 vdd.n2893 vss 0.00394f
C4317 vdd.n2894 vss 0.00423f
C4318 vdd.n2895 vss 0.00524f
C4319 vdd.n2896 vss 0.00722f
C4320 vdd.n2897 vss 0.00594f
C4321 vdd.n2898 vss 0.00297f
C4322 vdd.n2899 vss 0.00877f
C4323 vdd.n2900 vss 0.00877f
C4324 vdd.n2901 vss 0.0115f
C4325 vdd.n2903 vss 0.00248f
C4326 vdd.n2904 vss 0.00933f
C4327 vdd.n2905 vss 2.83e-19
C4328 vdd.n2906 vss 0.00311f
C4329 vdd.n2907 vss 4.25e-19
C4330 vdd.n2908 vss 0.00437f
C4331 vdd.n2909 vss 0.00714f
C4332 vdd.n2910 vss 0.00836f
C4333 vdd.n2911 vss 0.0082f
C4334 vdd.n2912 vss 0.00502f
C4335 vdd.n2913 vss -0.0674f
C4336 vdd.n2914 vss -0.189f
C4337 vdd.n2915 vss 0.00524f
C4338 vdd.n2916 vss 0.00722f
C4339 vdd.n2917 vss 0.00594f
C4340 vdd.n2918 vss 0.00297f
C4341 vdd.n2919 vss 0.00877f
C4342 vdd.n2920 vss 0.00877f
C4343 vdd.n2921 vss 0.0115f
C4344 vdd.n2922 vss 0.00248f
C4345 vdd.n2923 vss 0.021f
C4346 vdd.n2924 vss 4.73e-19
C4347 vdd.n2925 vss 0.00311f
C4348 vdd.n2926 vss 4.25e-19
C4349 vdd.n2927 vss 0.00437f
C4350 vdd.n2928 vss 0.0257f
C4351 vdd.n2929 vss 0.0296f
C4352 vdd.n2930 vss 0.0294f
C4353 vdd.n2931 vss 0.00518f
C4354 vdd.n2932 vss 0.00502f
C4355 vdd.n2933 vss 2.92e-19
C4356 vdd.n2934 vss 0.00423f
C4357 vdd.n2935 vss 4.25e-19
C4358 vdd.n2936 vss 0.00311f
C4359 vdd.n2937 vss 4.73e-19
C4360 vdd.n2938 vss 0.021f
C4361 vdd.n2939 vss 0.00248f
C4362 vdd.n2940 vss 0.0115f
C4363 vdd.n2943 vss 0.00248f
C4364 vdd.n2944 vss 0.00933f
C4365 vdd.n2945 vss 2.83e-19
C4366 vdd.n2946 vss 0.00241f
C4367 vdd.n2947 vss 0.00877f
C4368 vdd.n2948 vss 0.00297f
C4369 vdd.n2949 vss 0.00594f
C4370 vdd.n2950 vss 0.00722f
C4371 vdd.n2951 vss 0.00524f
C4372 vdd.n2952 vss -0.189f
C4373 vdd.n2953 vss 0.0035f
C4374 vdd.n2954 vss 0.00423f
C4375 vdd.n2955 vss 0.007f
C4376 vdd.n2956 vss 0.0082f
C4377 vdd.n2957 vss 0.00502f
C4378 vdd.n2958 vss -0.175f
C4379 vdd.n2959 vss 0.00423f
C4380 vdd.n2960 vss 0.007f
C4381 vdd.n2961 vss 0.0035f
C4382 vdd.n2962 vss 0.00836f
C4383 vdd.n2963 vss 0.00518f
C4384 vdd.n2964 vss 0.00394f
C4385 vdd.n2965 vss 0.00297f
C4386 vdd.n2966 vss 0.00368f
C4387 vdd.n2967 vss 0.00821f
C4388 vdd.n2968 vss 0.00594f
C4389 vdd.n2969 vss 0.00722f
C4390 vdd.n2970 vss 0.00311f
C4391 vdd.n2971 vss 0.00241f
C4392 vdd.n2972 vss 0.00241f
C4393 vdd.n2973 vss 2.83e-19
C4394 vdd.n2974 vss 0.00933f
C4395 vdd.n2976 vss 0.00248f
C4396 vdd.n2978 vss 0.0115f
C4397 vdd.n2979 vss 0.00877f
C4398 vdd.n2980 vss 0.00877f
C4399 vdd.n2981 vss 0.00297f
C4400 vdd.n2982 vss 0.00311f
C4401 vdd.n2983 vss 0.00722f
C4402 vdd.n2984 vss 0.00594f
C4403 vdd.n2985 vss 0.00821f
C4404 vdd.n2986 vss 0.00368f
C4405 vdd.n2987 vss 0.00297f
C4406 vdd.n2988 vss 0.00394f
C4407 vdd.n2989 vss 0.00518f
C4408 vdd.n2990 vss 0.00836f
C4409 vdd.n2991 vss 0.0035f
C4410 vdd.n2992 vss 0.007f
C4411 vdd.n2993 vss 0.00423f
C4412 vdd.n2994 vss 2.92e-19
C4413 vdd.n2995 vss 0.00502f
C4414 vdd.n2996 vss 0.00518f
C4415 vdd.n2997 vss 0.00836f
C4416 vdd.n2998 vss 0.0035f
C4417 vdd.n2999 vss -0.189f
C4418 vdd.n3000 vss 0.00524f
C4419 vdd.n3001 vss 0.00368f
C4420 vdd.n3002 vss 0.00821f
C4421 vdd.n3003 vss 0.00311f
C4422 vdd.n3004 vss 2.83e-19
C4423 vdd.n3005 vss 0.00241f
C4424 vdd.n3006 vss 0.00248f
C4425 vdd.n3008 vss 0.0115f
C4426 vdd.n3010 vss 0.00933f
C4427 vdd.n3011 vss 2.83e-19
C4428 vdd.n3012 vss 0.00311f
C4429 vdd.n3013 vss 4.25e-19
C4430 vdd.n3014 vss 0.00423f
C4431 vdd.n3015 vss 2.92e-19
C4432 vdd.n3016 vss 0.00502f
C4433 vdd.n3017 vss 0.00518f
C4434 vdd.n3018 vss 0.00836f
C4435 vdd.n3019 vss 0.0035f
C4436 vdd.n3020 vss 0.00437f
C4437 vdd.n3021 vss 0.00524f
C4438 vdd.n3022 vss 0.00722f
C4439 vdd.n3023 vss 0.00594f
C4440 vdd.n3024 vss 0.00297f
C4441 vdd.n3025 vss 0.00877f
C4442 vdd.n3026 vss 0.00877f
C4443 vdd.n3027 vss 0.0115f
C4444 vdd.n3029 vss 0.0155f
C4445 vdd.n3030 vss 0.028f
C4446 vdd.n3031 vss 0.028f
C4447 vdd.n3032 vss 0.0155f
C4448 vdd.n3033 vss 0.00248f
C4449 vdd.n3034 vss 0.00933f
C4450 vdd.n3035 vss 2.83e-19
C4451 vdd.n3036 vss 0.00311f
C4452 vdd.n3037 vss 4.25e-19
C4453 vdd.n3038 vss 0.00423f
C4454 vdd.n3039 vss 2.92e-19
C4455 vdd.n3040 vss -0.0772f
C4456 vdd.n3041 vss 0.00518f
C4457 vdd.n3042 vss 0.0221f
C4458 vdd.n3043 vss 0.0217f
C4459 vdd.n3044 vss 0.00437f
C4460 vdd.n3045 vss 0.0225f
C4461 vdd.n3046 vss 0.00368f
C4462 vdd.n3047 vss 0.0225f
C4463 vdd.n3048 vss 0.00423f
C4464 vdd.n3049 vss 0.00394f
C4465 vdd.n3050 vss 0.00502f
C4466 vdd.n3051 vss -0.0832f
C4467 vdd.n3052 vss -0.168f
C4468 vdd.n3053 vss 0.00714f
C4469 vdd.n3054 vss 0.00437f
C4470 vdd.n3055 vss 4.25e-19
C4471 vdd.n3056 vss 0.00311f
C4472 vdd.n3057 vss 2.83e-19
C4473 vdd.n3058 vss 0.00933f
C4474 vdd.n3060 vss 0.0115f
C4475 vdd.n3061 vss 0.00877f
C4476 vdd.n3062 vss 0.00877f
C4477 vdd.n3063 vss 0.00297f
C4478 vdd.n3064 vss 0.00594f
C4479 vdd.n3065 vss 0.00722f
C4480 vdd.n3066 vss 0.00368f
C4481 vdd.n3067 vss 0.00524f
C4482 vdd.n3068 vss 0.00423f
C4483 vdd.n3069 vss 0.00394f
C4484 vdd.n3070 vss 0.00502f
C4485 vdd.n3071 vss 0.00518f
C4486 vdd.n3072 vss 0.0082f
C4487 vdd.n3073 vss 0.00836f
C4488 vdd.n3074 vss 0.00714f
C4489 vdd.n3075 vss 0.00437f
C4490 vdd.n3076 vss 4.25e-19
C4491 vdd.n3077 vss 0.00311f
C4492 vdd.n3078 vss 2.83e-19
C4493 vdd.n3079 vss 0.00933f
C4494 vdd.n3081 vss 0.0115f
C4495 vdd.n3082 vss 0.00877f
C4496 vdd.n3083 vss 0.00877f
C4497 vdd.n3084 vss 0.00297f
C4498 vdd.n3085 vss 0.00594f
C4499 vdd.n3086 vss 0.00722f
C4500 vdd.n3087 vss 0.00524f
C4501 vdd.n3088 vss 0.00368f
C4502 vdd.n3089 vss 0.00297f
C4503 vdd.n3090 vss -0.0674f
C4504 vdd.n3091 vss 2.92e-19
C4505 vdd.n3092 vss 0.00437f
C4506 vdd.n3093 vss 0.00714f
C4507 vdd.n3094 vss 0.00836f
C4508 vdd.n3095 vss 0.0082f
C4509 vdd.n3096 vss 0.00502f
C4510 vdd.n3097 vss 0.00394f
C4511 vdd.n3098 vss 0.00423f
C4512 vdd.n3099 vss 0.00524f
C4513 vdd.n3100 vss 0.00594f
C4514 vdd.n3101 vss 0.00722f
C4515 vdd.n3102 vss 0.00311f
C4516 vdd.n3103 vss 0.00241f
C4517 vdd.n3104 vss 0.00311f
C4518 vdd.n3105 vss 2.83e-19
C4519 vdd.n3106 vss 0.00933f
C4520 vdd.n3107 vss 0.0115f
C4521 vdd.n3109 vss 0.00248f
C4522 vdd.n3110 vss 0.00241f
C4523 vdd.n3111 vss 2.83e-19
C4524 vdd.n3112 vss 0.00311f
C4525 vdd.n3113 vss 4.25e-19
C4526 vdd.n3114 vss 0.00437f
C4527 vdd.n3115 vss 0.00714f
C4528 vdd.n3116 vss -0.168f
C4529 vdd.n3117 vss 0.0082f
C4530 vdd.n3118 vss 0.00502f
C4531 vdd.n3119 vss 0.00394f
C4532 vdd.n3120 vss 0.00423f
C4533 vdd.n3121 vss 0.00524f
C4534 vdd.n3122 vss 0.00722f
C4535 vdd.n3123 vss 0.00594f
C4536 vdd.n3124 vss 0.00297f
C4537 vdd.n3125 vss 0.00877f
C4538 vdd.n3126 vss 0.00877f
C4539 vdd.n3127 vss 0.0115f
C4540 vdd.n3129 vss 0.00248f
C4541 vdd.n3130 vss 0.00933f
C4542 vdd.n3131 vss 2.83e-19
C4543 vdd.n3132 vss 0.00311f
C4544 vdd.n3133 vss 4.25e-19
C4545 vdd.n3134 vss 0.00437f
C4546 vdd.n3135 vss 0.00714f
C4547 vdd.n3136 vss 0.00836f
C4548 vdd.n3137 vss 0.0082f
C4549 vdd.n3138 vss 0.00502f
C4550 vdd.n3139 vss -0.0674f
C4551 vdd.n3140 vss -0.189f
C4552 vdd.n3141 vss 0.00524f
C4553 vdd.n3142 vss 0.00722f
C4554 vdd.n3143 vss 0.00594f
C4555 vdd.n3144 vss 0.00297f
C4556 vdd.n3145 vss 0.00877f
C4557 vdd.n3146 vss 0.00877f
C4558 vdd.n3147 vss 0.0115f
C4559 vdd.n3148 vss 0.00248f
C4560 vdd.n3149 vss 0.021f
C4561 vdd.n3150 vss 4.73e-19
C4562 vdd.n3151 vss 0.00311f
C4563 vdd.n3152 vss 4.25e-19
C4564 vdd.n3153 vss 0.00437f
C4565 vdd.n3154 vss 0.0257f
C4566 vdd.n3155 vss 0.0296f
C4567 vdd.n3156 vss 0.0294f
C4568 vdd.n3157 vss 0.00518f
C4569 vdd.n3158 vss 0.00502f
C4570 vdd.n3159 vss 2.92e-19
C4571 vdd.n3160 vss 0.00423f
C4572 vdd.n3161 vss 4.25e-19
C4573 vdd.n3162 vss 0.00311f
C4574 vdd.n3163 vss 4.73e-19
C4575 vdd.n3164 vss 0.021f
C4576 vdd.n3165 vss 0.00248f
C4577 vdd.n3166 vss 0.0115f
C4578 vdd.n3169 vss 0.00248f
C4579 vdd.n3170 vss 0.00933f
C4580 vdd.n3171 vss 2.83e-19
C4581 vdd.n3172 vss 0.00241f
C4582 vdd.n3173 vss 0.00877f
C4583 vdd.n3174 vss 0.00297f
C4584 vdd.n3175 vss 0.00594f
C4585 vdd.n3176 vss 0.00722f
C4586 vdd.n3177 vss 0.00524f
C4587 vdd.n3178 vss -0.189f
C4588 vdd.n3179 vss 0.0035f
C4589 vdd.n3180 vss 0.00423f
C4590 vdd.n3181 vss 0.007f
C4591 vdd.n3182 vss 0.0082f
C4592 vdd.n3183 vss 0.00502f
C4593 vdd.n3184 vss -0.175f
C4594 vdd.n3185 vss 0.00423f
C4595 vdd.n3186 vss 0.007f
C4596 vdd.n3187 vss 0.0035f
C4597 vdd.n3188 vss 0.00836f
C4598 vdd.n3189 vss 0.00518f
C4599 vdd.n3190 vss 0.00394f
C4600 vdd.n3191 vss 0.00297f
C4601 vdd.n3192 vss 0.00368f
C4602 vdd.n3193 vss 0.00821f
C4603 vdd.n3194 vss 0.00594f
C4604 vdd.n3195 vss 0.00722f
C4605 vdd.n3196 vss 0.00311f
C4606 vdd.n3197 vss 0.00241f
C4607 vdd.n3198 vss 0.00241f
C4608 vdd.n3199 vss 2.83e-19
C4609 vdd.n3200 vss 0.00933f
C4610 vdd.n3202 vss 0.00248f
C4611 vdd.n3204 vss 0.0115f
C4612 vdd.n3205 vss 0.00877f
C4613 vdd.n3206 vss 0.00877f
C4614 vdd.n3207 vss 0.00297f
C4615 vdd.n3208 vss 0.00311f
C4616 vdd.n3209 vss 0.00722f
C4617 vdd.n3210 vss 0.00594f
C4618 vdd.n3211 vss 0.00821f
C4619 vdd.n3212 vss 0.00368f
C4620 vdd.n3213 vss 0.00297f
C4621 vdd.n3214 vss 0.00394f
C4622 vdd.n3215 vss 0.00518f
C4623 vdd.n3216 vss 0.00836f
C4624 vdd.n3217 vss 0.0035f
C4625 vdd.n3218 vss 0.007f
C4626 vdd.n3219 vss 0.00423f
C4627 vdd.n3220 vss 2.92e-19
C4628 vdd.n3221 vss 0.00502f
C4629 vdd.n3222 vss 0.00518f
C4630 vdd.n3223 vss 0.00836f
C4631 vdd.n3224 vss 0.0035f
C4632 vdd.n3225 vss -0.189f
C4633 vdd.n3226 vss 0.00524f
C4634 vdd.n3227 vss 0.00368f
C4635 vdd.n3228 vss 0.00821f
C4636 vdd.n3229 vss 0.00311f
C4637 vdd.n3230 vss 2.83e-19
C4638 vdd.n3231 vss 0.00241f
C4639 vdd.n3232 vss 0.00248f
C4640 vdd.n3234 vss 0.0115f
C4641 vdd.n3236 vss 0.00933f
C4642 vdd.n3237 vss 2.83e-19
C4643 vdd.n3238 vss 0.00311f
C4644 vdd.n3239 vss 4.25e-19
C4645 vdd.n3240 vss 0.00423f
C4646 vdd.n3241 vss 2.92e-19
C4647 vdd.n3242 vss 0.00502f
C4648 vdd.n3243 vss 0.00518f
C4649 vdd.n3244 vss 0.00836f
C4650 vdd.n3245 vss 0.0035f
C4651 vdd.n3246 vss 0.00437f
C4652 vdd.n3247 vss 0.00524f
C4653 vdd.n3248 vss 0.00722f
C4654 vdd.n3249 vss 0.00594f
C4655 vdd.n3250 vss 0.00297f
C4656 vdd.n3251 vss 0.00877f
C4657 vdd.n3252 vss 0.00877f
C4658 vdd.n3253 vss 0.0115f
C4659 vdd.n3255 vss 0.0155f
C4660 vdd.n3256 vss 0.028f
C4661 vdd.n3257 vss 0.028f
C4662 vdd.n3258 vss 0.0155f
C4663 vdd.n3259 vss 0.00248f
C4664 vdd.n3260 vss 0.00933f
C4665 vdd.n3261 vss 2.83e-19
C4666 vdd.n3262 vss 0.00311f
C4667 vdd.n3263 vss 4.25e-19
C4668 vdd.n3264 vss 0.00423f
C4669 vdd.n3265 vss 2.92e-19
C4670 vdd.n3266 vss -0.0772f
C4671 vdd.n3267 vss 0.00518f
C4672 vdd.n3268 vss 0.0221f
C4673 vdd.n3269 vss 0.0217f
C4674 vdd.n3270 vss 0.00437f
C4675 vdd.n3271 vss 0.0225f
C4676 vdd.n3272 vss 0.00368f
C4677 vdd.n3273 vss 0.0225f
C4678 vdd.n3274 vss 0.00423f
C4679 vdd.n3275 vss 0.00394f
C4680 vdd.n3276 vss 0.00502f
C4681 vdd.n3277 vss -0.0832f
C4682 vdd.n3278 vss -0.168f
C4683 vdd.n3279 vss 0.00714f
C4684 vdd.n3280 vss 0.00437f
C4685 vdd.n3281 vss 4.25e-19
C4686 vdd.n3282 vss 0.00311f
C4687 vdd.n3283 vss 2.83e-19
C4688 vdd.n3284 vss 0.00933f
C4689 vdd.n3286 vss 0.0115f
C4690 vdd.n3287 vss 0.00877f
C4691 vdd.n3288 vss 0.00877f
C4692 vdd.n3289 vss 0.00297f
C4693 vdd.n3290 vss 0.00594f
C4694 vdd.n3291 vss 0.00722f
C4695 vdd.n3292 vss 0.00368f
C4696 vdd.n3293 vss 0.00524f
C4697 vdd.n3294 vss 0.00423f
C4698 vdd.n3295 vss 0.00394f
C4699 vdd.n3296 vss 0.00502f
C4700 vdd.n3297 vss 0.00518f
C4701 vdd.n3298 vss 0.0082f
C4702 vdd.n3299 vss 0.00836f
C4703 vdd.n3300 vss 0.00714f
C4704 vdd.n3301 vss 0.00437f
C4705 vdd.n3302 vss 4.25e-19
C4706 vdd.n3303 vss 0.00311f
C4707 vdd.n3304 vss 2.83e-19
C4708 vdd.n3305 vss 0.00933f
C4709 vdd.n3307 vss 0.0115f
C4710 vdd.n3308 vss 0.00877f
C4711 vdd.n3309 vss 0.00877f
C4712 vdd.n3310 vss 0.00297f
C4713 vdd.n3311 vss 0.00594f
C4714 vdd.n3312 vss 0.00722f
C4715 vdd.n3313 vss 0.00524f
C4716 vdd.n3314 vss 0.00368f
C4717 vdd.n3315 vss 0.00297f
C4718 vdd.n3316 vss -0.0674f
C4719 vdd.n3317 vss 2.92e-19
C4720 vdd.n3318 vss 0.00437f
C4721 vdd.n3319 vss 0.00714f
C4722 vdd.n3320 vss 0.00836f
C4723 vdd.n3321 vss 0.0082f
C4724 vdd.n3322 vss 0.00502f
C4725 vdd.n3323 vss 0.00394f
C4726 vdd.n3324 vss 0.00423f
C4727 vdd.n3325 vss 0.00524f
C4728 vdd.n3326 vss 0.00594f
C4729 vdd.n3327 vss 0.00722f
C4730 vdd.n3328 vss 0.00311f
C4731 vdd.n3329 vss 0.00241f
C4732 vdd.n3330 vss 0.00311f
C4733 vdd.n3331 vss 2.83e-19
C4734 vdd.n3332 vss 0.00933f
C4735 vdd.n3333 vss 0.0115f
C4736 vdd.n3335 vss 0.00248f
C4737 vdd.n3336 vss 0.00241f
C4738 vdd.n3337 vss 2.83e-19
C4739 vdd.n3338 vss 0.00311f
C4740 vdd.n3339 vss 4.25e-19
C4741 vdd.n3340 vss 0.00437f
C4742 vdd.n3341 vss 0.00714f
C4743 vdd.n3342 vss -0.168f
C4744 vdd.n3343 vss 0.0082f
C4745 vdd.n3344 vss 0.00502f
C4746 vdd.n3345 vss 0.00394f
C4747 vdd.n3346 vss 0.00423f
C4748 vdd.n3347 vss 0.00524f
C4749 vdd.n3348 vss 0.00722f
C4750 vdd.n3349 vss 0.00594f
C4751 vdd.n3350 vss 0.00297f
C4752 vdd.n3351 vss 0.00877f
C4753 vdd.n3352 vss 0.00877f
C4754 vdd.n3353 vss 0.0115f
C4755 vdd.n3355 vss 0.00248f
C4756 vdd.n3356 vss 0.00933f
C4757 vdd.n3357 vss 2.83e-19
C4758 vdd.n3358 vss 0.00311f
C4759 vdd.n3359 vss 4.25e-19
C4760 vdd.n3360 vss 0.00437f
C4761 vdd.n3361 vss 0.00714f
C4762 vdd.n3362 vss 0.00836f
C4763 vdd.n3363 vss 0.0082f
C4764 vdd.n3364 vss 0.00502f
C4765 vdd.n3365 vss -0.0674f
C4766 vdd.n3366 vss -0.189f
C4767 vdd.n3367 vss 0.00524f
C4768 vdd.n3368 vss 0.00722f
C4769 vdd.n3369 vss 0.00594f
C4770 vdd.n3370 vss 0.00297f
C4771 vdd.n3371 vss 0.00877f
C4772 vdd.n3372 vss 0.00877f
C4773 vdd.n3373 vss 0.0115f
C4774 vdd.n3374 vss 0.00248f
C4775 vdd.n3375 vss 0.021f
C4776 vdd.n3376 vss 4.73e-19
C4777 vdd.n3377 vss 0.00311f
C4778 vdd.n3378 vss 4.25e-19
C4779 vdd.n3379 vss 0.00437f
C4780 vdd.n3380 vss 0.0257f
C4781 vdd.n3381 vss 0.0296f
C4782 vdd.n3382 vss 0.0294f
C4783 vdd.n3383 vss 0.00518f
C4784 vdd.n3384 vss 0.00502f
C4785 vdd.n3385 vss 2.92e-19
C4786 vdd.n3386 vss 0.00423f
C4787 vdd.n3387 vss 4.25e-19
C4788 vdd.n3388 vss 0.00311f
C4789 vdd.n3389 vss 4.73e-19
C4790 vdd.n3390 vss 0.021f
C4791 vdd.n3391 vss 0.00248f
C4792 vdd.n3392 vss 0.0115f
C4793 vdd.n3395 vss 0.00248f
C4794 vdd.n3396 vss 0.00933f
C4795 vdd.n3397 vss 2.83e-19
C4796 vdd.n3398 vss 0.00241f
C4797 vdd.n3399 vss 0.00877f
C4798 vdd.n3400 vss 0.00297f
C4799 vdd.n3401 vss 0.00594f
C4800 vdd.n3402 vss 0.00722f
C4801 vdd.n3403 vss 0.00524f
C4802 vdd.n3404 vss -0.189f
C4803 vdd.n3405 vss 0.0035f
C4804 vdd.n3406 vss 0.00423f
C4805 vdd.n3407 vss 0.007f
C4806 vdd.n3408 vss 0.0082f
C4807 vdd.n3409 vss 0.00502f
C4808 vdd.n3410 vss -0.175f
C4809 vdd.n3411 vss 0.00423f
C4810 vdd.n3412 vss 0.007f
C4811 vdd.n3413 vss 0.0035f
C4812 vdd.n3414 vss 0.00836f
C4813 vdd.n3415 vss 0.00518f
C4814 vdd.n3416 vss 0.00394f
C4815 vdd.n3417 vss 0.00297f
C4816 vdd.n3418 vss 0.00368f
C4817 vdd.n3419 vss 0.00821f
C4818 vdd.n3420 vss 0.00594f
C4819 vdd.n3421 vss 0.00722f
C4820 vdd.n3422 vss 0.00311f
C4821 vdd.n3423 vss 0.00241f
C4822 vdd.n3424 vss 0.00241f
C4823 vdd.n3425 vss 2.83e-19
C4824 vdd.n3426 vss 0.00933f
C4825 vdd.n3428 vss 0.00248f
C4826 vdd.n3430 vss 0.0115f
C4827 vdd.n3431 vss 0.00877f
C4828 vdd.n3432 vss 0.00877f
C4829 vdd.n3433 vss 0.00297f
C4830 vdd.n3434 vss 0.00311f
C4831 vdd.n3435 vss 0.00722f
C4832 vdd.n3436 vss 0.00594f
C4833 vdd.n3437 vss 0.00821f
C4834 vdd.n3438 vss 0.00368f
C4835 vdd.n3439 vss 0.00297f
C4836 vdd.n3440 vss 0.00394f
C4837 vdd.n3441 vss 0.00518f
C4838 vdd.n3442 vss 0.00836f
C4839 vdd.n3443 vss 0.0035f
C4840 vdd.n3444 vss 0.007f
C4841 vdd.n3445 vss 0.00423f
C4842 vdd.n3446 vss 2.92e-19
C4843 vdd.n3447 vss 0.00502f
C4844 vdd.n3448 vss 0.00518f
C4845 vdd.n3449 vss 0.00836f
C4846 vdd.n3450 vss 0.0035f
C4847 vdd.n3451 vss -0.189f
C4848 vdd.n3452 vss 0.00524f
C4849 vdd.n3453 vss 0.00368f
C4850 vdd.n3454 vss 0.00821f
C4851 vdd.n3455 vss 0.00311f
C4852 vdd.n3456 vss 2.83e-19
C4853 vdd.n3457 vss 0.00241f
C4854 vdd.n3458 vss 0.00248f
C4855 vdd.n3460 vss 0.0115f
C4856 vdd.n3462 vss 0.00933f
C4857 vdd.n3463 vss 2.83e-19
C4858 vdd.n3464 vss 0.00311f
C4859 vdd.n3465 vss 4.25e-19
C4860 vdd.n3466 vss 0.00423f
C4861 vdd.n3467 vss 2.92e-19
C4862 vdd.n3468 vss 0.00502f
C4863 vdd.n3469 vss 0.00518f
C4864 vdd.n3470 vss 0.00836f
C4865 vdd.n3471 vss 0.0035f
C4866 vdd.n3472 vss 0.00437f
C4867 vdd.n3473 vss 0.00524f
C4868 vdd.n3474 vss 0.00722f
C4869 vdd.n3475 vss 0.00594f
C4870 vdd.n3476 vss 0.00297f
C4871 vdd.n3477 vss 0.00877f
C4872 vdd.n3478 vss 0.00877f
C4873 vdd.n3479 vss 0.0115f
C4874 vdd.n3481 vss 0.0155f
C4875 vdd.n3482 vss 0.028f
C4876 vdd.n3483 vss 0.028f
C4877 vdd.n3484 vss 0.0155f
C4878 vdd.n3485 vss 0.00248f
C4879 vdd.n3486 vss 0.00933f
C4880 vdd.n3487 vss 2.83e-19
C4881 vdd.n3488 vss 0.00311f
C4882 vdd.n3489 vss 4.25e-19
C4883 vdd.n3490 vss 0.00423f
C4884 vdd.n3491 vss 2.92e-19
C4885 vdd.n3492 vss -0.0772f
C4886 vdd.n3493 vss 0.00518f
C4887 vdd.n3494 vss 0.0221f
C4888 vdd.n3495 vss 0.0217f
C4889 vdd.n3496 vss 0.00437f
C4890 vdd.n3497 vss 0.0225f
C4891 vdd.n3498 vss 0.00368f
C4892 vdd.n3499 vss 0.0225f
C4893 vdd.n3500 vss 0.00423f
C4894 vdd.n3501 vss 0.00394f
C4895 vdd.n3502 vss 0.00502f
C4896 vdd.n3503 vss -0.0832f
C4897 vdd.n3504 vss -0.168f
C4898 vdd.n3505 vss 0.00714f
C4899 vdd.n3506 vss 0.00437f
C4900 vdd.n3507 vss 4.25e-19
C4901 vdd.n3508 vss 0.00311f
C4902 vdd.n3509 vss 2.83e-19
C4903 vdd.n3510 vss 0.00933f
C4904 vdd.n3512 vss 0.0115f
C4905 vdd.n3513 vss 0.00877f
C4906 vdd.n3514 vss 0.00877f
C4907 vdd.n3515 vss 0.00297f
C4908 vdd.n3516 vss 0.00594f
C4909 vdd.n3517 vss 0.00722f
C4910 vdd.n3518 vss 0.00368f
C4911 vdd.n3519 vss 0.00524f
C4912 vdd.n3520 vss 0.00423f
C4913 vdd.n3521 vss 0.00394f
C4914 vdd.n3522 vss 0.00502f
C4915 vdd.n3523 vss 0.00518f
C4916 vdd.n3524 vss 0.0082f
C4917 vdd.n3525 vss 0.00836f
C4918 vdd.n3526 vss 0.00714f
C4919 vdd.n3527 vss 0.00437f
C4920 vdd.n3528 vss 4.25e-19
C4921 vdd.n3529 vss 0.00311f
C4922 vdd.n3530 vss 2.83e-19
C4923 vdd.n3531 vss 0.00933f
C4924 vdd.n3533 vss 0.0115f
C4925 vdd.n3534 vss 0.00877f
C4926 vdd.n3535 vss 0.00877f
C4927 vdd.n3536 vss 0.00297f
C4928 vdd.n3537 vss 0.00594f
C4929 vdd.n3538 vss 0.00722f
C4930 vdd.n3539 vss 0.00524f
C4931 vdd.n3540 vss 0.00368f
C4932 vdd.n3541 vss 0.00297f
C4933 vdd.n3542 vss -0.0674f
C4934 vdd.n3543 vss 2.92e-19
C4935 vdd.n3544 vss 0.00437f
C4936 vdd.n3545 vss 0.00714f
C4937 vdd.n3546 vss 0.00836f
C4938 vdd.n3547 vss 0.0082f
C4939 vdd.n3548 vss 0.00502f
C4940 vdd.n3549 vss 0.00394f
C4941 vdd.n3550 vss 0.00423f
C4942 vdd.n3551 vss 0.00524f
C4943 vdd.n3552 vss 0.00594f
C4944 vdd.n3553 vss 0.00722f
C4945 vdd.n3554 vss 0.00311f
C4946 vdd.n3555 vss 0.00241f
C4947 vdd.n3556 vss 0.00311f
C4948 vdd.n3557 vss 2.83e-19
C4949 vdd.n3558 vss 0.00933f
C4950 vdd.n3559 vss 0.0115f
C4951 vdd.n3561 vss 0.00248f
C4952 vdd.n3562 vss 0.00241f
C4953 vdd.n3563 vss 2.83e-19
C4954 vdd.n3564 vss 0.00311f
C4955 vdd.n3565 vss 4.25e-19
C4956 vdd.n3566 vss 0.00437f
C4957 vdd.n3567 vss 0.00714f
C4958 vdd.n3568 vss -0.168f
C4959 vdd.n3569 vss 0.0082f
C4960 vdd.n3570 vss 0.00502f
C4961 vdd.n3571 vss 0.00394f
C4962 vdd.n3572 vss 0.00423f
C4963 vdd.n3573 vss 0.00524f
C4964 vdd.n3574 vss 0.00722f
C4965 vdd.n3575 vss 0.00594f
C4966 vdd.n3576 vss 0.00297f
C4967 vdd.n3577 vss 0.00877f
C4968 vdd.n3578 vss 0.00877f
C4969 vdd.n3579 vss 0.0115f
C4970 vdd.n3581 vss 0.00248f
C4971 vdd.n3582 vss 0.00933f
C4972 vdd.n3583 vss 2.83e-19
C4973 vdd.n3584 vss 0.00311f
C4974 vdd.n3585 vss 4.25e-19
C4975 vdd.n3586 vss 0.00437f
C4976 vdd.n3587 vss 0.00714f
C4977 vdd.n3588 vss 0.00836f
C4978 vdd.n3589 vss 0.0082f
C4979 vdd.n3590 vss 0.00502f
C4980 vdd.n3591 vss -0.0674f
C4981 vdd.n3592 vss -0.189f
C4982 vdd.n3593 vss 0.00524f
C4983 vdd.n3594 vss 0.00722f
C4984 vdd.n3595 vss 0.00594f
C4985 vdd.n3596 vss 0.00297f
C4986 vdd.n3597 vss 0.00877f
C4987 vdd.n3598 vss 0.00877f
C4988 vdd.n3599 vss 0.0115f
C4989 vdd.n3600 vss 0.00248f
C4990 vdd.n3601 vss 0.021f
C4991 vdd.n3602 vss 4.73e-19
C4992 vdd.n3603 vss 0.00311f
C4993 vdd.n3604 vss 4.25e-19
C4994 vdd.n3605 vss 0.00437f
C4995 vdd.n3606 vss 0.0257f
C4996 vdd.n3607 vss 0.0296f
C4997 vdd.n3608 vss 0.0294f
C4998 vdd.n3609 vss 0.00518f
C4999 vdd.n3610 vss 0.00502f
C5000 vdd.n3611 vss 2.92e-19
C5001 vdd.n3612 vss 0.00423f
C5002 vdd.n3613 vss 4.25e-19
C5003 vdd.n3614 vss 0.00311f
C5004 vdd.n3615 vss 4.73e-19
C5005 vdd.n3616 vss 0.021f
C5006 vdd.n3617 vss 0.00248f
C5007 vdd.n3618 vss 0.0115f
C5008 vdd.n3621 vss 0.00248f
C5009 vdd.n3622 vss 0.00933f
C5010 vdd.n3623 vss 2.83e-19
C5011 vdd.n3624 vss 0.00241f
C5012 vdd.n3625 vss 0.00877f
C5013 vdd.n3626 vss 0.00297f
C5014 vdd.n3627 vss 0.00594f
C5015 vdd.n3628 vss 0.00722f
C5016 vdd.n3629 vss 0.00524f
C5017 vdd.n3630 vss -0.189f
C5018 vdd.n3631 vss 0.0035f
C5019 vdd.n3632 vss 0.00423f
C5020 vdd.n3633 vss 0.007f
C5021 vdd.n3634 vss 0.0082f
C5022 vdd.n3635 vss 0.00502f
C5023 vdd.n3636 vss -0.175f
C5024 vdd.n3637 vss 0.00423f
C5025 vdd.n3638 vss 0.007f
C5026 vdd.n3639 vss 0.0035f
C5027 vdd.n3640 vss 0.00836f
C5028 vdd.n3641 vss 0.00518f
C5029 vdd.n3642 vss 0.00394f
C5030 vdd.n3643 vss 0.00297f
C5031 vdd.n3644 vss 0.00368f
C5032 vdd.n3645 vss 0.00821f
C5033 vdd.n3646 vss 0.00594f
C5034 vdd.n3647 vss 0.00722f
C5035 vdd.n3648 vss 0.00311f
C5036 vdd.n3649 vss 0.00241f
C5037 vdd.n3650 vss 0.00241f
C5038 vdd.n3651 vss 2.83e-19
C5039 vdd.n3652 vss 0.00933f
C5040 vdd.n3654 vss 0.00248f
C5041 vdd.n3656 vss 0.0115f
C5042 vdd.n3657 vss 0.00877f
C5043 vdd.n3658 vss 0.00877f
C5044 vdd.n3659 vss 0.00297f
C5045 vdd.n3660 vss 0.00311f
C5046 vdd.n3661 vss 0.00722f
C5047 vdd.n3662 vss 0.00594f
C5048 vdd.n3663 vss 0.00821f
C5049 vdd.n3664 vss 0.00368f
C5050 vdd.n3665 vss 0.00297f
C5051 vdd.n3666 vss 0.00394f
C5052 vdd.n3667 vss 0.00518f
C5053 vdd.n3668 vss 0.00836f
C5054 vdd.n3669 vss 0.0035f
C5055 vdd.n3670 vss 0.007f
C5056 vdd.n3671 vss 0.00423f
C5057 vdd.n3672 vss 2.92e-19
C5058 vdd.n3673 vss 0.00502f
C5059 vdd.n3674 vss 0.00518f
C5060 vdd.n3675 vss 0.00836f
C5061 vdd.n3676 vss 0.0035f
C5062 vdd.n3677 vss -0.189f
C5063 vdd.n3678 vss 0.00524f
C5064 vdd.n3679 vss 0.00368f
C5065 vdd.n3680 vss 0.00821f
C5066 vdd.n3681 vss 0.00311f
C5067 vdd.n3682 vss 2.83e-19
C5068 vdd.n3683 vss 0.00241f
C5069 vdd.n3684 vss 0.00248f
C5070 vdd.n3686 vss 0.0115f
C5071 vdd.n3688 vss 0.00933f
C5072 vdd.n3689 vss 2.83e-19
C5073 vdd.n3690 vss 0.00311f
C5074 vdd.n3691 vss 4.25e-19
C5075 vdd.n3692 vss 0.00423f
C5076 vdd.n3693 vss 2.92e-19
C5077 vdd.n3694 vss 0.00502f
C5078 vdd.n3695 vss 0.00518f
C5079 vdd.n3696 vss 0.00423f
C5080 vdd.n3697 vss 2.92e-19
C5081 vdd.n3698 vss -0.0772f
C5082 vdd.n3699 vss -0.175f
C5083 vdd.n3700 vss 0.00836f
C5084 vdd.n3701 vss 0.0035f
C5085 vdd.n3702 vss 0.00437f
C5086 vdd.n3703 vss 0.00524f
C5087 vdd.n3704 vss 0.00311f
C5088 vdd.n3705 vss 0.00722f
C5089 vdd.n3706 vss 0.00594f
C5090 vdd.n3707 vss 0.00297f
C5091 vdd.n3708 vss 0.00877f
C5092 vdd.n3709 vss 0.00877f
C5093 vdd.n3710 vss 0.0115f
C5094 vdd.n3711 vss 0.0181f
C5095 vdd.n3712 vss 0.0462f
C5096 vdd.n3713 vss 0.0378f
C5097 vdd.n3714 vss 0.0349f
C5098 vdd.n3715 vss 0.0357f
C5099 vdd.n3716 vss 0.0221f
C5100 vdd.n3717 vss 0.0349f
C5101 vdd.n3718 vss 0.00297f
C5102 vdd.n3719 vss 0.00248f
C5103 vdd.n3720 vss 0.0211f
C5104 vdd.n3721 vss 0.0282f
C5105 vdd.n3722 vss 0.0516f
C5106 vdd.n3723 vss 0.0388f
C5107 vdd.n3724 vss 0.0393f
C5108 vdd.n3725 vss 2.92e-19
C5109 vdd.n3726 vss 0.00521f
C5110 vdd.n3727 vss 0.00538f
C5111 vdd.n3728 vss 0.00868f
C5112 vdd.n3729 vss 0.0035f
C5113 vdd.n3730 vss -0.189f
C5114 vdd.n3731 vss 0.00524f
C5115 vdd.n3732 vss 0.00722f
C5116 vdd.n3733 vss 0.00594f
C5117 vdd.n3734 vss 0.00297f
C5118 vdd.n3735 vss 0.00877f
C5119 vdd.n3736 vss 0.00877f
C5120 vdd.n3737 vss 0.0115f
C5121 vdd.n3739 vss 0.00933f
C5122 vdd.n3740 vss 2.83e-19
C5123 vdd.n3741 vss 0.00311f
C5124 vdd.n3742 vss 4.25e-19
C5125 vdd.n3743 vss 0.00423f
C5126 vdd.n3744 vss 2.92e-19
C5127 vdd.n3745 vss 0.00521f
C5128 vdd.n3746 vss 0.00538f
C5129 vdd.n3747 vss 0.00868f
C5130 vdd.n3748 vss 0.0035f
C5131 vdd.n3749 vss 0.00437f
C5132 vdd.n3750 vss 0.00524f
C5133 vdd.n3751 vss 0.00722f
C5134 vdd.n3752 vss 0.00594f
C5135 vdd.n3753 vss 0.00297f
C5136 vdd.n3754 vss 0.00877f
C5137 vdd.n3755 vss 0.00877f
C5138 vdd.n3756 vss 0.0115f
C5139 vdd.n3758 vss 0.00933f
C5140 vdd.n3759 vss 2.83e-19
C5141 vdd.n3760 vss 0.00311f
C5142 vdd.n3761 vss 4.25e-19
C5143 vdd.n3762 vss 0.00423f
C5144 vdd.n3763 vss 2.92e-19
C5145 vdd.n3764 vss -0.077f
C5146 vdd.n3765 vss 0.00538f
C5147 vdd.n3766 vss 0.00868f
C5148 vdd.n3767 vss 0.0035f
C5149 vdd.n3768 vss 0.00437f
C5150 vdd.n3769 vss 0.00524f
C5151 vdd.n3770 vss 0.00722f
C5152 vdd.n3771 vss 0.00594f
C5153 vdd.n3772 vss 0.00297f
C5154 vdd.n3773 vss 0.00877f
C5155 vdd.n3774 vss 0.00877f
C5156 vdd.n3775 vss 0.0115f
C5157 vdd.n3777 vss 0.00933f
C5158 vdd.n3778 vss 2.83e-19
C5159 vdd.n3779 vss 0.00311f
C5160 vdd.n3780 vss 4.25e-19
C5161 vdd.n3781 vss 0.00423f
C5162 vdd.n3782 vss 2.92e-19
C5163 vdd.n3783 vss 0.00521f
C5164 vdd.n3784 vss 0.00538f
C5165 vdd.n3785 vss 0.00868f
C5166 vdd.n3786 vss 0.0035f
C5167 vdd.n3787 vss -0.189f
C5168 vdd.n3788 vss 0.00524f
C5169 vdd.n3789 vss 0.00722f
C5170 vdd.n3790 vss 0.00594f
C5171 vdd.n3791 vss 0.00297f
C5172 vdd.n3792 vss 0.00877f
C5173 vdd.n3793 vss 0.00877f
C5174 vdd.n3794 vss 0.0115f
C5175 vdd.n3796 vss 0.00933f
C5176 vdd.n3797 vss 2.83e-19
C5177 vdd.n3798 vss 0.00311f
C5178 vdd.n3799 vss 4.25e-19
C5179 vdd.n3800 vss 0.00423f
C5180 vdd.n3801 vss 2.92e-19
C5181 vdd.n3802 vss 0.00521f
C5182 vdd.n3803 vss 0.00538f
C5183 vdd.n3804 vss 0.00868f
C5184 vdd.n3805 vss 0.0035f
C5185 vdd.n3806 vss 0.00437f
C5186 vdd.n3807 vss 0.00524f
C5187 vdd.n3808 vss 0.00722f
C5188 vdd.n3809 vss 0.00594f
C5189 vdd.n3810 vss 0.00297f
C5190 vdd.n3811 vss 0.00877f
C5191 vdd.n3812 vss 0.00877f
C5192 vdd.n3813 vss 0.0115f
C5193 vdd.n3815 vss 0.00933f
C5194 vdd.n3816 vss 2.83e-19
C5195 vdd.n3817 vss 0.00311f
C5196 vdd.n3818 vss 4.25e-19
C5197 vdd.n3819 vss 0.00423f
C5198 vdd.n3820 vss 2.92e-19
C5199 vdd.n3821 vss -0.077f
C5200 vdd.n3822 vss 0.00538f
C5201 vdd.n3823 vss 0.0116f
C5202 vdd.n3824 vss 0.0238f
C5203 vdd.n3825 vss 0.00573f
C5204 vdd.n3826 vss 0.00687f
C5205 vdd.n3827 vss 0.00437f
C5206 vdd.n3828 vss 0.00698f
C5207 vdd.n3829 vss 0.0109f
C5208 vdd.n3830 vss 0.00553f
C5209 vdd.n3831 vss 0.00996f
C5210 vdd.n3832 vss 9.51e-19
C5211 vdd.n3833 vss 0.00664f
C5212 vdd.n3834 vss 3.74f
C5213 x4.x5[7].floating.n0 vss -7.99f
C5214 x4.x5[7].floating.n1 vss -28.9f
C5215 x4.x5[7].floating.n2 vss 3.83f
C5216 x4.x5[7].floating.n3 vss -7.07f
C5217 x4.x5[7].floating.n4 vss -28.3f
C5218 x4.x5[7].floating.n5 vss 52.7f
C5219 x4.x5[7].floating.n6 vss -28.3f
C5220 x4.x5[7].floating.n7 vss -7.07f
C5221 x4.x5[7].floating.n8 vss 3.83f
C5222 x4.x5[7].floating.n9 vss -28.9f
C5223 x4.x5[7].floating.n10 vss -8.01f
C5224 x4.x5[7].floating.n11 vss 2.21f
C5225 x4.x5[7].floating.t1 vss 0.859f
C5226 x4.x5[7].floating.n12 vss 6.65f
C5227 x4.x5[7].floating.n13 vss 1.21f
C5228 x4.x5[7].floating.n14 vss 1.17f
C5229 x4.x5[7].floating.n15 vss 2.18f
C5230 x4.x5[7].floating.n16 vss 1.06f
C5231 x4.x5[7].floating.n17 vss 0.366f
C5232 x4.x5[7].floating.n18 vss 1.06f
C5233 x4.x5[7].floating.n19 vss 2.8f
C5234 x4.x5[7].floating.n20 vss 51.4f
C5235 x4.x5[7].floating.n21 vss 2.79f
C5236 x4.x5[7].floating.n22 vss 1.06f
C5237 x4.x5[7].floating.n23 vss 0.364f
C5238 x4.x5[7].floating.t7 vss 0.859f
C5239 x4.x5[7].floating.n24 vss 6.48f
C5240 x4.x5[7].floating.n25 vss 1.15f
C5241 x4.x5[7].floating.n26 vss 1.36f
C5242 x4.x5[7].floating.n27 vss 2.2f
C5243 x4.x5[7].floating.n28 vss 1.06f
C5244 x4.x5[7].floating.n29 vss 2.23f
C5245 x4.x5[7].floating.n30 vss -7.99f
C5246 x4.x5[7].floating.n31 vss -28.9f
C5247 x4.x5[7].floating.n32 vss 3.83f
C5248 x4.x5[7].floating.n33 vss -7.07f
C5249 x4.x5[7].floating.n34 vss -28.3f
C5250 x4.x5[7].floating.n35 vss 52.7f
C5251 x4.x5[7].floating.n36 vss -28.3f
C5252 x4.x5[7].floating.n37 vss -7.07f
C5253 x4.x5[7].floating.n38 vss 3.83f
C5254 x4.x5[7].floating.n39 vss -28.9f
C5255 x4.x5[7].floating.n40 vss -8.01f
C5256 x4.x5[7].floating.n41 vss 2.21f
C5257 x4.x5[7].floating.t6 vss 0.859f
C5258 x4.x5[7].floating.n42 vss 6.65f
C5259 x4.x5[7].floating.n43 vss 1.21f
C5260 x4.x5[7].floating.n44 vss 1.17f
C5261 x4.x5[7].floating.n45 vss 2.18f
C5262 x4.x5[7].floating.n46 vss 1.06f
C5263 x4.x5[7].floating.n47 vss 0.366f
C5264 x4.x5[7].floating.n48 vss 1.06f
C5265 x4.x5[7].floating.n49 vss 2.8f
C5266 x4.x5[7].floating.n50 vss 51.4f
C5267 x4.x5[7].floating.n51 vss 2.79f
C5268 x4.x5[7].floating.n52 vss 1.06f
C5269 x4.x5[7].floating.n53 vss 0.364f
C5270 x4.x5[7].floating.t4 vss 0.859f
C5271 x4.x5[7].floating.n54 vss 6.48f
C5272 x4.x5[7].floating.n55 vss 1.15f
C5273 x4.x5[7].floating.n56 vss 1.36f
C5274 x4.x5[7].floating.n57 vss 2.2f
C5275 x4.x5[7].floating.n58 vss 1.06f
C5276 x4.x5[7].floating.n59 vss 2.23f
C5277 x4.x5[7].floating.n60 vss -7.99f
C5278 x4.x5[7].floating.n61 vss -28.9f
C5279 x4.x5[7].floating.n62 vss 3.83f
C5280 x4.x5[7].floating.n63 vss -7.07f
C5281 x4.x5[7].floating.n64 vss -28.3f
C5282 x4.x5[7].floating.n65 vss 52.7f
C5283 x4.x5[7].floating.n66 vss -28.3f
C5284 x4.x5[7].floating.n67 vss -7.07f
C5285 x4.x5[7].floating.n68 vss 3.83f
C5286 x4.x5[7].floating.n69 vss -28.9f
C5287 x4.x5[7].floating.n70 vss -8.01f
C5288 x4.x5[7].floating.n71 vss 2.21f
C5289 x4.x5[7].floating.t3 vss 0.859f
C5290 x4.x5[7].floating.n72 vss 6.65f
C5291 x4.x5[7].floating.n73 vss 1.21f
C5292 x4.x5[7].floating.n74 vss 1.17f
C5293 x4.x5[7].floating.n75 vss 2.18f
C5294 x4.x5[7].floating.n76 vss 1.06f
C5295 x4.x5[7].floating.n77 vss 0.366f
C5296 x4.x5[7].floating.n78 vss 1.06f
C5297 x4.x5[7].floating.n79 vss 2.8f
C5298 x4.x5[7].floating.n80 vss 51.4f
C5299 x4.x5[7].floating.n81 vss 2.79f
C5300 x4.x5[7].floating.n82 vss 1.06f
C5301 x4.x5[7].floating.n83 vss 0.364f
C5302 x4.x5[7].floating.t0 vss 0.859f
C5303 x4.x5[7].floating.n84 vss 6.48f
C5304 x4.x5[7].floating.n85 vss 1.15f
C5305 x4.x5[7].floating.n86 vss 1.36f
C5306 x4.x5[7].floating.n87 vss 2.2f
C5307 x4.x5[7].floating.n88 vss 1.06f
C5308 x4.x5[7].floating.n89 vss -15.2f
C5309 x4.x5[7].floating.n90 vss -15.2f
C5310 x4.x5[7].floating.n91 vss -41.6f
C5311 x4.x5[7].floating.n92 vss 0.766f
C5312 x4.x5[7].floating.n93 vss 2.47f
C5313 x4.x5[7].floating.n94 vss 51.5f
C5314 x4.x5[7].floating.n95 vss 2.47f
C5315 x4.x5[7].floating.n96 vss 0.766f
C5316 x4.x5[7].floating.n97 vss -33.5f
C5317 x4.x5[7].floating.n98 vss -4.56f
C5318 x4.x5[7].floating.n99 vss 3.83f
C5319 x4.x5[7].floating.n100 vss -28.9f
C5320 x4.x5[7].floating.n101 vss -7.07f
C5321 x4.x5[7].floating.n102 vss 2.68f
C5322 x4.x5[7].floating.n103 vss 52f
C5323 x4.x5[7].floating.n104 vss 3.23f
C5324 x4.x5[7].floating.n105 vss -7.84f
C5325 x4.x5[7].floating.n106 vss -28.9f
C5326 x4.x5[7].floating.n107 vss 3.83f
C5327 x4.x5[7].floating.n108 vss -5.01f
C5328 x4.x5[7].floating.n109 vss -33f
C5329 x4.x5[7].floating.n110 vss 0.766f
C5330 x4.x5[7].floating.n111 vss 2.47f
C5331 x4.x5[7].floating.n112 vss 51.5f
C5332 x4.x5[7].floating.n113 vss 2.47f
C5333 x4.x5[7].floating.n114 vss 0.766f
C5334 x4.x5[7].floating.n115 vss -33.5f
C5335 x4.x5[7].floating.n116 vss -4.56f
C5336 x4.x5[7].floating.n117 vss 3.83f
C5337 x4.x5[7].floating.n118 vss -28.9f
C5338 x4.x5[7].floating.n119 vss -7.07f
C5339 x4.x5[7].floating.n120 vss 2.68f
C5340 x4.x5[7].floating.n121 vss 52f
C5341 x4.x5[7].floating.n122 vss 3.23f
C5342 x4.x5[7].floating.n123 vss -7.84f
C5343 x4.x5[7].floating.n124 vss -28.9f
C5344 x4.x5[7].floating.n125 vss 3.83f
C5345 x4.x5[7].floating.n126 vss -5.01f
C5346 x4.x5[7].floating.n127 vss -33f
C5347 x4.x5[7].floating.n128 vss 0.766f
C5348 x4.x5[7].floating.n129 vss 2.47f
C5349 x4.x5[7].floating.n130 vss 51.5f
C5350 x4.x5[7].floating.n131 vss 2.47f
C5351 x4.x5[7].floating.n132 vss 0.766f
C5352 x4.x5[7].floating.n133 vss -33.5f
C5353 x4.x5[7].floating.n134 vss -4.56f
C5354 x4.x5[7].floating.n135 vss 3.83f
C5355 x4.x5[7].floating.n136 vss -28.9f
C5356 x4.x5[7].floating.n137 vss -7.07f
C5357 x4.x5[7].floating.n138 vss 2.68f
C5358 x4.x5[7].floating.n139 vss 52f
C5359 x4.x5[7].floating.n140 vss 3.23f
C5360 x4.x5[7].floating.n141 vss 2.23f
C5361 x4.x5[7].floating.t2 vss 0.859f
C5362 x4.x5[7].floating.n142 vss 6.48f
C5363 x4.x5[7].floating.n143 vss 1.15f
C5364 x4.x5[7].floating.n144 vss 1.36f
C5365 x4.x5[7].floating.n145 vss 2.2f
C5366 x4.x5[7].floating.n146 vss 1.06f
C5367 x4.x5[7].floating.n147 vss 0.364f
C5368 x4.x5[7].floating.n148 vss 1.06f
C5369 x4.x5[7].floating.n149 vss 2.79f
C5370 x4.x5[7].floating.n150 vss 51.4f
C5371 x4.x5[7].floating.n151 vss 2.8f
C5372 x4.x5[7].floating.n152 vss 1.06f
C5373 x4.x5[7].floating.n153 vss 0.366f
C5374 x4.x5[7].floating.t5 vss 0.859f
C5375 x4.x5[7].floating.n154 vss 7.16f
C5376 x4.x5[7].floating.n155 vss 1.21f
C5377 x4.x5[7].floating.n156 vss 1.17f
C5378 x4.x5[7].floating.n157 vss 1.67f
C5379 x4.x5[7].floating.n158 vss 1.06f
C5380 x4.x5[7].floating.n159 vss -17.4f
C5381 x4.x5[7].floating.n160 vss -17.2f
C5382 x4.x5[7].floating.n161 vss -43.6f
C5383 x4.x5[7].floating.n162 vss 0.766f
C5384 x4.x5[7].floating.n163 vss 2.47f
C5385 x4.x5[7].floating.n164 vss 51.5f
C5386 x4.x5[7].floating.n165 vss 2.47f
C5387 x4.x5[7].floating.n166 vss 0.766f
C5388 x4.x5[7].floating.n167 vss -33f
C5389 x4.x5[7].floating.n168 vss -5.01f
C5390 x4.x5[7].floating.n169 vss 3.83f
C5391 x4.x5[7].floating.n170 vss -28.9f
C5392 x4.x5[7].floating.n171 vss -7.84f
C5393 x4.x10.Y.t0 vss 0.0462f
C5394 x4.x10.Y.t9 vss 0.0167f
C5395 x4.x10.Y.t6 vss 0.0167f
C5396 x4.x10.Y.t5 vss 0.0167f
C5397 x4.x10.Y.t3 vss 0.0167f
C5398 x4.x10.Y.t2 vss 0.0167f
C5399 x4.x10.Y.t8 vss 0.0167f
C5400 x4.x10.Y.t7 vss 0.0167f
C5401 x4.x10.Y.t4 vss 0.0167f
C5402 x4.x10.Y.n0 vss 0.222f
C5403 x4.x10.Y.n1 vss 0.0366f
C5404 x4.x10.Y.t1 vss 0.0174f
C5405 x4.x10.Y.n2 vss 0.0188f
C5406 x4.x10.Y.n3 vss 0.0186f
C5407 x4.x10.Y.n4 vss 0.0151f
C5408 x4.x10.Y.n5 vss 0.0211f
.ends

