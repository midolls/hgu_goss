magic
tech sky130A
timestamp 1698045514
<< checkpaint >>
rect -630 -1630 730 730
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 SAMPLE_CLK
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 CLK
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 VDD
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 VSS
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 SET
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 RESET
port 5 nsew
<< end >>
