magic
tech sky130A
magscale 1 2
timestamp 1700648830
<< nwell >>
rect 511 1081 933 1603
<< pwell >>
rect 518 570 940 1074
<< nmos >>
rect 714 780 744 864
<< pmos >>
rect 707 1300 737 1384
<< ndiff >>
rect 656 852 714 864
rect 656 792 668 852
rect 702 792 714 852
rect 656 780 714 792
rect 744 852 802 864
rect 744 792 756 852
rect 790 792 802 852
rect 744 780 802 792
<< pdiff >>
rect 649 1372 707 1384
rect 649 1312 661 1372
rect 695 1312 707 1372
rect 649 1300 707 1312
rect 737 1372 795 1384
rect 737 1312 749 1372
rect 783 1312 795 1372
rect 737 1300 795 1312
<< ndiffc >>
rect 668 792 702 852
rect 756 792 790 852
<< pdiffc >>
rect 661 1312 695 1372
rect 749 1312 783 1372
<< psubdiff >>
rect 554 1004 650 1038
rect 808 1004 904 1038
rect 554 942 588 1004
rect 870 942 904 1004
rect 554 640 588 702
rect 870 640 904 702
rect 554 606 650 640
rect 808 606 904 640
<< nsubdiff >>
rect 547 1533 643 1567
rect 801 1533 897 1567
rect 547 1471 581 1533
rect 863 1471 897 1533
rect 547 1151 581 1213
rect 863 1151 897 1213
rect 547 1117 643 1151
rect 801 1117 897 1151
<< psubdiffcont >>
rect 650 1004 808 1038
rect 554 702 588 942
rect 870 702 904 942
rect 650 606 808 640
<< nsubdiffcont >>
rect 643 1533 801 1567
rect 547 1213 581 1471
rect 863 1213 897 1471
rect 643 1117 801 1151
<< poly >>
rect 707 1384 737 1414
rect 707 1269 737 1300
rect 689 1253 755 1269
rect 689 1219 705 1253
rect 739 1219 755 1253
rect 689 1203 755 1219
rect 696 936 762 952
rect 696 902 712 936
rect 746 902 762 936
rect 696 886 762 902
rect 714 864 744 886
rect 714 754 744 780
<< polycont >>
rect 705 1219 739 1253
rect 712 902 746 936
<< locali >>
rect 547 1533 643 1567
rect 801 1533 897 1567
rect 547 1471 581 1533
rect 660 1512 750 1533
rect 660 1382 696 1512
rect 863 1471 897 1533
rect 660 1380 695 1382
rect 661 1372 695 1380
rect 661 1296 695 1312
rect 749 1372 783 1388
rect 749 1296 783 1312
rect 689 1219 705 1253
rect 739 1219 755 1253
rect 547 1151 581 1213
rect 863 1151 897 1213
rect 547 1117 643 1151
rect 801 1117 897 1151
rect 554 1004 650 1038
rect 808 1004 904 1038
rect 554 942 588 1004
rect 870 942 904 1004
rect 696 902 712 936
rect 746 902 762 936
rect 554 640 588 702
rect 668 852 702 868
rect 668 716 702 792
rect 756 852 790 868
rect 756 776 790 792
rect 668 674 758 716
rect 700 640 758 674
rect 870 640 904 702
rect 554 606 650 640
rect 808 606 904 640
<< viali >>
rect 661 1312 695 1372
rect 749 1312 783 1372
rect 705 1219 739 1253
rect 712 902 746 936
rect 668 792 702 852
rect 756 792 790 852
<< metal1 >>
rect 655 1372 701 1384
rect 655 1312 661 1372
rect 695 1312 701 1372
rect 655 1300 701 1312
rect 743 1382 789 1384
rect 743 1372 816 1382
rect 743 1312 749 1372
rect 783 1312 828 1372
rect 743 1300 828 1312
rect 776 1298 828 1300
rect 693 1253 751 1259
rect 693 1232 705 1253
rect 692 1219 705 1232
rect 739 1232 751 1253
rect 739 1219 762 1232
rect 692 936 762 1219
rect 692 904 712 936
rect 700 902 712 904
rect 746 904 762 936
rect 746 902 758 904
rect 700 896 758 902
rect 790 864 828 1298
rect 662 852 708 864
rect 662 792 668 852
rect 702 792 708 852
rect 662 780 708 792
rect 750 852 828 864
rect 750 792 756 852
rect 790 792 828 852
rect 750 786 828 792
rect 750 780 796 786
<< labels >>
flabel metal1 692 904 762 1232 0 FreeSans 320 0 0 0 input
port 10 nsew
flabel metal1 790 786 828 1372 0 FreeSans 320 0 0 0 output
port 12 nsew
flabel locali 660 1382 696 1533 0 FreeSans 320 0 0 0 vdd
port 13 nsew
flabel locali 668 674 702 792 0 FreeSans 320 0 0 0 vss
port 15 nsew
<< end >>
