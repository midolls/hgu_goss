magic
tech sky130A
magscale 1 2
timestamp 1698241761
<< pwell >>
rect 320 1438 346 1470
rect 926 1438 952 1470
rect 320 416 346 448
rect 926 416 952 448
<< metal3 >>
rect 0 2110 1278 2112
rect 0 2046 104 2110
rect 168 2046 184 2110
rect 248 2046 264 2110
rect 328 2046 344 2110
rect 408 2046 424 2110
rect 488 2046 504 2110
rect 568 2046 710 2110
rect 774 2046 790 2110
rect 854 2046 870 2110
rect 934 2046 950 2110
rect 1014 2046 1030 2110
rect 1094 2046 1110 2110
rect 1174 2046 1278 2110
rect 0 2044 1278 2046
rect 0 1998 66 2044
rect 0 1934 1 1998
rect 65 1934 66 1998
rect 0 1918 66 1934
rect 0 1854 1 1918
rect 65 1854 66 1918
rect 0 1838 66 1854
rect 0 1774 1 1838
rect 65 1774 66 1838
rect 0 1758 66 1774
rect 0 1694 1 1758
rect 65 1694 66 1758
rect 0 1678 66 1694
rect 0 1614 1 1678
rect 65 1614 66 1678
rect 0 1598 66 1614
rect 0 1534 1 1598
rect 65 1534 66 1598
rect 0 1518 66 1534
rect 0 1454 1 1518
rect 65 1454 66 1518
rect 0 1438 66 1454
rect 0 1374 1 1438
rect 65 1374 66 1438
rect 0 1358 66 1374
rect 0 1294 1 1358
rect 65 1294 66 1358
rect 0 1278 66 1294
rect 0 1214 1 1278
rect 65 1214 66 1278
rect 0 1150 66 1214
rect 126 1150 186 2044
rect 246 1090 306 1984
rect 366 1150 426 2044
rect 606 1998 672 2044
rect 486 1090 546 1984
rect 606 1934 607 1998
rect 671 1934 672 1998
rect 606 1918 672 1934
rect 606 1854 607 1918
rect 671 1854 672 1918
rect 606 1838 672 1854
rect 606 1774 607 1838
rect 671 1774 672 1838
rect 606 1758 672 1774
rect 606 1694 607 1758
rect 671 1694 672 1758
rect 606 1678 672 1694
rect 606 1614 607 1678
rect 671 1614 672 1678
rect 606 1598 672 1614
rect 606 1534 607 1598
rect 671 1534 672 1598
rect 606 1518 672 1534
rect 606 1454 607 1518
rect 671 1454 672 1518
rect 606 1438 672 1454
rect 606 1374 607 1438
rect 671 1374 672 1438
rect 606 1358 672 1374
rect 606 1294 607 1358
rect 671 1294 672 1358
rect 606 1278 672 1294
rect 606 1214 607 1278
rect 671 1214 672 1278
rect 606 1150 672 1214
rect 732 1150 792 2044
rect 852 1090 912 1984
rect 972 1150 1032 2044
rect 1212 1998 1278 2044
rect 1092 1090 1152 1984
rect 1212 1934 1213 1998
rect 1277 1934 1278 1998
rect 1212 1918 1278 1934
rect 1212 1854 1213 1918
rect 1277 1854 1278 1918
rect 1212 1838 1278 1854
rect 1212 1774 1213 1838
rect 1277 1774 1278 1838
rect 1212 1758 1278 1774
rect 1212 1694 1213 1758
rect 1277 1694 1278 1758
rect 1212 1678 1278 1694
rect 1212 1614 1213 1678
rect 1277 1614 1278 1678
rect 1212 1598 1278 1614
rect 1212 1534 1213 1598
rect 1277 1534 1278 1598
rect 1212 1518 1278 1534
rect 1212 1454 1213 1518
rect 1277 1454 1278 1518
rect 1212 1438 1278 1454
rect 1212 1374 1213 1438
rect 1277 1374 1278 1438
rect 1212 1358 1278 1374
rect 1212 1294 1213 1358
rect 1277 1294 1278 1358
rect 1212 1278 1278 1294
rect 1212 1214 1213 1278
rect 1277 1214 1278 1278
rect 1212 1150 1278 1214
rect 0 1088 1278 1090
rect 0 1024 104 1088
rect 168 1024 184 1088
rect 248 1024 264 1088
rect 328 1024 344 1088
rect 408 1024 424 1088
rect 488 1024 504 1088
rect 568 1024 710 1088
rect 774 1024 790 1088
rect 854 1024 870 1088
rect 934 1024 950 1088
rect 1014 1024 1030 1088
rect 1094 1024 1110 1088
rect 1174 1024 1278 1088
rect 0 1022 1278 1024
rect 0 976 66 1022
rect 0 912 1 976
rect 65 912 66 976
rect 0 896 66 912
rect 0 832 1 896
rect 65 832 66 896
rect 0 816 66 832
rect 0 752 1 816
rect 65 752 66 816
rect 0 736 66 752
rect 0 672 1 736
rect 65 672 66 736
rect 0 656 66 672
rect 0 592 1 656
rect 65 592 66 656
rect 0 576 66 592
rect 0 512 1 576
rect 65 512 66 576
rect 0 496 66 512
rect 0 432 1 496
rect 65 432 66 496
rect 0 416 66 432
rect 0 352 1 416
rect 65 352 66 416
rect 0 336 66 352
rect 0 272 1 336
rect 65 272 66 336
rect 0 256 66 272
rect 0 192 1 256
rect 65 192 66 256
rect 0 128 66 192
rect 126 128 186 1022
rect 246 68 306 962
rect 366 128 426 1022
rect 606 976 672 1022
rect 486 68 546 962
rect 606 912 607 976
rect 671 912 672 976
rect 606 896 672 912
rect 606 832 607 896
rect 671 832 672 896
rect 606 816 672 832
rect 606 752 607 816
rect 671 752 672 816
rect 606 736 672 752
rect 606 672 607 736
rect 671 672 672 736
rect 606 656 672 672
rect 606 592 607 656
rect 671 592 672 656
rect 606 576 672 592
rect 606 512 607 576
rect 671 512 672 576
rect 606 496 672 512
rect 606 432 607 496
rect 671 432 672 496
rect 606 416 672 432
rect 606 352 607 416
rect 671 352 672 416
rect 606 336 672 352
rect 606 272 607 336
rect 671 272 672 336
rect 606 256 672 272
rect 606 192 607 256
rect 671 192 672 256
rect 606 128 672 192
rect 732 128 792 1022
rect 852 68 912 962
rect 972 128 1032 1022
rect 1212 976 1278 1022
rect 1092 68 1152 962
rect 1212 912 1213 976
rect 1277 912 1278 976
rect 1212 896 1278 912
rect 1212 832 1213 896
rect 1277 832 1278 896
rect 1212 816 1278 832
rect 1212 752 1213 816
rect 1277 752 1278 816
rect 1212 736 1278 752
rect 1212 672 1213 736
rect 1277 672 1278 736
rect 1212 656 1278 672
rect 1212 592 1213 656
rect 1277 592 1278 656
rect 1212 576 1278 592
rect 1212 512 1213 576
rect 1277 512 1278 576
rect 1212 496 1278 512
rect 1212 432 1213 496
rect 1277 432 1278 496
rect 1212 416 1278 432
rect 1212 352 1213 416
rect 1277 352 1278 416
rect 1212 336 1278 352
rect 1212 272 1213 336
rect 1277 272 1278 336
rect 1212 256 1278 272
rect 1212 192 1213 256
rect 1277 192 1278 256
rect 1212 128 1278 192
rect 126 66 1152 68
rect 126 2 184 66
rect 248 2 264 66
rect 328 2 344 66
rect 408 2 424 66
rect 488 2 790 66
rect 854 2 870 66
rect 934 2 950 66
rect 1014 2 1030 66
rect 1094 2 1152 66
rect 126 0 1152 2
<< via3 >>
rect 104 2046 168 2110
rect 184 2046 248 2110
rect 264 2046 328 2110
rect 344 2046 408 2110
rect 424 2046 488 2110
rect 504 2046 568 2110
rect 710 2046 774 2110
rect 790 2046 854 2110
rect 870 2046 934 2110
rect 950 2046 1014 2110
rect 1030 2046 1094 2110
rect 1110 2046 1174 2110
rect 1 1934 65 1998
rect 1 1854 65 1918
rect 1 1774 65 1838
rect 1 1694 65 1758
rect 1 1614 65 1678
rect 1 1534 65 1598
rect 1 1454 65 1518
rect 1 1374 65 1438
rect 1 1294 65 1358
rect 1 1214 65 1278
rect 607 1934 671 1998
rect 607 1854 671 1918
rect 607 1774 671 1838
rect 607 1694 671 1758
rect 607 1614 671 1678
rect 607 1534 671 1598
rect 607 1454 671 1518
rect 607 1374 671 1438
rect 607 1294 671 1358
rect 607 1214 671 1278
rect 1213 1934 1277 1998
rect 1213 1854 1277 1918
rect 1213 1774 1277 1838
rect 1213 1694 1277 1758
rect 1213 1614 1277 1678
rect 1213 1534 1277 1598
rect 1213 1454 1277 1518
rect 1213 1374 1277 1438
rect 1213 1294 1277 1358
rect 1213 1214 1277 1278
rect 104 1024 168 1088
rect 184 1024 248 1088
rect 264 1024 328 1088
rect 344 1024 408 1088
rect 424 1024 488 1088
rect 504 1024 568 1088
rect 710 1024 774 1088
rect 790 1024 854 1088
rect 870 1024 934 1088
rect 950 1024 1014 1088
rect 1030 1024 1094 1088
rect 1110 1024 1174 1088
rect 1 912 65 976
rect 1 832 65 896
rect 1 752 65 816
rect 1 672 65 736
rect 1 592 65 656
rect 1 512 65 576
rect 1 432 65 496
rect 1 352 65 416
rect 1 272 65 336
rect 1 192 65 256
rect 607 912 671 976
rect 607 832 671 896
rect 607 752 671 816
rect 607 672 671 736
rect 607 592 671 656
rect 607 512 671 576
rect 607 432 671 496
rect 607 352 671 416
rect 607 272 671 336
rect 607 192 671 256
rect 1213 912 1277 976
rect 1213 832 1277 896
rect 1213 752 1277 816
rect 1213 672 1277 736
rect 1213 592 1277 656
rect 1213 512 1277 576
rect 1213 432 1277 496
rect 1213 352 1277 416
rect 1213 272 1277 336
rect 1213 192 1277 256
rect 184 2 248 66
rect 264 2 328 66
rect 344 2 408 66
rect 424 2 488 66
rect 790 2 854 66
rect 870 2 934 66
rect 950 2 1014 66
rect 1030 2 1094 66
<< metal4 >>
rect 0 2110 1278 2112
rect 0 2046 104 2110
rect 168 2046 184 2110
rect 248 2046 264 2110
rect 328 2046 344 2110
rect 408 2046 424 2110
rect 488 2046 504 2110
rect 568 2046 710 2110
rect 774 2046 790 2110
rect 854 2046 870 2110
rect 934 2046 950 2110
rect 1014 2046 1030 2110
rect 1094 2046 1110 2110
rect 1174 2046 1278 2110
rect 0 2044 1278 2046
rect 0 1998 66 2044
rect 0 1934 1 1998
rect 65 1934 66 1998
rect 0 1918 66 1934
rect 0 1854 1 1918
rect 65 1854 66 1918
rect 0 1838 66 1854
rect 0 1774 1 1838
rect 65 1774 66 1838
rect 0 1758 66 1774
rect 0 1694 1 1758
rect 65 1694 66 1758
rect 0 1678 66 1694
rect 0 1614 1 1678
rect 65 1614 66 1678
rect 0 1598 66 1614
rect 0 1534 1 1598
rect 65 1534 66 1598
rect 0 1518 66 1534
rect 0 1454 1 1518
rect 65 1454 66 1518
rect 0 1438 66 1454
rect 0 1374 1 1438
rect 65 1374 66 1438
rect 0 1358 66 1374
rect 0 1294 1 1358
rect 65 1294 66 1358
rect 0 1278 66 1294
rect 0 1214 1 1278
rect 65 1214 66 1278
rect 0 1150 66 1214
rect 126 1090 186 1984
rect 246 1150 306 2044
rect 366 1090 426 1984
rect 486 1150 546 2044
rect 606 1998 672 2044
rect 606 1934 607 1998
rect 671 1934 672 1998
rect 606 1918 672 1934
rect 606 1854 607 1918
rect 671 1854 672 1918
rect 606 1838 672 1854
rect 606 1774 607 1838
rect 671 1774 672 1838
rect 606 1758 672 1774
rect 606 1694 607 1758
rect 671 1694 672 1758
rect 606 1678 672 1694
rect 606 1614 607 1678
rect 671 1614 672 1678
rect 606 1598 672 1614
rect 606 1534 607 1598
rect 671 1534 672 1598
rect 606 1518 672 1534
rect 606 1454 607 1518
rect 671 1454 672 1518
rect 606 1438 672 1454
rect 606 1374 607 1438
rect 671 1374 672 1438
rect 606 1358 672 1374
rect 606 1294 607 1358
rect 671 1294 672 1358
rect 606 1278 672 1294
rect 606 1214 607 1278
rect 671 1214 672 1278
rect 606 1150 672 1214
rect 732 1090 792 1984
rect 852 1150 912 2044
rect 972 1090 1032 1984
rect 1092 1150 1152 2044
rect 1212 1998 1278 2044
rect 1212 1934 1213 1998
rect 1277 1934 1278 1998
rect 1212 1918 1278 1934
rect 1212 1854 1213 1918
rect 1277 1854 1278 1918
rect 1212 1838 1278 1854
rect 1212 1774 1213 1838
rect 1277 1774 1278 1838
rect 1212 1758 1278 1774
rect 1212 1694 1213 1758
rect 1277 1694 1278 1758
rect 1212 1678 1278 1694
rect 1212 1614 1213 1678
rect 1277 1614 1278 1678
rect 1212 1598 1278 1614
rect 1212 1534 1213 1598
rect 1277 1534 1278 1598
rect 1212 1518 1278 1534
rect 1212 1454 1213 1518
rect 1277 1454 1278 1518
rect 1212 1438 1278 1454
rect 1212 1374 1213 1438
rect 1277 1374 1278 1438
rect 1212 1358 1278 1374
rect 1212 1294 1213 1358
rect 1277 1294 1278 1358
rect 1212 1278 1278 1294
rect 1212 1214 1213 1278
rect 1277 1214 1278 1278
rect 1212 1150 1278 1214
rect 0 1088 1278 1090
rect 0 1024 104 1088
rect 168 1024 184 1088
rect 248 1024 264 1088
rect 328 1024 344 1088
rect 408 1024 424 1088
rect 488 1024 504 1088
rect 568 1024 710 1088
rect 774 1024 790 1088
rect 854 1024 870 1088
rect 934 1024 950 1088
rect 1014 1024 1030 1088
rect 1094 1024 1110 1088
rect 1174 1024 1278 1088
rect 0 1022 1278 1024
rect 0 976 66 1022
rect 0 912 1 976
rect 65 912 66 976
rect 0 896 66 912
rect 0 832 1 896
rect 65 832 66 896
rect 0 816 66 832
rect 0 752 1 816
rect 65 752 66 816
rect 0 736 66 752
rect 0 672 1 736
rect 65 672 66 736
rect 0 656 66 672
rect 0 592 1 656
rect 65 592 66 656
rect 0 576 66 592
rect 0 512 1 576
rect 65 512 66 576
rect 0 496 66 512
rect 0 432 1 496
rect 65 432 66 496
rect 0 416 66 432
rect 0 352 1 416
rect 65 352 66 416
rect 0 336 66 352
rect 0 272 1 336
rect 65 272 66 336
rect 0 256 66 272
rect 0 192 1 256
rect 65 192 66 256
rect 0 128 66 192
rect 126 68 186 962
rect 246 128 306 1022
rect 366 68 426 962
rect 486 128 546 1022
rect 606 976 672 1022
rect 606 912 607 976
rect 671 912 672 976
rect 606 896 672 912
rect 606 832 607 896
rect 671 832 672 896
rect 606 816 672 832
rect 606 752 607 816
rect 671 752 672 816
rect 606 736 672 752
rect 606 672 607 736
rect 671 672 672 736
rect 606 656 672 672
rect 606 592 607 656
rect 671 592 672 656
rect 606 576 672 592
rect 606 512 607 576
rect 671 512 672 576
rect 606 496 672 512
rect 606 432 607 496
rect 671 432 672 496
rect 606 416 672 432
rect 606 352 607 416
rect 671 352 672 416
rect 606 336 672 352
rect 606 272 607 336
rect 671 272 672 336
rect 606 256 672 272
rect 606 192 607 256
rect 671 192 672 256
rect 606 128 672 192
rect 732 68 792 962
rect 852 128 912 1022
rect 972 68 1032 962
rect 1092 128 1152 1022
rect 1212 976 1278 1022
rect 1212 912 1213 976
rect 1277 912 1278 976
rect 1212 896 1278 912
rect 1212 832 1213 896
rect 1277 832 1278 896
rect 1212 816 1278 832
rect 1212 752 1213 816
rect 1277 752 1278 816
rect 1212 736 1278 752
rect 1212 672 1213 736
rect 1277 672 1278 736
rect 1212 656 1278 672
rect 1212 592 1213 656
rect 1277 592 1278 656
rect 1212 576 1278 592
rect 1212 512 1213 576
rect 1277 512 1278 576
rect 1212 496 1278 512
rect 1212 432 1213 496
rect 1277 432 1278 496
rect 1212 416 1278 432
rect 1212 352 1213 416
rect 1277 352 1278 416
rect 1212 336 1278 352
rect 1212 272 1213 336
rect 1277 272 1278 336
rect 1212 256 1278 272
rect 1212 192 1213 256
rect 1277 192 1278 256
rect 1212 128 1278 192
rect 126 66 1152 68
rect 126 2 184 66
rect 248 2 264 66
rect 328 2 344 66
rect 408 2 424 66
rect 488 2 790 66
rect 854 2 870 66
rect 934 2 950 66
rect 1014 2 1030 66
rect 1094 2 1152 66
rect 126 0 1152 2
<< labels >>
flabel space 926 1440 952 1472 0 FreeSans 160 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_0.SUB
flabel metal4 868 1772 894 1804 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_0.C1
flabel metal4 986 1182 1012 1214 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_0.C0
flabel space 926 418 952 450 0 FreeSans 160 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_1.SUB
flabel metal4 868 750 894 782 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_1.C1
flabel metal4 986 160 1012 192 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_0.hgu_cdac_unit_1.C0
flabel space 320 1440 346 1472 0 FreeSans 160 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_0.SUB
flabel metal4 262 1772 288 1804 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_0.C1
flabel metal4 380 1182 406 1214 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_0.C0
flabel space 320 418 346 450 0 FreeSans 160 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_1.SUB
flabel metal4 262 750 288 782 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C1
flabel metal4 380 160 406 192 0 FreeSans 320 0 0 0 hgu_cdac_cap_2_1.hgu_cdac_unit_1.C0
<< end >>
