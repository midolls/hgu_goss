* NGSPICE file created from hgu_tah_flat.ext - technology: sky130A

.subckt hgu_tah_flat sw VDD GND sw_n tah_vp vip vin tah_vn
X0 vip.t7 sw_n tah_vp.t8 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X1 tah_vn.t11 sw_n.t0 vin.t6 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X2 vin.t7 sw_n.t1 tah_vn.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X3 tah_vn.t2 sw.t0 tah_vn.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.908 ps=5.83 w=5.5 l=0.15
X4 vin.t4 sw_n.t2 tah_vn.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
X5 tah_vn.t8 sw_n.t3 vin.t5 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X6 tah_vn.t4 sw.t1 tah_vn.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0 ps=0 w=5.5 l=0.15
X7 tah_vp.t3 sw vip.t3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X8 tah_vp.t7 sw_n tah_vp.t7 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.454 ps=3.08 w=2.75 l=0.15
X9 tah_vn.t5 sw.t2 vin.t3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X10 tah_vp.t10 sw_n vip.t6 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X11 tah_vn.t7 sw_n.t4 tah_vn.t7 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.454 ps=3.08 w=2.75 l=0.15
X12 tah_vp.t2 sw tah_vp.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.908 ps=5.83 w=5.5 l=0.15
X13 vip.t2 sw tah_vp.t0 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.853 ps=6.12 w=2.75 l=0.15
X14 tah_vp.t5 sw vip.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X15 vin.t1 sw.t3 tah_vn.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.853 ps=6.12 w=2.75 l=0.15
X16 vip.t5 sw_n tah_vp.t11 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=1.71 ps=11.6 w=5.5 l=0.15
X17 tah_vn.t0 sw.t4 vin.t0 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X18 tah_vp.t9 sw_n vip.t4 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0.908 ps=5.83 w=5.5 l=0.15
X19 tah_vp.t6 sw_n tah_vp.t6 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0 ps=0 w=2.75 l=0.15
X20 tah_vn.t6 sw_n.t5 tah_vn.t6 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0 ps=0 w=2.75 l=0.15
X21 tah_vp.t1 sw tah_vp.t1 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.908 pd=5.83 as=0 ps=0 w=5.5 l=0.15
X22 vip.t0 sw tah_vp.t4 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
X23 vin.t2 sw.t5 tah_vn.t3 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.454 pd=3.08 as=0.454 ps=3.08 w=2.75 l=0.15
R0 sw_n.t5 sw_n.t4 1121.45
R1 sw_n.n2 sw_n.t2 1074.7
R2 sw_n.n3 sw_n.t1 925.441
R3 sw_n.n2 sw_n.t0 925.441
R4 sw_n.n4 sw_n.t3 925.441
R5 sw_n.t1 sw_n.n1 923.833
R6 sw_n sw_n.t5 582.713
R7 sw_n.n1 sw_n.n0 149.266
R8 sw_n.n4 sw_n.n3 149.266
R9 sw_n.n3 sw_n.n2 149.266
R10 sw_n sw_n.n4 67.8268
R11 tah_vp.n10 tah_vp.t0 8.79834
R12 tah_vp.n3 tah_vp.t11 8.25495
R13 tah_vp.n13 tah_vp.t6 7.20179
R14 tah_vp.n7 tah_vp.t7 7.2005
R15 tah_vp.n8 tah_vp.t5 7.2005
R16 tah_vp.n9 tah_vp.t4 7.2005
R17 tah_vp.n9 tah_vp.t3 7.2005
R18 tah_vp.n6 tah_vp.t1 5.91112
R19 tah_vp.n2 tah_vp.t8 5.9105
R20 tah_vp.n2 tah_vp.t10 5.9105
R21 tah_vp.n1 tah_vp.t9 5.9105
R22 tah_vp.n0 tah_vp.t2 5.9105
R23 tah_vp tah_vp.n6 2.79078
R24 tah_vp.n6 tah_vp.n5 1.99139
R25 tah_vp tah_vp.n13 1.77996
R26 tah_vp.n3 tah_vp.n2 1.63907
R27 tah_vp.n4 tah_vp.n1 1.63907
R28 tah_vp.n5 tah_vp.n0 1.63907
R29 tah_vp.n13 tah_vp.n12 1.24411
R30 tah_vp.n12 tah_vp.n7 0.892459
R31 tah_vp.n11 tah_vp.n8 0.892459
R32 tah_vp.n10 tah_vp.n9 0.892459
R33 tah_vp.n4 tah_vp.n3 0.706382
R34 tah_vp.n11 tah_vp.n10 0.706382
R35 tah_vp.n5 tah_vp.n4 0.353441
R36 tah_vp.n12 tah_vp.n11 0.353441
R37 vip.n4 vip.t3 7.2005
R38 vip.n4 vip.t2 7.2005
R39 vip.n3 vip.t1 7.2005
R40 vip.n3 vip.t0 7.2005
R41 vip.n1 vip.t4 5.9105
R42 vip.n1 vip.t7 5.9105
R43 vip.n0 vip.t6 5.9105
R44 vip.n0 vip.t5 5.9105
R45 vip.n2 vip.n1 1.95341
R46 vip.n2 vip.n0 1.94448
R47 vip.n5 vip.n3 1.20864
R48 vip.n5 vip.n4 1.20128
R49 vip vip.n2 0.706382
R50 vip vip.n5 0.695353
R51 VDD.n88 VDD.n84 68.0281
R52 VDD.n39 VDD.n36 67.9094
R53 VDD.n54 VDD.n51 66.2697
R54 VDD.n6 VDD.n3 66.2697
R55 VDD.n91 VDD.n90 42.9181
R56 VDD.n43 VDD.n42 42.9181
R57 VDD.n74 VDD.n73 36.1417
R58 VDD.n75 VDD.n74 36.1417
R59 VDD.n76 VDD.n75 36.1417
R60 VDD.n77 VDD.n76 36.1417
R61 VDD.n78 VDD.n77 36.1417
R62 VDD.n60 VDD.n56 36.1417
R63 VDD.n64 VDD.n60 36.1417
R64 VDD.n68 VDD.n64 36.1417
R65 VDD.n72 VDD.n68 36.1417
R66 VDD.n82 VDD.n72 36.1417
R67 VDD.n90 VDD.n82 36.1417
R68 VDD.n14 VDD.n13 36.1417
R69 VDD.n15 VDD.n14 36.1417
R70 VDD.n30 VDD.n29 36.1417
R71 VDD.n12 VDD.n8 36.1417
R72 VDD.n19 VDD.n12 36.1417
R73 VDD.n24 VDD.n19 36.1417
R74 VDD.n28 VDD.n24 36.1417
R75 VDD.n34 VDD.n28 36.1417
R76 VDD.n42 VDD.n34 36.1417
R77 VDD.n58 VDD.t3 29.3064
R78 VDD.n62 VDD.t0 29.3064
R79 VDD.n66 VDD.t7 29.3064
R80 VDD.n70 VDD.t9 29.3064
R81 VDD.n80 VDD.t10 29.3064
R82 VDD.n87 VDD.t8 29.3064
R83 VDD.n10 VDD.t1 29.3064
R84 VDD.n17 VDD.t2 29.3064
R85 VDD.n22 VDD.t4 29.3064
R86 VDD.n26 VDD.t11 29.3064
R87 VDD.n32 VDD.t6 29.3064
R88 VDD.n40 VDD.t5 29.3064
R89 VDD.n44 VDD.n43 6.00467
R90 VDD.n92 VDD.n91 5.78843
R91 VDD.n86 VDD.n85 0.267071
R92 VDD.n87 VDD.n86 0.267071
R93 VDD.n79 VDD.n78 0.267071
R94 VDD.n80 VDD.n79 0.267071
R95 VDD.n70 VDD.n69 0.267071
R96 VDD.n66 VDD.n65 0.267071
R97 VDD.n62 VDD.n61 0.267071
R98 VDD.n58 VDD.n57 0.267071
R99 VDD.n53 VDD.n52 0.267071
R100 VDD.n56 VDD.n55 0.267071
R101 VDD.n60 VDD.n59 0.267071
R102 VDD.n59 VDD.n58 0.267071
R103 VDD.n64 VDD.n63 0.267071
R104 VDD.n63 VDD.n62 0.267071
R105 VDD.n68 VDD.n67 0.267071
R106 VDD.n67 VDD.n66 0.267071
R107 VDD.n72 VDD.n71 0.267071
R108 VDD.n71 VDD.n70 0.267071
R109 VDD.n82 VDD.n81 0.267071
R110 VDD.n81 VDD.n80 0.267071
R111 VDD.n90 VDD.n89 0.267071
R112 VDD.n5 VDD.n4 0.267071
R113 VDD.n10 VDD.n9 0.267071
R114 VDD.n16 VDD.n15 0.267071
R115 VDD.n17 VDD.n16 0.267071
R116 VDD.n21 VDD.n20 0.267071
R117 VDD.n22 VDD.n21 0.267071
R118 VDD.n26 VDD.n25 0.267071
R119 VDD.n31 VDD.n30 0.267071
R120 VDD.n32 VDD.n31 0.267071
R121 VDD.n38 VDD.n37 0.267071
R122 VDD.n42 VDD.n41 0.267071
R123 VDD.n41 VDD.n40 0.267071
R124 VDD.n34 VDD.n33 0.267071
R125 VDD.n33 VDD.n32 0.267071
R126 VDD.n28 VDD.n27 0.267071
R127 VDD.n27 VDD.n26 0.267071
R128 VDD.n24 VDD.n23 0.267071
R129 VDD.n23 VDD.n22 0.267071
R130 VDD.n19 VDD.n18 0.267071
R131 VDD.n18 VDD.n17 0.267071
R132 VDD.n12 VDD.n11 0.267071
R133 VDD.n11 VDD.n10 0.267071
R134 VDD.n8 VDD.n7 0.267071
R135 VDD.n55 VDD.n54 0.261652
R136 VDD.n7 VDD.n6 0.261652
R137 VDD.n89 VDD.n88 0.26153
R138 VDD.n39 VDD.n38 0.261076
R139 VDD VDD.n47 0.257835
R140 VDD VDD.n95 0.205622
R141 VDD.n49 VDD.n48 0.0199714
R142 VDD.n46 VDD.n1 0.0199714
R143 VDD.n95 VDD.n94 0.00852938
R144 VDD.n40 VDD.n39 0.00771967
R145 VDD.n88 VDD.n87 0.00726749
R146 VDD.n54 VDD.n53 0.00689537
R147 VDD.n6 VDD.n5 0.00689537
R148 VDD.n84 VDD.n83 0.00407322
R149 VDD.n36 VDD.n35 0.00407322
R150 VDD.n51 VDD.n50 0.00407019
R151 VDD.n3 VDD.n2 0.00407019
R152 VDD.n94 VDD.n93 0.00200216
R153 VDD.n47 VDD.n46 0.00100125
R154 VDD.n93 VDD.n92 0.00100116
R155 VDD.n45 VDD.n44 0.00100116
R156 VDD.n46 VDD.n45 0.00100001
R157 VDD.n47 VDD.n0 0.00100001
R158 VDD.n93 VDD.n49 0.001
R159 vin.n0 vin.t0 7.2005
R160 vin.n0 vin.t2 7.2005
R161 vin.n1 vin.t3 7.2005
R162 vin.n1 vin.t1 7.2005
R163 vin.n4 vin.t5 5.9105
R164 vin.n4 vin.t7 5.9105
R165 vin.n3 vin.t6 5.9105
R166 vin.n3 vin.t4 5.9105
R167 vin.n5 vin.n4 1.95341
R168 vin.n5 vin.n3 1.94448
R169 vin.n2 vin.n0 1.20864
R170 vin.n2 vin.n1 1.20128
R171 vin vin.n5 0.728441
R172 vin vin.n2 0.673294
R173 tah_vn.n3 tah_vn.t1 8.79834
R174 tah_vn.n10 tah_vn.t9 8.25495
R175 tah_vn.n6 tah_vn.t6 7.20179
R176 tah_vn.n2 tah_vn.t3 7.2005
R177 tah_vn.n2 tah_vn.t5 7.2005
R178 tah_vn.n1 tah_vn.t0 7.2005
R179 tah_vn.n0 tah_vn.t7 7.2005
R180 tah_vn.n13 tah_vn.t4 5.91112
R181 tah_vn.n7 tah_vn.t2 5.9105
R182 tah_vn.n8 tah_vn.t8 5.9105
R183 tah_vn.n9 tah_vn.t10 5.9105
R184 tah_vn.n9 tah_vn.t11 5.9105
R185 tah_vn tah_vn.n13 2.57755
R186 tah_vn.n13 tah_vn.n12 1.99139
R187 tah_vn tah_vn.n6 1.90012
R188 tah_vn.n12 tah_vn.n7 1.63907
R189 tah_vn.n11 tah_vn.n8 1.63907
R190 tah_vn.n10 tah_vn.n9 1.63907
R191 tah_vn.n6 tah_vn.n5 1.24411
R192 tah_vn.n3 tah_vn.n2 0.892459
R193 tah_vn.n4 tah_vn.n1 0.892459
R194 tah_vn.n5 tah_vn.n0 0.892459
R195 tah_vn.n4 tah_vn.n3 0.706382
R196 tah_vn.n11 tah_vn.n10 0.706382
R197 tah_vn.n5 tah_vn.n4 0.353441
R198 tah_vn.n12 tah_vn.n11 0.353441
R199 sw.t1 sw.t0 2005.12
R200 sw sw.t1 965.894
R201 sw.n0 sw.t3 632.871
R202 sw.n2 sw.t4 483.608
R203 sw.n1 sw.t5 483.608
R204 sw.n0 sw.t2 483.608
R205 sw.n2 sw.n1 149.266
R206 sw.n1 sw.n0 149.266
R207 sw sw.n2 102.927
R208 VSS.n15 VSS.n11 660.529
R209 VSS.n60 VSS.n51 660.529
R210 VSS.n10 VSS.n7 156.236
R211 VSS.n10 VSS.n9 156.236
R212 VSS.n62 VSS.n1 156.236
R213 VSS.n62 VSS.n4 156.236
R214 VSS.n19 VSS.t4 108.531
R215 VSS.n30 VSS.t5 108.531
R216 VSS.n35 VSS.t1 108.531
R217 VSS.n40 VSS.t0 108.531
R218 VSS.n48 VSS.t3 108.531
R219 VSS.n59 VSS.t2 108.531
R220 VSS.n16 VSS.n10 42.9181
R221 VSS.n62 VSS.n61 42.9181
R222 VSS.n23 VSS.n22 36.1417
R223 VSS.n24 VSS.n23 36.1417
R224 VSS.n53 VSS.n52 36.1417
R225 VSS.n54 VSS.n53 36.1417
R226 VSS.n55 VSS.n54 36.1417
R227 VSS.n27 VSS.n26 36.1417
R228 VSS.n28 VSS.n27 36.1417
R229 VSS.n45 VSS.n44 36.1417
R230 VSS.n46 VSS.n45 36.1417
R231 VSS.n21 VSS.n16 36.1417
R232 VSS.n32 VSS.n21 36.1417
R233 VSS.n37 VSS.n32 36.1417
R234 VSS.n42 VSS.n37 36.1417
R235 VSS.n50 VSS.n42 36.1417
R236 VSS.n61 VSS.n50 36.1417
R237 VSS VSS.n62 2.25932
R238 VSS.n56 VSS.n55 0.843439
R239 VSS.n59 VSS.n56 0.843439
R240 VSS.n48 VSS.n43 0.843439
R241 VSS.n40 VSS.n38 0.843439
R242 VSS.n35 VSS.n33 0.843439
R243 VSS.n25 VSS.n24 0.843439
R244 VSS.n30 VSS.n25 0.843439
R245 VSS.n19 VSS.n17 0.843439
R246 VSS.n14 VSS.n12 0.843439
R247 VSS.n14 VSS.n13 0.843439
R248 VSS.n19 VSS.n18 0.843439
R249 VSS.n29 VSS.n28 0.843439
R250 VSS.n30 VSS.n29 0.843439
R251 VSS.n35 VSS.n34 0.843439
R252 VSS.n40 VSS.n39 0.843439
R253 VSS.n47 VSS.n46 0.843439
R254 VSS.n48 VSS.n47 0.843439
R255 VSS.n58 VSS.n57 0.843439
R256 VSS.n59 VSS.n58 0.843439
R257 VSS.n16 VSS.n15 0.843439
R258 VSS.n15 VSS.n14 0.843439
R259 VSS.n21 VSS.n20 0.843439
R260 VSS.n20 VSS.n19 0.843439
R261 VSS.n32 VSS.n31 0.843439
R262 VSS.n31 VSS.n30 0.843439
R263 VSS.n37 VSS.n36 0.843439
R264 VSS.n36 VSS.n35 0.843439
R265 VSS.n42 VSS.n41 0.843439
R266 VSS.n41 VSS.n40 0.843439
R267 VSS.n50 VSS.n49 0.843439
R268 VSS.n49 VSS.n48 0.843439
R269 VSS.n61 VSS.n60 0.843439
R270 VSS.n60 VSS.n59 0.843439
R271 VSS.n7 VSS.n6 0.0206266
R272 VSS.n6 VSS.n5 0.0206266
R273 VSS.n9 VSS.n8 0.0206266
R274 VSS.n1 VSS.n0 0.0206266
R275 VSS.n4 VSS.n3 0.0206266
R276 VSS.n3 VSS.n2 0.0206266
C0 tah_vp vip 5.1f
C1 VDD sw_n 1.24f
C2 VDD tah_vn 1.03f
C3 tah_vn vin 5.11f
C4 VDD tah_vp 1.03f
C5 sw sw_n 17.1f
.ends

