* NGSPICE file created from hgu_comp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_MQX2PY a_n73_n84# a_15_n84# a_n15_n115# w_n211_n303#
X0 a_15_n84# a_n15_n115# a_n73_n84# w_n211_n303# sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_9NW3WL a_n73_n84# a_15_n84# a_n15_n110# VSUBS
X0 a_15_n84# a_n15_n110# a_n73_n84# VSUBS sky130_fd_pr__nfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_MQP8BZ w_n311_n303# a_111_n84# a_n81_n84# a_n111_n129#
+ a_15_n84# a_n173_n84#
X0 a_15_n84# a_n111_n129# a_n81_n84# w_n311_n303# sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.139 ps=1.17 w=0.84 l=0.15
X1 a_n81_n84# a_n111_n129# a_n173_n84# w_n311_n303# sky130_fd_pr__pfet_01v8 ad=0.139 pd=1.17 as=0.26 ps=2.3 w=0.84 l=0.15
X2 a_111_n84# a_n111_n129# a_15_n84# w_n311_n303# sky130_fd_pr__pfet_01v8 ad=0.26 pd=2.3 as=0.139 ps=1.17 w=0.84 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_L7T3GD a_15_n42# a_n15_n68# a_n73_n42# VSUBS
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_PK34ES a_111_n46# a_n111_n72# a_n81_n46# a_15_n46#
+ a_n173_n46# VSUBS
X0 a_15_n46# a_n111_n72# a_n81_n46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.0759 ps=0.79 w=0.46 l=0.15
X1 a_111_n46# a_n111_n72# a_15_n46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.54 as=0.0759 ps=0.79 w=0.46 l=0.15
X2 a_n81_n46# a_n111_n72# a_n173_n46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0759 pd=0.79 as=0.143 ps=1.54 w=0.46 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_HNLS5R a_n159_n126# a_n129_n100# a_n221_n100# a_63_n100#
+ a_n33_n100# VSUBS
X0 a_n129_n100# a_n159_n126# a_n221_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1 a_63_n100# a_n159_n126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_n33_n100# a_n159_n126# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_159_n100# a_n159_n126# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z a_159_n100# a_n413_n100# a_255_n100# a_351_n100#
+ a_n129_n100# a_63_n100# a_n225_n100# a_n321_n100# a_n33_n100# a_n417_126# VSUBS
X0 a_63_n100# a_n417_126# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1 a_n33_n100# a_n417_126# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_351_n100# a_n417_126# a_255_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X3 a_159_n100# a_n417_126# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4 a_255_n100# a_n417_126# a_159_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_n321_n100# a_n417_126# a_n413_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X6 a_n225_n100# a_n417_126# a_n321_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7 a_n129_n100# a_n417_126# a_n225_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n15_n131#
X0 a_15_n100# a_n15_n131# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt hgu_comp cdac_vn cdac_vp comp_outp comp_outn clk VDD VSS
XXM12 VDD a_1716_n1348# a_1712_n8# VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM23 RS_p VSS a_1716_n1348# VSS sky130_fd_pr__nfet_01v8_9NW3WL
XXM34 VDD a_2060_n1456# RS_p VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM14 VDD a_534_n1522# a_534_n1522# a_1716_n1348# VDD VDD sky130_fd_pr__pfet_01v8_MQP8BZ
XXM13 a_1716_n1348# a_1712_n8# VSS VSS sky130_fd_pr__nfet_01v8_L7T3GD
XXM35 a_2060_n1456# RS_p VSS VSS sky130_fd_pr__nfet_01v8_L7T3GD
XXM36 VDD comp_outp comp_outp a_2060_n1456# VDD VDD sky130_fd_pr__pfet_01v8_MQP8BZ
XXM25 a_622_n1522# a_768_n1356# a_534_n1522# VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM24 a_768_n1356# a_534_n1522# a_622_n1522# VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM15 a_534_n1522# a_1716_n1348# a_534_n1522# VSS VSS VSS sky130_fd_pr__nfet_01v8_PK34ES
XXM26 XM27/a_15_n84# VSS a_622_n1522# VSS sky130_fd_pr__nfet_01v8_9NW3WL
XXM37 comp_outp a_2060_n1456# comp_outp VSS VSS VSS sky130_fd_pr__nfet_01v8_PK34ES
XXM27 a_768_n1356# XM27/a_15_n84# a_534_n1522# VSS sky130_fd_pr__nfet_01v8_9NW3WL
XXM16 RS_p VDD RS_n VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM17 VDD RS_n RS_p VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM28 VDD m1_864_n1556# a_768_n1356# VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM18 a_1040_n132# VDD a_1248_n152# VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM29 m1_864_n1556# a_768_n1356# VSS VSS sky130_fd_pr__nfet_01v8_L7T3GD
XXM19 VSS RS_n a_1040_n132# VSS sky130_fd_pr__nfet_01v8_9NW3WL
XXM1 clk VSS m1_594_n764# VSS m1_594_n764# VSS sky130_fd_pr__nfet_01v8_HNLS5R
XXM2 m1_594_n764# m1_594_n764# m1_690_n502# m1_594_n764# m1_690_n502# m1_690_n502#
+ m1_594_n764# m1_690_n502# m1_594_n764# cdac_vp VSS sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z
XXM3 m1_594_n764# m1_594_n764# m1_1842_n474# m1_594_n764# m1_1842_n474# m1_1842_n474#
+ m1_594_n764# m1_1842_n474# m1_594_n764# cdac_vn VSS sky130_fd_pr__nfet_01v8_lvt_Y5HS5Z
XXM4 m1_690_n502# a_1712_n8# a_1248_n152# VSS sky130_fd_pr__nfet_01v8_648S5X
XXM5 a_1248_n152# m1_1842_n474# a_1712_n8# VSS sky130_fd_pr__nfet_01v8_648S5X
XXM6 a_1712_n8# VDD VDD a_1248_n152# sky130_fd_pr__pfet_01v8_XGS3BL
XXM7 VDD a_1248_n152# VDD a_1712_n8# sky130_fd_pr__pfet_01v8_XGS3BL
XXM8 VDD a_1712_n8# VDD clk sky130_fd_pr__pfet_01v8_XGS3BL
XXM9 XM9/a_n73_n100# VDD VDD clk sky130_fd_pr__pfet_01v8_XGS3BL
XXM30 VDD a_1216_n1508# RS_n VDD sky130_fd_pr__pfet_01v8_MQX2PY
XXM20 a_1040_n132# a_1248_n152# VSS VSS sky130_fd_pr__nfet_01v8_L7T3GD
XXM31 a_1216_n1508# RS_n VSS VSS sky130_fd_pr__nfet_01v8_L7T3GD
XXM10 a_1248_n152# VDD VDD clk sky130_fd_pr__pfet_01v8_XGS3BL
XXM21 VDD a_622_n1522# a_622_n1522# a_1040_n132# VDD VDD sky130_fd_pr__pfet_01v8_MQP8BZ
XXM32 VDD comp_outn comp_outn a_1216_n1508# VDD VDD sky130_fd_pr__pfet_01v8_MQP8BZ
XXM11 VDD XM11/a_15_n100# VDD clk sky130_fd_pr__pfet_01v8_XGS3BL
XXM22 VSS a_1040_n132# VSS a_622_n1522# a_622_n1522# VSS sky130_fd_pr__nfet_01v8_PK34ES
XXM33 comp_outn a_1216_n1508# comp_outn VSS VSS VSS sky130_fd_pr__nfet_01v8_PK34ES
.ends

