* SPICE3 file created from ringoscill.ext - technology: sky130A

*.subckt ringoscill enable
Xx1 x5/Y x4/VGND VSUBS x5/VPB x4/VPWR x2/A sky130_fd_sc_hd__inv_2
Xx3 x3/A x4/VGND VSUBS x5/VPB x4/VPWR x4/A sky130_fd_sc_hd__inv_2
Xx2 x2/A x4/VGND VSUBS x5/VPB x4/VPWR x3/A sky130_fd_sc_hd__inv_2
Xx4 x4/A x4/VGND VSUBS x5/VPB x4/VPWR x5/B sky130_fd_sc_hd__inv_2
Xx5 enable x5/B x5/VGND VSUBS x5/VPB x5/VPWR x5/Y sky130_fd_sc_hd__nand2_1
*.ends
