** sch_path: /foss/designs/hgu_goss/hgu/tutorial/ringoscill.sch
**.subckt ringoscill enable out
*.ipin enable
*.opin out
x1 net1 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__inv_2
x2 net2 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_2
x3 net3 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_2
x4 net4 VGND VNB VPB VPWR out sky130_fd_sc_hd__inv_2
x5 enable out VGND VNB VPB VPWR net1 sky130_fd_sc_hd__nand2_1
**.ends
.end
