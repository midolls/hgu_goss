* NGSPICE file created from hgu_cdac_cap_4.ext - technology: sky130A

.subckt hgu_cdac_cap_4 CBOT CTOP SUB
C0 CBOT CTOP 20.3f
C1 CTOP SUB 1.95f
C2 CBOT SUB 2.64f
.ends

