magic
tech sky130A
timestamp 1699599968
<< checkpaint >>
rect -649 1202 1845 1226
rect -649 1178 2002 1202
rect -649 -354 2159 1178
rect -630 -402 2159 -354
rect -630 -1630 730 -402
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use sky130_fd_sc_hd__dfbbp_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699530450
transform 1 0 0 0 1 300
box -19 -24 1215 296
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 1215 0 1 276
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x4
timestamp 1697965495
transform 1 0 1372 0 1 252
box -19 -24 157 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 VSS
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 CLK
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 DIV_CLK
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 RESET
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 SET
port 5 nsew
<< end >>
