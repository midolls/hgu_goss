* NGSPICE file created from origin_state.ext - technology: sky130A

.subckt origin_state in out VSS VDD
X0 out.t0 x2.A VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 x2.A in.t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2 x2.A in.t1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3 out.t1 x2.A VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
R0 VSS.n0 VSS 1754.68
R1 VSS VSS.t0 1409.06
R2 VSS.t2 VSS 1409.06
R3 VSS.n1 VSS.n0 585
R4 VSS.n0 VSS.t2 505.137
R5 VSS.n6 VSS.t1 111.924
R6 VSS.n3 VSS.t3 111.924
R7 VSS.n10 VSS.n9 34.6358
R8 VSS.n4 VSS.n3 11.427
R9 VSS.n2 VSS.n1 6.89281
R10 VSS.n9 VSS.n6 6.77697
R11 VSS.n9 VSS.n8 4.6505
R12 VSS.n11 VSS.n10 4.6505
R13 VSS.n5 VSS.n2 4.6505
R14 VSS.n7 VSS 0.491331
R15 VSS.n8 VSS.n7 0.108749
R16 VSS.n11 VSS.n5 0.0979576
R17 VSS.n5 VSS.n4 0.0979576
R18 VSS VSS.n11 0.0492288
R19 VSS.n8 VSS 0.0185085
R20 VSS.n4 VSS 0.0185085
R21 out.n0 out.t1 137.917
R22 out out.t0 106.635
R23 out.n1 out 13.357
R24 out out.n1 5.56572
R25 out.n1 out 4.66888
R26 out out.n0 2.22659
R27 out.n0 out 1.55202
R28 in.n0 in.t0 230.502
R29 in.n0 in.t1 157.821
R30 in.n1 in.n0 8.66327
R31 in in.n1 3.61504
R32 in.n1 in 2.02684
R33 VDD.n10 VDD 366.325
R34 VDD VDD.t0 258.87
R35 VDD.t2 VDD 258.87
R36 VDD.n16 VDD.t1 158.06
R37 VDD.n2 VDD.t3 152.88
R38 VDD.n9 VDD.n8 50.5268
R39 VDD.n11 VDD.n10 39.0751
R40 VDD.n18 VDD.n17 34.6358
R41 VDD.n3 VDD.n2 20.8387
R42 VDD.n5 VDD.n4 9.3005
R43 VDD.n14 VDD.n13 9.3005
R44 VDD.n13 VDD.n12 9.3005
R45 VDD.n17 VDD.n16 8.28285
R46 VDD.n12 VDD.t2 7.32698
R47 VDD.n7 VDD.n6 6.02403
R48 VDD.n17 VDD.n1 4.6505
R49 VDD.n19 VDD.n18 4.6505
R50 VDD.n13 VDD.n9 3.15839
R51 VDD.n15 VDD.n14 3.1005
R52 VDD.n12 VDD.n11 2.44266
R53 VDD.n0 VDD 0.50103
R54 VDD.n14 VDD.n7 0.376971
R55 VDD.n1 VDD.n0 0.116584
R56 VDD.n19 VDD.n15 0.105045
R57 VDD.n5 VDD.n3 0.0857273
R58 VDD VDD.n19 0.0527727
R59 VDD VDD.n1 0.0198182
R60 VDD.n15 VDD.n5 0.0198182
R61 VDD.n3 VDD 0.0198182
.ends

