magic
tech sky130A
timestamp 1698147819
<< checkpaint >>
rect -630 -330 43302 1476
<< error_s >>
rect 1183 1857 1215 1858
rect 1223 1857 1255 1858
rect 1263 1857 1295 1858
rect 1303 1857 1335 1858
rect 1343 1857 1375 1858
rect 1546 1857 1578 1858
rect 1586 1857 1618 1858
rect 1626 1857 1658 1858
rect 1666 1857 1698 1858
rect 1706 1857 1738 1858
rect 1909 1857 1941 1858
rect 1949 1857 1981 1858
rect 1989 1857 2021 1858
rect 2029 1857 2061 1858
rect 2069 1857 2101 1858
rect 1162 1826 1394 1857
rect 1162 1825 1194 1826
rect 1202 1825 1234 1826
rect 1242 1825 1274 1826
rect 1282 1825 1314 1826
rect 1322 1825 1354 1826
rect 1362 1825 1394 1826
rect 1525 1826 1757 1857
rect 1525 1825 1557 1826
rect 1565 1825 1597 1826
rect 1605 1825 1637 1826
rect 1645 1825 1677 1826
rect 1685 1825 1717 1826
rect 1725 1825 1757 1826
rect 1888 1826 2120 1857
rect 1888 1825 1920 1826
rect 1928 1825 1960 1826
rect 1968 1825 2000 1826
rect 2008 1825 2040 1826
rect 2048 1825 2080 1826
rect 2088 1825 2120 1826
use save  hg
timestamp 1698132400
transform 1 0 46557 0 1 1100
box 343 298 739 758
use save  save_0
timestamp 1698132400
transform 1 0 47296 0 1 1100
box 343 298 739 758
use save  save_1
timestamp 1698132400
transform 1 0 48035 0 1 1100
box 343 298 739 758
use save  save_2
timestamp 1698132400
transform 1 0 48774 0 1 1100
box 343 298 739 758
use save  save_3
timestamp 1698132400
transform 1 0 49513 0 1 1100
box 343 298 739 758
use save  save_4
timestamp 1698132400
transform 1 0 50252 0 1 1100
box 343 298 739 758
use save  save_5
timestamp 1698132400
transform 1 0 50991 0 1 1100
box 343 298 739 758
use save  save_6
timestamp 1698132400
transform 1 0 51730 0 1 1100
box 343 298 739 758
use save  save_7
timestamp 1698132400
transform 1 0 52469 0 1 1100
box 343 298 739 758
use save  save_8
timestamp 1698132400
transform 1 0 53208 0 1 1100
box 343 298 739 758
use save  save_9
timestamp 1698132400
transform 1 0 53947 0 1 1100
box 343 298 739 758
use save  save_10
timestamp 1698132400
transform 1 0 54686 0 1 1100
box 343 298 739 758
use save  save_11
timestamp 1698132400
transform 1 0 55425 0 1 1100
box 343 298 739 758
use save  save_12
timestamp 1698132400
transform 1 0 56164 0 1 1100
box 343 298 739 758
use save  save_13
timestamp 1698132400
transform 1 0 56903 0 1 1100
box 343 298 739 758
use save  save_14
timestamp 1698132400
transform 1 0 57642 0 1 1100
box 343 298 739 758
use save  save_15
timestamp 1698132400
transform 1 0 58381 0 1 1100
box 343 298 739 758
use save  save_16
timestamp 1698132400
transform 1 0 59120 0 1 1100
box 343 298 739 758
use save  save_17
timestamp 1698132400
transform 1 0 59859 0 1 1100
box 343 298 739 758
use save  save_18
timestamp 1698132400
transform 1 0 60598 0 1 1100
box 343 298 739 758
use save  save_19
timestamp 1698132400
transform 1 0 61337 0 1 1100
box 343 298 739 758
use save  save_20
timestamp 1698132400
transform 1 0 62076 0 1 1100
box 343 298 739 758
use save  save_21
timestamp 1698132400
transform 1 0 62815 0 1 1100
box 343 298 739 758
use save  save_22
timestamp 1698132400
transform 1 0 63554 0 1 1100
box 343 298 739 758
use save  save_23
timestamp 1698132400
transform 1 0 64293 0 1 1100
box 343 298 739 758
use save  save_24
timestamp 1698132400
transform 1 0 65032 0 1 1100
box 343 298 739 758
use save  save_25
timestamp 1698132400
transform 1 0 65771 0 1 1100
box 343 298 739 758
use save  save_26
timestamp 1698132400
transform 1 0 66510 0 1 1100
box 343 298 739 758
use save  save_27
timestamp 1698132400
transform 1 0 67249 0 1 1100
box 343 298 739 758
use save  save_28
timestamp 1698132400
transform 1 0 67988 0 1 1100
box 343 298 739 758
use save  save_29
timestamp 1698132400
transform 1 0 68727 0 1 1100
box 343 298 739 758
use save  save_30
timestamp 1698132400
transform 1 0 69466 0 1 1100
box 343 298 739 758
use save  save_31
timestamp 1698132400
transform 1 0 70205 0 1 1100
box 343 298 739 758
use save  save_32
timestamp 1698132400
transform 1 0 70944 0 1 1100
box 343 298 739 758
use save  save_33
timestamp 1698132400
transform 1 0 71683 0 1 1100
box 343 298 739 758
use save  save_34
timestamp 1698132400
transform 1 0 72422 0 1 1100
box 343 298 739 758
use save  save_35
timestamp 1698132400
transform 1 0 73161 0 1 1100
box 343 298 739 758
use save  save_36
timestamp 1698132400
transform 1 0 73900 0 1 1100
box 343 298 739 758
use save  save_37
timestamp 1698132400
transform 1 0 74639 0 1 1100
box 343 298 739 758
use save  save_38
timestamp 1698132400
transform 1 0 75378 0 1 1100
box 343 298 739 758
use save  save_39
timestamp 1698132400
transform 1 0 76117 0 1 1100
box 343 298 739 758
use save  save_40
timestamp 1698132400
transform 1 0 76856 0 1 1100
box 343 298 739 758
use save  save_41
timestamp 1698132400
transform 1 0 77595 0 1 1100
box 343 298 739 758
use save  save_42
timestamp 1698132400
transform 1 0 78334 0 1 1100
box 343 298 739 758
use save  save_43
timestamp 1698132400
transform 1 0 79073 0 1 1100
box 343 298 739 758
use save  save_44
timestamp 1698132400
transform 1 0 79812 0 1 1100
box 343 298 739 758
use save  save_45
timestamp 1698132400
transform 1 0 80551 0 1 1100
box 343 298 739 758
use save  save_46
timestamp 1698132400
transform 1 0 81290 0 1 1100
box 343 298 739 758
use save  save_47
timestamp 1698132400
transform 1 0 82029 0 1 1100
box 343 298 739 758
use save  save_48
timestamp 1698132400
transform 1 0 82768 0 1 1100
box 343 298 739 758
use save  save_49
timestamp 1698132400
transform 1 0 83507 0 1 1100
box 343 298 739 758
use save  save_50
timestamp 1698132400
transform 1 0 84246 0 1 1100
box 343 298 739 758
use save  save_51
timestamp 1698132400
transform 1 0 84985 0 1 1100
box 343 298 739 758
use save  save_52
timestamp 1698132400
transform 1 0 85724 0 1 1100
box 343 298 739 758
use save  save_53
timestamp 1698132400
transform 1 0 86463 0 1 1100
box 343 298 739 758
use save  save_54
timestamp 1698132400
transform 1 0 87202 0 1 1100
box 343 298 739 758
use save  save_55
timestamp 1698132400
transform 1 0 87941 0 1 1100
box 343 298 739 758
use save  save_56
timestamp 1698132400
transform 1 0 88680 0 1 1100
box 343 298 739 758
use save  save_57
timestamp 1698132400
transform 1 0 89419 0 1 1100
box 343 298 739 758
use save  save_58
timestamp 1698132400
transform 1 0 90158 0 1 1100
box 343 298 739 758
use save  save_59
timestamp 1698132400
transform 1 0 90897 0 1 1100
box 343 298 739 758
use save  save_60
timestamp 1698132400
transform 1 0 91636 0 1 1100
box 343 298 739 758
use save  save_61
timestamp 1698132400
transform 1 0 92375 0 1 1100
box 343 298 739 758
use save  save_62
timestamp 1698132400
transform 1 0 93114 0 1 1100
box 343 298 739 758
use save  save_63
timestamp 1698132400
transform 1 0 22909 0 1 1100
box 343 298 739 758
use save  save_64
timestamp 1698132400
transform 1 0 23648 0 1 1100
box 343 298 739 758
use save  save_65
timestamp 1698132400
transform 1 0 24387 0 1 1100
box 343 298 739 758
use save  save_66
timestamp 1698132400
transform 1 0 25126 0 1 1100
box 343 298 739 758
use save  save_67
timestamp 1698132400
transform 1 0 25865 0 1 1100
box 343 298 739 758
use save  save_68
timestamp 1698132400
transform 1 0 26604 0 1 1100
box 343 298 739 758
use save  save_69
timestamp 1698132400
transform 1 0 27343 0 1 1100
box 343 298 739 758
use save  save_70
timestamp 1698132400
transform 1 0 28082 0 1 1100
box 343 298 739 758
use save  save_71
timestamp 1698132400
transform 1 0 28821 0 1 1100
box 343 298 739 758
use save  save_72
timestamp 1698132400
transform 1 0 29560 0 1 1100
box 343 298 739 758
use save  save_73
timestamp 1698132400
transform 1 0 30299 0 1 1100
box 343 298 739 758
use save  save_74
timestamp 1698132400
transform 1 0 31038 0 1 1100
box 343 298 739 758
use save  save_75
timestamp 1698132400
transform 1 0 31777 0 1 1100
box 343 298 739 758
use save  save_76
timestamp 1698132400
transform 1 0 32516 0 1 1100
box 343 298 739 758
use save  save_77
timestamp 1698132400
transform 1 0 33255 0 1 1100
box 343 298 739 758
use save  save_78
timestamp 1698132400
transform 1 0 33994 0 1 1100
box 343 298 739 758
use save  save_79
timestamp 1698132400
transform 1 0 34733 0 1 1100
box 343 298 739 758
use save  save_80
timestamp 1698132400
transform 1 0 35472 0 1 1100
box 343 298 739 758
use save  save_81
timestamp 1698132400
transform 1 0 36211 0 1 1100
box 343 298 739 758
use save  save_82
timestamp 1698132400
transform 1 0 36950 0 1 1100
box 343 298 739 758
use save  save_83
timestamp 1698132400
transform 1 0 37689 0 1 1100
box 343 298 739 758
use save  save_84
timestamp 1698132400
transform 1 0 38428 0 1 1100
box 343 298 739 758
use save  save_85
timestamp 1698132400
transform 1 0 39167 0 1 1100
box 343 298 739 758
use save  save_86
timestamp 1698132400
transform 1 0 39906 0 1 1100
box 343 298 739 758
use save  save_87
timestamp 1698132400
transform 1 0 40645 0 1 1100
box 343 298 739 758
use save  save_88
timestamp 1698132400
transform 1 0 41384 0 1 1100
box 343 298 739 758
use save  save_89
timestamp 1698132400
transform 1 0 42123 0 1 1100
box 343 298 739 758
use save  save_90
timestamp 1698132400
transform 1 0 42862 0 1 1100
box 343 298 739 758
use save  save_91
timestamp 1698132400
transform 1 0 43601 0 1 1100
box 343 298 739 758
use save  save_92
timestamp 1698132400
transform 1 0 44340 0 1 1100
box 343 298 739 758
use save  save_93
timestamp 1698132400
transform 1 0 45079 0 1 1100
box 343 298 739 758
use save  save_94
timestamp 1698132400
transform 1 0 45818 0 1 1100
box 343 298 739 758
use save  save_95
timestamp 1698132400
transform 1 0 11085 0 1 1100
box 343 298 739 758
use save  save_96
timestamp 1698132400
transform 1 0 11824 0 1 1100
box 343 298 739 758
use save  save_97
timestamp 1698132400
transform 1 0 12563 0 1 1100
box 343 298 739 758
use save  save_98
timestamp 1698132400
transform 1 0 13302 0 1 1100
box 343 298 739 758
use save  save_99
timestamp 1698132400
transform 1 0 14041 0 1 1100
box 343 298 739 758
use save  save_100
timestamp 1698132400
transform 1 0 14780 0 1 1100
box 343 298 739 758
use save  save_101
timestamp 1698132400
transform 1 0 15519 0 1 1100
box 343 298 739 758
use save  save_102
timestamp 1698132400
transform 1 0 16258 0 1 1100
box 343 298 739 758
use save  save_103
timestamp 1698132400
transform 1 0 16997 0 1 1100
box 343 298 739 758
use save  save_104
timestamp 1698132400
transform 1 0 17736 0 1 1100
box 343 298 739 758
use save  save_105
timestamp 1698132400
transform 1 0 18475 0 1 1100
box 343 298 739 758
use save  save_106
timestamp 1698132400
transform 1 0 19214 0 1 1100
box 343 298 739 758
use save  save_107
timestamp 1698132400
transform 1 0 19953 0 1 1100
box 343 298 739 758
use save  save_108
timestamp 1698132400
transform 1 0 20692 0 1 1100
box 343 298 739 758
use save  save_109
timestamp 1698132400
transform 1 0 21431 0 1 1100
box 343 298 739 758
use save  save_110
timestamp 1698132400
transform 1 0 22170 0 1 1100
box 343 298 739 758
use save  save_111
timestamp 1698132400
transform 1 0 -1407 0 1 255
box 343 298 739 758
use save  save_112
timestamp 1698132400
transform 1 0 -668 0 1 255
box 343 298 739 758
use save  save_113
timestamp 1698132400
transform 1 0 71 0 1 255
box 343 298 739 758
use save  save_114
timestamp 1698132400
transform 1 0 810 0 1 255
box 343 298 739 758
use save  save_115
timestamp 1698132400
transform 1 0 1549 0 1 255
box 343 298 739 758
use save  save_116
timestamp 1698132400
transform 1 0 2288 0 1 255
box 343 298 739 758
use save  save_117
timestamp 1698132400
transform 1 0 3034 0 1 233
box 343 298 739 758
use save  save_118
timestamp 1698132400
transform 1 0 10346 0 1 1100
box 343 298 739 758
use save  save_119
timestamp 1698132400
transform 1 0 1465 0 1 1100
box 343 298 739 758
use save  save_120
timestamp 1698132400
transform 1 0 1465 0 1 1526
box 343 298 739 758
use save  save_121
timestamp 1698132400
transform 1 0 1102 0 1 1100
box 343 298 739 758
use save  save_122
timestamp 1698132400
transform 1 0 1102 0 1 1526
box 343 298 739 758
use save  save_123
timestamp 1698132400
transform 1 0 739 0 1 1100
box 343 298 739 758
use save  save_124
timestamp 1698132400
transform 1 0 739 0 1 1526
box 343 298 739 758
use save  save_125
timestamp 1698132400
transform 1 0 376 0 1 1100
box 343 298 739 758
use hgu_cdac_unit  x1
timestamp 1698146599
transform 1 0 -343 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x2[0]
timestamp 1698146599
transform 1 0 329 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x2[1]
timestamp 1698146599
transform 1 0 -7 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x3[0]
timestamp 1698146599
transform 1 0 1673 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x3[1]
timestamp 1698146599
transform 1 0 1337 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x3[2]
timestamp 1698146599
transform 1 0 1001 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x3[3]
timestamp 1698146599
transform 1 0 665 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[0]
timestamp 1698146599
transform 1 0 4361 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[1]
timestamp 1698146599
transform 1 0 4025 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[2]
timestamp 1698146599
transform 1 0 3689 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[3]
timestamp 1698146599
transform 1 0 3353 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[4]
timestamp 1698146599
transform 1 0 3017 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[5]
timestamp 1698146599
transform 1 0 2681 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[6]
timestamp 1698146599
transform 1 0 2345 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x4[7]
timestamp 1698146599
transform 1 0 2009 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[0]
timestamp 1698146599
transform 1 0 9737 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[1]
timestamp 1698146599
transform 1 0 9401 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[2]
timestamp 1698146599
transform 1 0 9065 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[3]
timestamp 1698146599
transform 1 0 8729 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[4]
timestamp 1698146599
transform 1 0 8393 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[5]
timestamp 1698146599
transform 1 0 8057 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[6]
timestamp 1698146599
transform 1 0 7721 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[7]
timestamp 1698146599
transform 1 0 7385 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[8]
timestamp 1698146599
transform 1 0 7049 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[9]
timestamp 1698146599
transform 1 0 6713 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[10]
timestamp 1698146599
transform 1 0 6377 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[11]
timestamp 1698146599
transform 1 0 6041 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[12]
timestamp 1698146599
transform 1 0 5705 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[13]
timestamp 1698146599
transform 1 0 5369 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[14]
timestamp 1698146599
transform 1 0 5033 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x5[15]
timestamp 1698146599
transform 1 0 4697 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[0]
timestamp 1698146599
transform 1 0 20489 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[1]
timestamp 1698146599
transform 1 0 20153 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[2]
timestamp 1698146599
transform 1 0 19817 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[3]
timestamp 1698146599
transform 1 0 19481 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[4]
timestamp 1698146599
transform 1 0 19145 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[5]
timestamp 1698146599
transform 1 0 18809 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[6]
timestamp 1698146599
transform 1 0 18473 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[7]
timestamp 1698146599
transform 1 0 18137 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[8]
timestamp 1698146599
transform 1 0 17801 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[9]
timestamp 1698146599
transform 1 0 17465 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[10]
timestamp 1698146599
transform 1 0 17129 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[11]
timestamp 1698146599
transform 1 0 16793 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[12]
timestamp 1698146599
transform 1 0 16457 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[13]
timestamp 1698146599
transform 1 0 16121 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[14]
timestamp 1698146599
transform 1 0 15785 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[15]
timestamp 1698146599
transform 1 0 15449 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[16]
timestamp 1698146599
transform 1 0 15113 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[17]
timestamp 1698146599
transform 1 0 14777 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[18]
timestamp 1698146599
transform 1 0 14441 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[19]
timestamp 1698146599
transform 1 0 14105 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[20]
timestamp 1698146599
transform 1 0 13769 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[21]
timestamp 1698146599
transform 1 0 13433 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[22]
timestamp 1698146599
transform 1 0 13097 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[23]
timestamp 1698146599
transform 1 0 12761 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[24]
timestamp 1698146599
transform 1 0 12425 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[25]
timestamp 1698146599
transform 1 0 12089 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[26]
timestamp 1698146599
transform 1 0 11753 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[27]
timestamp 1698146599
transform 1 0 11417 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[28]
timestamp 1698146599
transform 1 0 11081 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[29]
timestamp 1698146599
transform 1 0 10745 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[30]
timestamp 1698146599
transform 1 0 10409 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x6[31]
timestamp 1698146599
transform 1 0 10073 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[0]
timestamp 1698146599
transform 1 0 41993 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[1]
timestamp 1698146599
transform 1 0 41657 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[2]
timestamp 1698146599
transform 1 0 41321 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[3]
timestamp 1698146599
transform 1 0 40985 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[4]
timestamp 1698146599
transform 1 0 40649 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[5]
timestamp 1698146599
transform 1 0 40313 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[6]
timestamp 1698146599
transform 1 0 39977 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[7]
timestamp 1698146599
transform 1 0 39641 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[8]
timestamp 1698146599
transform 1 0 39305 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[9]
timestamp 1698146599
transform 1 0 38969 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[10]
timestamp 1698146599
transform 1 0 38633 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[11]
timestamp 1698146599
transform 1 0 38297 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[12]
timestamp 1698146599
transform 1 0 37961 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[13]
timestamp 1698146599
transform 1 0 37625 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[14]
timestamp 1698146599
transform 1 0 37289 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[15]
timestamp 1698146599
transform 1 0 36953 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[16]
timestamp 1698146599
transform 1 0 36617 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[17]
timestamp 1698146599
transform 1 0 36281 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[18]
timestamp 1698146599
transform 1 0 35945 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[19]
timestamp 1698146599
transform 1 0 35609 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[20]
timestamp 1698146599
transform 1 0 35273 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[21]
timestamp 1698146599
transform 1 0 34937 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[22]
timestamp 1698146599
transform 1 0 34601 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[23]
timestamp 1698146599
transform 1 0 34265 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[24]
timestamp 1698146599
transform 1 0 33929 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[25]
timestamp 1698146599
transform 1 0 33593 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[26]
timestamp 1698146599
transform 1 0 33257 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[27]
timestamp 1698146599
transform 1 0 32921 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[28]
timestamp 1698146599
transform 1 0 32585 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[29]
timestamp 1698146599
transform 1 0 32249 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[30]
timestamp 1698146599
transform 1 0 31913 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[31]
timestamp 1698146599
transform 1 0 31577 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[32]
timestamp 1698146599
transform 1 0 31241 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[33]
timestamp 1698146599
transform 1 0 30905 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[34]
timestamp 1698146599
transform 1 0 30569 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[35]
timestamp 1698146599
transform 1 0 30233 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[36]
timestamp 1698146599
transform 1 0 29897 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[37]
timestamp 1698146599
transform 1 0 29561 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[38]
timestamp 1698146599
transform 1 0 29225 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[39]
timestamp 1698146599
transform 1 0 28889 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[40]
timestamp 1698146599
transform 1 0 28553 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[41]
timestamp 1698146599
transform 1 0 28217 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[42]
timestamp 1698146599
transform 1 0 27881 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[43]
timestamp 1698146599
transform 1 0 27545 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[44]
timestamp 1698146599
transform 1 0 27209 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[45]
timestamp 1698146599
transform 1 0 26873 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[46]
timestamp 1698146599
transform 1 0 26537 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[47]
timestamp 1698146599
transform 1 0 26201 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[48]
timestamp 1698146599
transform 1 0 25865 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[49]
timestamp 1698146599
transform 1 0 25529 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[50]
timestamp 1698146599
transform 1 0 25193 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[51]
timestamp 1698146599
transform 1 0 24857 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[52]
timestamp 1698146599
transform 1 0 24521 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[53]
timestamp 1698146599
transform 1 0 24185 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[54]
timestamp 1698146599
transform 1 0 23849 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[55]
timestamp 1698146599
transform 1 0 23513 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[56]
timestamp 1698146599
transform 1 0 23177 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[57]
timestamp 1698146599
transform 1 0 22841 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[58]
timestamp 1698146599
transform 1 0 22505 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[59]
timestamp 1698146599
transform 1 0 22169 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[60]
timestamp 1698146599
transform 1 0 21833 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[61]
timestamp 1698146599
transform 1 0 21497 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[62]
timestamp 1698146599
transform 1 0 21161 0 1 2
box 343 298 679 844
use hgu_cdac_unit  x7[63]
timestamp 1698146599
transform 1 0 20825 0 1 2
box 343 298 679 844
<< end >>
