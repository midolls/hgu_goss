magic
tech sky130A
magscale 1 2
timestamp 1698859995
<< nwell >>
rect 522 3138 6705 3326
rect 7211 3138 13394 3326
rect 522 2675 13394 3138
rect 24 2354 13394 2675
rect 522 2344 13394 2354
rect 522 2146 6705 2344
rect 522 1995 6751 2146
rect 7211 2146 13394 2344
rect 7211 1995 13440 2146
rect 1198 1962 1416 1995
rect 1930 1962 2274 1995
rect 3142 1962 3486 1995
rect 4354 1962 4698 1995
rect 5566 1962 5910 1995
rect 6340 1977 6751 1995
rect 6340 1976 6559 1977
rect 7887 1962 8105 1995
rect 8619 1962 8963 1995
rect 9831 1962 10175 1995
rect 11043 1962 11387 1995
rect 12255 1962 12599 1995
rect 13029 1977 13440 1995
rect 13029 1976 13248 1977
rect 290 -1029 509 -1028
rect 98 -1047 509 -1029
rect 939 -1047 1283 -1014
rect 2151 -1047 2495 -1014
rect 3363 -1047 3707 -1014
rect 4575 -1047 4919 -1014
rect 5433 -1047 5651 -1014
rect 7045 -1029 7264 -1028
rect 6853 -1047 7264 -1029
rect 7694 -1047 8038 -1014
rect 8906 -1047 9250 -1014
rect 10118 -1047 10462 -1014
rect 11330 -1047 11674 -1014
rect 12188 -1047 12406 -1014
rect 98 -1198 6327 -1047
rect 144 -1406 6327 -1198
rect 6853 -1198 13082 -1047
rect 6899 -1406 13082 -1198
rect 144 -1727 6825 -1406
rect 6899 -1727 13580 -1406
rect 144 -2378 6327 -1727
rect 6899 -2378 13082 -1727
<< pwell >>
rect 104 2114 290 2296
rect 294 2114 480 2296
rect 104 2110 125 2114
rect 91 2076 125 2110
rect 459 2110 480 2114
rect 459 2076 493 2110
rect 6793 2114 6979 2296
rect 6983 2114 7169 2296
rect 6793 2110 6814 2114
rect 6780 2076 6814 2110
rect 7148 2110 7169 2114
rect 7148 2076 7182 2110
rect 1337 1002 1507 1172
rect 2069 1002 2239 1172
rect 2673 1002 2843 1172
rect 3281 1002 3451 1172
rect 3885 1002 4055 1172
rect 4619 1002 4789 1172
rect 5223 1002 5393 1172
rect 5955 1002 6125 1172
rect 8026 1002 8196 1172
rect 8758 1002 8928 1172
rect 9362 1002 9532 1172
rect 9970 1002 10140 1172
rect 10574 1002 10744 1172
rect 11308 1002 11478 1172
rect 11912 1002 12082 1172
rect 12644 1002 12814 1172
rect 724 -224 894 -54
rect 1456 -224 1626 -54
rect 2060 -224 2230 -54
rect 2794 -224 2964 -54
rect 3398 -224 3568 -54
rect 4006 -224 4176 -54
rect 4610 -224 4780 -54
rect 5342 -224 5512 -54
rect 7479 -224 7649 -54
rect 8211 -224 8381 -54
rect 8815 -224 8985 -54
rect 9549 -224 9719 -54
rect 10153 -224 10323 -54
rect 10761 -224 10931 -54
rect 11365 -224 11535 -54
rect 12097 -224 12267 -54
rect 6356 -1162 6390 -1128
rect 6369 -1166 6390 -1162
rect 6724 -1162 6758 -1128
rect 6724 -1166 6745 -1162
rect 6369 -1348 6555 -1166
rect 6559 -1348 6745 -1166
rect 13111 -1162 13145 -1128
rect 13124 -1166 13145 -1162
rect 13479 -1162 13513 -1128
rect 13479 -1166 13500 -1162
rect 13124 -1348 13310 -1166
rect 13314 -1348 13500 -1166
<< nmos >>
rect 1647 1810 1677 1894
rect 2379 1810 2409 1894
rect 2503 1810 2533 1894
rect 3591 1810 3621 1894
rect 3715 1810 3745 1894
rect 4929 1810 4959 1894
rect 5053 1810 5083 1894
rect 5785 1810 5815 1894
rect 6435 1811 6465 1895
rect 6527 1811 6557 1895
rect 6623 1811 6653 1895
rect 8336 1810 8366 1894
rect 9068 1810 9098 1894
rect 9192 1810 9222 1894
rect 10280 1810 10310 1894
rect 10404 1810 10434 1894
rect 11618 1810 11648 1894
rect 11742 1810 11772 1894
rect 12474 1810 12504 1894
rect 13124 1811 13154 1895
rect 13216 1811 13246 1895
rect 13312 1811 13342 1895
rect 625 1626 655 1710
rect 697 1626 727 1710
rect 6435 1673 6465 1757
rect 7314 1626 7344 1710
rect 7386 1626 7416 1710
rect 13124 1673 13154 1757
rect 625 1488 655 1572
rect 697 1488 727 1572
rect 7314 1488 7344 1572
rect 7386 1488 7416 1572
rect 625 1350 655 1434
rect 697 1350 727 1434
rect 7314 1350 7344 1434
rect 7386 1350 7416 1434
rect 625 1212 655 1296
rect 697 1212 727 1296
rect 7314 1212 7344 1296
rect 7386 1212 7416 1296
rect 625 1074 655 1158
rect 697 1074 727 1158
rect 7314 1074 7344 1158
rect 7386 1074 7416 1158
rect 625 936 655 1020
rect 697 936 727 1020
rect 7314 936 7344 1020
rect 7386 936 7416 1020
rect 625 798 655 882
rect 697 798 727 882
rect 7314 798 7344 882
rect 7386 798 7416 882
rect 625 660 655 744
rect 697 660 727 744
rect 7314 660 7344 744
rect 7386 660 7416 744
rect 6122 204 6152 288
rect 6194 204 6224 288
rect 12877 204 12907 288
rect 12949 204 12979 288
rect 6122 66 6152 150
rect 6194 66 6224 150
rect 12877 66 12907 150
rect 12949 66 12979 150
rect 6122 -72 6152 12
rect 6194 -72 6224 12
rect 12877 -72 12907 12
rect 12949 -72 12979 12
rect 6122 -210 6152 -126
rect 6194 -210 6224 -126
rect 12877 -210 12907 -126
rect 12949 -210 12979 -126
rect 6122 -348 6152 -264
rect 6194 -348 6224 -264
rect 12877 -348 12907 -264
rect 12949 -348 12979 -264
rect 6122 -486 6152 -402
rect 6194 -486 6224 -402
rect 12877 -486 12907 -402
rect 12949 -486 12979 -402
rect 6122 -624 6152 -540
rect 6194 -624 6224 -540
rect 12877 -624 12907 -540
rect 12949 -624 12979 -540
rect 384 -809 414 -725
rect 6122 -762 6152 -678
rect 6194 -762 6224 -678
rect 7139 -809 7169 -725
rect 12877 -762 12907 -678
rect 12949 -762 12979 -678
rect 196 -947 226 -863
rect 292 -947 322 -863
rect 384 -947 414 -863
rect 1034 -946 1064 -862
rect 1766 -946 1796 -862
rect 1890 -946 1920 -862
rect 3104 -946 3134 -862
rect 3228 -946 3258 -862
rect 4316 -946 4346 -862
rect 4440 -946 4470 -862
rect 5172 -946 5202 -862
rect 6951 -947 6981 -863
rect 7047 -947 7077 -863
rect 7139 -947 7169 -863
rect 7789 -946 7819 -862
rect 8521 -946 8551 -862
rect 8645 -946 8675 -862
rect 9859 -946 9889 -862
rect 9983 -946 10013 -862
rect 11071 -946 11101 -862
rect 11195 -946 11225 -862
rect 11927 -946 11957 -862
<< scnmos >>
rect 182 2140 212 2270
rect 372 2140 402 2270
rect 6871 2140 6901 2270
rect 7061 2140 7091 2270
rect 6447 -1322 6477 -1192
rect 6637 -1322 6667 -1192
rect 13202 -1322 13232 -1192
rect 13392 -1322 13422 -1192
<< pmos >>
rect 1292 2011 1322 2095
rect 2024 2011 2054 2095
rect 2150 2011 2180 2095
rect 3236 2011 3266 2095
rect 3362 2011 3392 2095
rect 4448 2011 4478 2095
rect 4574 2011 4604 2095
rect 5660 2011 5690 2095
rect 5786 2011 5816 2095
rect 7981 2011 8011 2095
rect 8713 2011 8743 2095
rect 8839 2011 8869 2095
rect 9925 2011 9955 2095
rect 10051 2011 10081 2095
rect 11137 2011 11167 2095
rect 11263 2011 11293 2095
rect 12349 2011 12379 2095
rect 12475 2011 12505 2095
rect 1033 -1147 1063 -1063
rect 1159 -1147 1189 -1063
rect 2245 -1147 2275 -1063
rect 2371 -1147 2401 -1063
rect 3457 -1147 3487 -1063
rect 3583 -1147 3613 -1063
rect 4669 -1147 4699 -1063
rect 4795 -1147 4825 -1063
rect 5527 -1147 5557 -1063
rect 7788 -1147 7818 -1063
rect 7914 -1147 7944 -1063
rect 9000 -1147 9030 -1063
rect 9126 -1147 9156 -1063
rect 10212 -1147 10242 -1063
rect 10338 -1147 10368 -1063
rect 11424 -1147 11454 -1063
rect 11550 -1147 11580 -1063
rect 12282 -1147 12312 -1063
<< scpmoshvt >>
rect 182 2390 212 2590
rect 372 2390 402 2590
rect 6871 2390 6901 2590
rect 7061 2390 7091 2590
rect 6447 -1642 6477 -1442
rect 6637 -1642 6667 -1442
rect 13202 -1642 13232 -1442
rect 13392 -1642 13422 -1442
<< pmoshvt >>
rect 671 3153 701 3237
rect 7360 3153 7390 3237
rect 671 3015 701 3099
rect 7360 3015 7390 3099
rect 671 2877 701 2961
rect 7360 2877 7390 2961
rect 671 2739 701 2823
rect 7360 2739 7390 2823
rect 671 2601 701 2685
rect 7360 2601 7390 2685
rect 671 2463 701 2547
rect 7360 2463 7390 2547
rect 6435 2152 6465 2236
rect 13124 2152 13154 2236
rect 6435 2014 6465 2098
rect 6527 2014 6557 2098
rect 6623 2014 6653 2098
rect 13124 2014 13154 2098
rect 13216 2014 13246 2098
rect 13312 2014 13342 2098
rect 196 -1150 226 -1066
rect 292 -1150 322 -1066
rect 384 -1150 414 -1066
rect 6951 -1150 6981 -1066
rect 7047 -1150 7077 -1066
rect 7139 -1150 7169 -1066
rect 384 -1288 414 -1204
rect 7139 -1288 7169 -1204
rect 6148 -1599 6178 -1515
rect 12903 -1599 12933 -1515
rect 6148 -1737 6178 -1653
rect 12903 -1737 12933 -1653
rect 6148 -1875 6178 -1791
rect 12903 -1875 12933 -1791
rect 6148 -2013 6178 -1929
rect 12903 -2013 12933 -1929
rect 6148 -2151 6178 -2067
rect 12903 -2151 12933 -2067
rect 6148 -2289 6178 -2205
rect 12903 -2289 12933 -2205
<< ndiff >>
rect 130 2258 182 2270
rect 130 2224 138 2258
rect 172 2224 182 2258
rect 130 2190 182 2224
rect 130 2156 138 2190
rect 172 2156 182 2190
rect 130 2140 182 2156
rect 212 2258 264 2270
rect 212 2224 222 2258
rect 256 2224 264 2258
rect 212 2190 264 2224
rect 212 2156 222 2190
rect 256 2156 264 2190
rect 212 2140 264 2156
rect 320 2258 372 2270
rect 320 2224 328 2258
rect 362 2224 372 2258
rect 320 2190 372 2224
rect 320 2156 328 2190
rect 362 2156 372 2190
rect 320 2140 372 2156
rect 402 2258 454 2270
rect 402 2224 412 2258
rect 446 2224 454 2258
rect 6819 2258 6871 2270
rect 402 2190 454 2224
rect 402 2156 412 2190
rect 446 2156 454 2190
rect 402 2140 454 2156
rect 6819 2224 6827 2258
rect 6861 2224 6871 2258
rect 6819 2190 6871 2224
rect 6819 2156 6827 2190
rect 6861 2156 6871 2190
rect 6819 2140 6871 2156
rect 6901 2258 6953 2270
rect 6901 2224 6911 2258
rect 6945 2224 6953 2258
rect 6901 2190 6953 2224
rect 6901 2156 6911 2190
rect 6945 2156 6953 2190
rect 6901 2140 6953 2156
rect 7009 2258 7061 2270
rect 7009 2224 7017 2258
rect 7051 2224 7061 2258
rect 7009 2190 7061 2224
rect 7009 2156 7017 2190
rect 7051 2156 7061 2190
rect 7009 2140 7061 2156
rect 7091 2258 7143 2270
rect 7091 2224 7101 2258
rect 7135 2224 7143 2258
rect 7091 2190 7143 2224
rect 7091 2156 7101 2190
rect 7135 2156 7143 2190
rect 7091 2140 7143 2156
rect 1589 1882 1647 1894
rect 1589 1822 1601 1882
rect 1635 1822 1647 1882
rect 1589 1810 1647 1822
rect 1677 1882 1735 1894
rect 1677 1822 1689 1882
rect 1723 1822 1735 1882
rect 1677 1810 1735 1822
rect 2321 1882 2379 1894
rect 2321 1822 2333 1882
rect 2367 1822 2379 1882
rect 2321 1810 2379 1822
rect 2409 1882 2503 1894
rect 2409 1822 2438 1882
rect 2472 1822 2503 1882
rect 2409 1810 2503 1822
rect 2533 1882 2591 1894
rect 2533 1822 2545 1882
rect 2579 1822 2591 1882
rect 2533 1810 2591 1822
rect 3533 1882 3591 1894
rect 3533 1822 3545 1882
rect 3579 1822 3591 1882
rect 3533 1810 3591 1822
rect 3621 1882 3715 1894
rect 3621 1822 3649 1882
rect 3683 1822 3715 1882
rect 3621 1810 3715 1822
rect 3745 1882 3803 1894
rect 3745 1822 3757 1882
rect 3791 1822 3803 1882
rect 3745 1810 3803 1822
rect 4871 1882 4929 1894
rect 4871 1822 4883 1882
rect 4917 1822 4929 1882
rect 4871 1810 4929 1822
rect 4959 1882 5053 1894
rect 4959 1822 4989 1882
rect 5023 1822 5053 1882
rect 4959 1810 5053 1822
rect 5083 1882 5141 1894
rect 5083 1822 5095 1882
rect 5129 1822 5141 1882
rect 5083 1810 5141 1822
rect 5726 1882 5785 1894
rect 5726 1822 5738 1882
rect 5772 1822 5785 1882
rect 5726 1810 5785 1822
rect 5815 1882 5873 1894
rect 5815 1822 5827 1882
rect 5861 1822 5873 1882
rect 5815 1810 5873 1822
rect 6377 1883 6435 1895
rect 6377 1823 6389 1883
rect 6423 1823 6435 1883
rect 6377 1811 6435 1823
rect 6465 1883 6527 1895
rect 6465 1823 6477 1883
rect 6511 1823 6527 1883
rect 6465 1811 6527 1823
rect 6557 1883 6623 1895
rect 6557 1823 6573 1883
rect 6607 1823 6623 1883
rect 6557 1811 6623 1823
rect 6653 1883 6715 1895
rect 6653 1823 6669 1883
rect 6703 1823 6715 1883
rect 6653 1811 6715 1823
rect 8278 1882 8336 1894
rect 8278 1822 8290 1882
rect 8324 1822 8336 1882
rect 8278 1810 8336 1822
rect 8366 1882 8424 1894
rect 8366 1822 8378 1882
rect 8412 1822 8424 1882
rect 8366 1810 8424 1822
rect 9010 1882 9068 1894
rect 9010 1822 9022 1882
rect 9056 1822 9068 1882
rect 9010 1810 9068 1822
rect 9098 1882 9192 1894
rect 9098 1822 9127 1882
rect 9161 1822 9192 1882
rect 9098 1810 9192 1822
rect 9222 1882 9280 1894
rect 9222 1822 9234 1882
rect 9268 1822 9280 1882
rect 9222 1810 9280 1822
rect 10222 1882 10280 1894
rect 10222 1822 10234 1882
rect 10268 1822 10280 1882
rect 10222 1810 10280 1822
rect 10310 1882 10404 1894
rect 10310 1822 10338 1882
rect 10372 1822 10404 1882
rect 10310 1810 10404 1822
rect 10434 1882 10492 1894
rect 10434 1822 10446 1882
rect 10480 1822 10492 1882
rect 10434 1810 10492 1822
rect 11560 1882 11618 1894
rect 11560 1822 11572 1882
rect 11606 1822 11618 1882
rect 11560 1810 11618 1822
rect 11648 1882 11742 1894
rect 11648 1822 11678 1882
rect 11712 1822 11742 1882
rect 11648 1810 11742 1822
rect 11772 1882 11830 1894
rect 11772 1822 11784 1882
rect 11818 1822 11830 1882
rect 11772 1810 11830 1822
rect 12415 1882 12474 1894
rect 12415 1822 12427 1882
rect 12461 1822 12474 1882
rect 12415 1810 12474 1822
rect 12504 1882 12562 1894
rect 12504 1822 12516 1882
rect 12550 1822 12562 1882
rect 12504 1810 12562 1822
rect 13066 1883 13124 1895
rect 13066 1823 13078 1883
rect 13112 1823 13124 1883
rect 13066 1811 13124 1823
rect 13154 1883 13216 1895
rect 13154 1823 13166 1883
rect 13200 1823 13216 1883
rect 13154 1811 13216 1823
rect 13246 1883 13312 1895
rect 13246 1823 13262 1883
rect 13296 1823 13312 1883
rect 13246 1811 13312 1823
rect 13342 1883 13404 1895
rect 13342 1823 13358 1883
rect 13392 1823 13404 1883
rect 13342 1811 13404 1823
rect 6377 1745 6435 1757
rect 567 1698 625 1710
rect 567 1638 579 1698
rect 613 1638 625 1698
rect 567 1626 625 1638
rect 655 1626 697 1710
rect 727 1698 785 1710
rect 727 1638 739 1698
rect 773 1638 785 1698
rect 6377 1685 6389 1745
rect 6423 1685 6435 1745
rect 6377 1673 6435 1685
rect 6465 1745 6523 1757
rect 6465 1685 6477 1745
rect 6511 1685 6523 1745
rect 13066 1745 13124 1757
rect 6465 1673 6523 1685
rect 7256 1698 7314 1710
rect 727 1626 785 1638
rect 7256 1638 7268 1698
rect 7302 1638 7314 1698
rect 7256 1626 7314 1638
rect 7344 1626 7386 1710
rect 7416 1698 7474 1710
rect 7416 1638 7428 1698
rect 7462 1638 7474 1698
rect 13066 1685 13078 1745
rect 13112 1685 13124 1745
rect 13066 1673 13124 1685
rect 13154 1745 13212 1757
rect 13154 1685 13166 1745
rect 13200 1685 13212 1745
rect 13154 1673 13212 1685
rect 7416 1626 7474 1638
rect 567 1560 625 1572
rect 567 1500 579 1560
rect 613 1500 625 1560
rect 567 1488 625 1500
rect 655 1488 697 1572
rect 727 1560 785 1572
rect 727 1500 739 1560
rect 773 1500 785 1560
rect 727 1488 785 1500
rect 7256 1560 7314 1572
rect 7256 1500 7268 1560
rect 7302 1500 7314 1560
rect 7256 1488 7314 1500
rect 7344 1488 7386 1572
rect 7416 1560 7474 1572
rect 7416 1500 7428 1560
rect 7462 1500 7474 1560
rect 7416 1488 7474 1500
rect 567 1422 625 1434
rect 567 1362 579 1422
rect 613 1362 625 1422
rect 567 1350 625 1362
rect 655 1350 697 1434
rect 727 1422 785 1434
rect 727 1362 739 1422
rect 773 1362 785 1422
rect 727 1350 785 1362
rect 7256 1422 7314 1434
rect 7256 1362 7268 1422
rect 7302 1362 7314 1422
rect 7256 1350 7314 1362
rect 7344 1350 7386 1434
rect 7416 1422 7474 1434
rect 7416 1362 7428 1422
rect 7462 1362 7474 1422
rect 7416 1350 7474 1362
rect 567 1284 625 1296
rect 567 1224 579 1284
rect 613 1224 625 1284
rect 567 1212 625 1224
rect 655 1212 697 1296
rect 727 1284 785 1296
rect 727 1224 739 1284
rect 773 1224 785 1284
rect 727 1212 785 1224
rect 7256 1284 7314 1296
rect 7256 1224 7268 1284
rect 7302 1224 7314 1284
rect 7256 1212 7314 1224
rect 7344 1212 7386 1296
rect 7416 1284 7474 1296
rect 7416 1224 7428 1284
rect 7462 1224 7474 1284
rect 7416 1212 7474 1224
rect 567 1146 625 1158
rect 567 1086 579 1146
rect 613 1086 625 1146
rect 567 1074 625 1086
rect 655 1074 697 1158
rect 727 1146 785 1158
rect 727 1086 739 1146
rect 773 1086 785 1146
rect 727 1074 785 1086
rect 7256 1146 7314 1158
rect 7256 1086 7268 1146
rect 7302 1086 7314 1146
rect 7256 1074 7314 1086
rect 7344 1074 7386 1158
rect 7416 1146 7474 1158
rect 7416 1086 7428 1146
rect 7462 1086 7474 1146
rect 7416 1074 7474 1086
rect 567 1008 625 1020
rect 567 948 579 1008
rect 613 948 625 1008
rect 567 936 625 948
rect 655 936 697 1020
rect 727 1008 785 1020
rect 727 948 739 1008
rect 773 948 785 1008
rect 727 936 785 948
rect 7256 1008 7314 1020
rect 7256 948 7268 1008
rect 7302 948 7314 1008
rect 7256 936 7314 948
rect 7344 936 7386 1020
rect 7416 1008 7474 1020
rect 7416 948 7428 1008
rect 7462 948 7474 1008
rect 7416 936 7474 948
rect 567 870 625 882
rect 567 810 579 870
rect 613 810 625 870
rect 567 798 625 810
rect 655 798 697 882
rect 727 870 785 882
rect 727 810 739 870
rect 773 810 785 870
rect 727 798 785 810
rect 7256 870 7314 882
rect 7256 810 7268 870
rect 7302 810 7314 870
rect 7256 798 7314 810
rect 7344 798 7386 882
rect 7416 870 7474 882
rect 7416 810 7428 870
rect 7462 810 7474 870
rect 7416 798 7474 810
rect 567 732 625 744
rect 567 672 579 732
rect 613 672 625 732
rect 567 660 625 672
rect 655 660 697 744
rect 727 732 785 744
rect 727 672 739 732
rect 773 672 785 732
rect 727 660 785 672
rect 7256 732 7314 744
rect 7256 672 7268 732
rect 7302 672 7314 732
rect 7256 660 7314 672
rect 7344 660 7386 744
rect 7416 732 7474 744
rect 7416 672 7428 732
rect 7462 672 7474 732
rect 7416 660 7474 672
rect 6064 276 6122 288
rect 6064 216 6076 276
rect 6110 216 6122 276
rect 6064 204 6122 216
rect 6152 204 6194 288
rect 6224 276 6282 288
rect 6224 216 6236 276
rect 6270 216 6282 276
rect 6224 204 6282 216
rect 12819 276 12877 288
rect 12819 216 12831 276
rect 12865 216 12877 276
rect 12819 204 12877 216
rect 12907 204 12949 288
rect 12979 276 13037 288
rect 12979 216 12991 276
rect 13025 216 13037 276
rect 12979 204 13037 216
rect 6064 138 6122 150
rect 6064 78 6076 138
rect 6110 78 6122 138
rect 6064 66 6122 78
rect 6152 66 6194 150
rect 6224 138 6282 150
rect 6224 78 6236 138
rect 6270 78 6282 138
rect 6224 66 6282 78
rect 12819 138 12877 150
rect 12819 78 12831 138
rect 12865 78 12877 138
rect 12819 66 12877 78
rect 12907 66 12949 150
rect 12979 138 13037 150
rect 12979 78 12991 138
rect 13025 78 13037 138
rect 12979 66 13037 78
rect 6064 0 6122 12
rect 6064 -60 6076 0
rect 6110 -60 6122 0
rect 6064 -72 6122 -60
rect 6152 -72 6194 12
rect 6224 0 6282 12
rect 6224 -60 6236 0
rect 6270 -60 6282 0
rect 6224 -72 6282 -60
rect 12819 0 12877 12
rect 12819 -60 12831 0
rect 12865 -60 12877 0
rect 12819 -72 12877 -60
rect 12907 -72 12949 12
rect 12979 0 13037 12
rect 12979 -60 12991 0
rect 13025 -60 13037 0
rect 12979 -72 13037 -60
rect 6064 -138 6122 -126
rect 6064 -198 6076 -138
rect 6110 -198 6122 -138
rect 6064 -210 6122 -198
rect 6152 -210 6194 -126
rect 6224 -138 6282 -126
rect 6224 -198 6236 -138
rect 6270 -198 6282 -138
rect 6224 -210 6282 -198
rect 12819 -138 12877 -126
rect 12819 -198 12831 -138
rect 12865 -198 12877 -138
rect 12819 -210 12877 -198
rect 12907 -210 12949 -126
rect 12979 -138 13037 -126
rect 12979 -198 12991 -138
rect 13025 -198 13037 -138
rect 12979 -210 13037 -198
rect 6064 -276 6122 -264
rect 6064 -336 6076 -276
rect 6110 -336 6122 -276
rect 6064 -348 6122 -336
rect 6152 -348 6194 -264
rect 6224 -276 6282 -264
rect 6224 -336 6236 -276
rect 6270 -336 6282 -276
rect 6224 -348 6282 -336
rect 12819 -276 12877 -264
rect 12819 -336 12831 -276
rect 12865 -336 12877 -276
rect 12819 -348 12877 -336
rect 12907 -348 12949 -264
rect 12979 -276 13037 -264
rect 12979 -336 12991 -276
rect 13025 -336 13037 -276
rect 12979 -348 13037 -336
rect 6064 -414 6122 -402
rect 6064 -474 6076 -414
rect 6110 -474 6122 -414
rect 6064 -486 6122 -474
rect 6152 -486 6194 -402
rect 6224 -414 6282 -402
rect 6224 -474 6236 -414
rect 6270 -474 6282 -414
rect 6224 -486 6282 -474
rect 12819 -414 12877 -402
rect 12819 -474 12831 -414
rect 12865 -474 12877 -414
rect 12819 -486 12877 -474
rect 12907 -486 12949 -402
rect 12979 -414 13037 -402
rect 12979 -474 12991 -414
rect 13025 -474 13037 -414
rect 12979 -486 13037 -474
rect 6064 -552 6122 -540
rect 6064 -612 6076 -552
rect 6110 -612 6122 -552
rect 6064 -624 6122 -612
rect 6152 -624 6194 -540
rect 6224 -552 6282 -540
rect 6224 -612 6236 -552
rect 6270 -612 6282 -552
rect 6224 -624 6282 -612
rect 12819 -552 12877 -540
rect 12819 -612 12831 -552
rect 12865 -612 12877 -552
rect 12819 -624 12877 -612
rect 12907 -624 12949 -540
rect 12979 -552 13037 -540
rect 12979 -612 12991 -552
rect 13025 -612 13037 -552
rect 12979 -624 13037 -612
rect 6064 -690 6122 -678
rect 326 -737 384 -725
rect 326 -797 338 -737
rect 372 -797 384 -737
rect 326 -809 384 -797
rect 414 -737 472 -725
rect 414 -797 426 -737
rect 460 -797 472 -737
rect 6064 -750 6076 -690
rect 6110 -750 6122 -690
rect 6064 -762 6122 -750
rect 6152 -762 6194 -678
rect 6224 -690 6282 -678
rect 6224 -750 6236 -690
rect 6270 -750 6282 -690
rect 12819 -690 12877 -678
rect 6224 -762 6282 -750
rect 7081 -737 7139 -725
rect 414 -809 472 -797
rect 7081 -797 7093 -737
rect 7127 -797 7139 -737
rect 7081 -809 7139 -797
rect 7169 -737 7227 -725
rect 7169 -797 7181 -737
rect 7215 -797 7227 -737
rect 12819 -750 12831 -690
rect 12865 -750 12877 -690
rect 12819 -762 12877 -750
rect 12907 -762 12949 -678
rect 12979 -690 13037 -678
rect 12979 -750 12991 -690
rect 13025 -750 13037 -690
rect 12979 -762 13037 -750
rect 7169 -809 7227 -797
rect 134 -875 196 -863
rect 134 -935 146 -875
rect 180 -935 196 -875
rect 134 -947 196 -935
rect 226 -875 292 -863
rect 226 -935 242 -875
rect 276 -935 292 -875
rect 226 -947 292 -935
rect 322 -875 384 -863
rect 322 -935 338 -875
rect 372 -935 384 -875
rect 322 -947 384 -935
rect 414 -875 472 -863
rect 414 -935 426 -875
rect 460 -935 472 -875
rect 414 -947 472 -935
rect 976 -874 1034 -862
rect 976 -934 988 -874
rect 1022 -934 1034 -874
rect 976 -946 1034 -934
rect 1064 -874 1123 -862
rect 1064 -934 1077 -874
rect 1111 -934 1123 -874
rect 1064 -946 1123 -934
rect 1708 -874 1766 -862
rect 1708 -934 1720 -874
rect 1754 -934 1766 -874
rect 1708 -946 1766 -934
rect 1796 -874 1890 -862
rect 1796 -934 1826 -874
rect 1860 -934 1890 -874
rect 1796 -946 1890 -934
rect 1920 -874 1978 -862
rect 1920 -934 1932 -874
rect 1966 -934 1978 -874
rect 1920 -946 1978 -934
rect 3046 -874 3104 -862
rect 3046 -934 3058 -874
rect 3092 -934 3104 -874
rect 3046 -946 3104 -934
rect 3134 -874 3228 -862
rect 3134 -934 3166 -874
rect 3200 -934 3228 -874
rect 3134 -946 3228 -934
rect 3258 -874 3316 -862
rect 3258 -934 3270 -874
rect 3304 -934 3316 -874
rect 3258 -946 3316 -934
rect 4258 -874 4316 -862
rect 4258 -934 4270 -874
rect 4304 -934 4316 -874
rect 4258 -946 4316 -934
rect 4346 -874 4440 -862
rect 4346 -934 4377 -874
rect 4411 -934 4440 -874
rect 4346 -946 4440 -934
rect 4470 -874 4528 -862
rect 4470 -934 4482 -874
rect 4516 -934 4528 -874
rect 4470 -946 4528 -934
rect 5114 -874 5172 -862
rect 5114 -934 5126 -874
rect 5160 -934 5172 -874
rect 5114 -946 5172 -934
rect 5202 -874 5260 -862
rect 5202 -934 5214 -874
rect 5248 -934 5260 -874
rect 5202 -946 5260 -934
rect 6889 -875 6951 -863
rect 6889 -935 6901 -875
rect 6935 -935 6951 -875
rect 6889 -947 6951 -935
rect 6981 -875 7047 -863
rect 6981 -935 6997 -875
rect 7031 -935 7047 -875
rect 6981 -947 7047 -935
rect 7077 -875 7139 -863
rect 7077 -935 7093 -875
rect 7127 -935 7139 -875
rect 7077 -947 7139 -935
rect 7169 -875 7227 -863
rect 7169 -935 7181 -875
rect 7215 -935 7227 -875
rect 7169 -947 7227 -935
rect 7731 -874 7789 -862
rect 7731 -934 7743 -874
rect 7777 -934 7789 -874
rect 7731 -946 7789 -934
rect 7819 -874 7878 -862
rect 7819 -934 7832 -874
rect 7866 -934 7878 -874
rect 7819 -946 7878 -934
rect 8463 -874 8521 -862
rect 8463 -934 8475 -874
rect 8509 -934 8521 -874
rect 8463 -946 8521 -934
rect 8551 -874 8645 -862
rect 8551 -934 8581 -874
rect 8615 -934 8645 -874
rect 8551 -946 8645 -934
rect 8675 -874 8733 -862
rect 8675 -934 8687 -874
rect 8721 -934 8733 -874
rect 8675 -946 8733 -934
rect 9801 -874 9859 -862
rect 9801 -934 9813 -874
rect 9847 -934 9859 -874
rect 9801 -946 9859 -934
rect 9889 -874 9983 -862
rect 9889 -934 9921 -874
rect 9955 -934 9983 -874
rect 9889 -946 9983 -934
rect 10013 -874 10071 -862
rect 10013 -934 10025 -874
rect 10059 -934 10071 -874
rect 10013 -946 10071 -934
rect 11013 -874 11071 -862
rect 11013 -934 11025 -874
rect 11059 -934 11071 -874
rect 11013 -946 11071 -934
rect 11101 -874 11195 -862
rect 11101 -934 11132 -874
rect 11166 -934 11195 -874
rect 11101 -946 11195 -934
rect 11225 -874 11283 -862
rect 11225 -934 11237 -874
rect 11271 -934 11283 -874
rect 11225 -946 11283 -934
rect 11869 -874 11927 -862
rect 11869 -934 11881 -874
rect 11915 -934 11927 -874
rect 11869 -946 11927 -934
rect 11957 -874 12015 -862
rect 11957 -934 11969 -874
rect 12003 -934 12015 -874
rect 11957 -946 12015 -934
rect 6395 -1208 6447 -1192
rect 6395 -1242 6403 -1208
rect 6437 -1242 6447 -1208
rect 6395 -1276 6447 -1242
rect 6395 -1310 6403 -1276
rect 6437 -1310 6447 -1276
rect 6395 -1322 6447 -1310
rect 6477 -1208 6529 -1192
rect 6477 -1242 6487 -1208
rect 6521 -1242 6529 -1208
rect 6477 -1276 6529 -1242
rect 6477 -1310 6487 -1276
rect 6521 -1310 6529 -1276
rect 6477 -1322 6529 -1310
rect 6585 -1208 6637 -1192
rect 6585 -1242 6593 -1208
rect 6627 -1242 6637 -1208
rect 6585 -1276 6637 -1242
rect 6585 -1310 6593 -1276
rect 6627 -1310 6637 -1276
rect 6585 -1322 6637 -1310
rect 6667 -1208 6719 -1192
rect 6667 -1242 6677 -1208
rect 6711 -1242 6719 -1208
rect 6667 -1276 6719 -1242
rect 6667 -1310 6677 -1276
rect 6711 -1310 6719 -1276
rect 13150 -1208 13202 -1192
rect 13150 -1242 13158 -1208
rect 13192 -1242 13202 -1208
rect 13150 -1276 13202 -1242
rect 6667 -1322 6719 -1310
rect 13150 -1310 13158 -1276
rect 13192 -1310 13202 -1276
rect 13150 -1322 13202 -1310
rect 13232 -1208 13284 -1192
rect 13232 -1242 13242 -1208
rect 13276 -1242 13284 -1208
rect 13232 -1276 13284 -1242
rect 13232 -1310 13242 -1276
rect 13276 -1310 13284 -1276
rect 13232 -1322 13284 -1310
rect 13340 -1208 13392 -1192
rect 13340 -1242 13348 -1208
rect 13382 -1242 13392 -1208
rect 13340 -1276 13392 -1242
rect 13340 -1310 13348 -1276
rect 13382 -1310 13392 -1276
rect 13340 -1322 13392 -1310
rect 13422 -1208 13474 -1192
rect 13422 -1242 13432 -1208
rect 13466 -1242 13474 -1208
rect 13422 -1276 13474 -1242
rect 13422 -1310 13432 -1276
rect 13466 -1310 13474 -1276
rect 13422 -1322 13474 -1310
<< pdiff >>
rect 613 3225 671 3237
rect 613 3165 625 3225
rect 659 3165 671 3225
rect 613 3153 671 3165
rect 701 3225 759 3237
rect 701 3165 713 3225
rect 747 3165 759 3225
rect 701 3153 759 3165
rect 7302 3225 7360 3237
rect 7302 3165 7314 3225
rect 7348 3165 7360 3225
rect 7302 3153 7360 3165
rect 7390 3225 7448 3237
rect 7390 3165 7402 3225
rect 7436 3165 7448 3225
rect 7390 3153 7448 3165
rect 613 3087 671 3099
rect 613 3027 625 3087
rect 659 3027 671 3087
rect 613 3015 671 3027
rect 701 3087 759 3099
rect 701 3027 713 3087
rect 747 3027 759 3087
rect 701 3015 759 3027
rect 7302 3087 7360 3099
rect 7302 3027 7314 3087
rect 7348 3027 7360 3087
rect 7302 3015 7360 3027
rect 7390 3087 7448 3099
rect 7390 3027 7402 3087
rect 7436 3027 7448 3087
rect 7390 3015 7448 3027
rect 613 2949 671 2961
rect 613 2889 625 2949
rect 659 2889 671 2949
rect 613 2877 671 2889
rect 701 2949 759 2961
rect 701 2889 713 2949
rect 747 2889 759 2949
rect 701 2877 759 2889
rect 7302 2949 7360 2961
rect 7302 2889 7314 2949
rect 7348 2889 7360 2949
rect 7302 2877 7360 2889
rect 7390 2949 7448 2961
rect 7390 2889 7402 2949
rect 7436 2889 7448 2949
rect 7390 2877 7448 2889
rect 613 2811 671 2823
rect 613 2751 625 2811
rect 659 2751 671 2811
rect 613 2739 671 2751
rect 701 2811 759 2823
rect 701 2751 713 2811
rect 747 2751 759 2811
rect 701 2739 759 2751
rect 7302 2811 7360 2823
rect 7302 2751 7314 2811
rect 7348 2751 7360 2811
rect 7302 2739 7360 2751
rect 7390 2811 7448 2823
rect 7390 2751 7402 2811
rect 7436 2751 7448 2811
rect 7390 2739 7448 2751
rect 613 2673 671 2685
rect 613 2613 625 2673
rect 659 2613 671 2673
rect 613 2601 671 2613
rect 701 2673 759 2685
rect 701 2613 713 2673
rect 747 2613 759 2673
rect 7302 2673 7360 2685
rect 701 2601 759 2613
rect 130 2578 182 2590
rect 130 2544 138 2578
rect 172 2544 182 2578
rect 130 2510 182 2544
rect 130 2476 138 2510
rect 172 2476 182 2510
rect 130 2442 182 2476
rect 130 2408 138 2442
rect 172 2408 182 2442
rect 130 2390 182 2408
rect 212 2578 264 2590
rect 212 2544 222 2578
rect 256 2544 264 2578
rect 212 2510 264 2544
rect 212 2476 222 2510
rect 256 2476 264 2510
rect 212 2442 264 2476
rect 212 2408 222 2442
rect 256 2408 264 2442
rect 212 2390 264 2408
rect 320 2578 372 2590
rect 320 2544 328 2578
rect 362 2544 372 2578
rect 320 2510 372 2544
rect 320 2476 328 2510
rect 362 2476 372 2510
rect 320 2442 372 2476
rect 320 2408 328 2442
rect 362 2408 372 2442
rect 320 2390 372 2408
rect 402 2578 454 2590
rect 402 2544 412 2578
rect 446 2544 454 2578
rect 7302 2613 7314 2673
rect 7348 2613 7360 2673
rect 7302 2601 7360 2613
rect 7390 2673 7448 2685
rect 7390 2613 7402 2673
rect 7436 2613 7448 2673
rect 7390 2601 7448 2613
rect 6819 2578 6871 2590
rect 402 2510 454 2544
rect 402 2476 412 2510
rect 446 2476 454 2510
rect 402 2442 454 2476
rect 613 2535 671 2547
rect 613 2475 625 2535
rect 659 2475 671 2535
rect 613 2463 671 2475
rect 701 2535 759 2547
rect 701 2475 713 2535
rect 747 2475 759 2535
rect 701 2463 759 2475
rect 6819 2544 6827 2578
rect 6861 2544 6871 2578
rect 6819 2510 6871 2544
rect 6819 2476 6827 2510
rect 6861 2476 6871 2510
rect 402 2408 412 2442
rect 446 2408 454 2442
rect 6819 2442 6871 2476
rect 402 2390 454 2408
rect 6819 2408 6827 2442
rect 6861 2408 6871 2442
rect 6819 2390 6871 2408
rect 6901 2578 6953 2590
rect 6901 2544 6911 2578
rect 6945 2544 6953 2578
rect 6901 2510 6953 2544
rect 6901 2476 6911 2510
rect 6945 2476 6953 2510
rect 6901 2442 6953 2476
rect 6901 2408 6911 2442
rect 6945 2408 6953 2442
rect 6901 2390 6953 2408
rect 7009 2578 7061 2590
rect 7009 2544 7017 2578
rect 7051 2544 7061 2578
rect 7009 2510 7061 2544
rect 7009 2476 7017 2510
rect 7051 2476 7061 2510
rect 7009 2442 7061 2476
rect 7009 2408 7017 2442
rect 7051 2408 7061 2442
rect 7009 2390 7061 2408
rect 7091 2578 7143 2590
rect 7091 2544 7101 2578
rect 7135 2544 7143 2578
rect 7091 2510 7143 2544
rect 7091 2476 7101 2510
rect 7135 2476 7143 2510
rect 7091 2442 7143 2476
rect 7302 2535 7360 2547
rect 7302 2475 7314 2535
rect 7348 2475 7360 2535
rect 7302 2463 7360 2475
rect 7390 2535 7448 2547
rect 7390 2475 7402 2535
rect 7436 2475 7448 2535
rect 7390 2463 7448 2475
rect 7091 2408 7101 2442
rect 7135 2408 7143 2442
rect 7091 2390 7143 2408
rect 6377 2224 6435 2236
rect 6377 2164 6389 2224
rect 6423 2164 6435 2224
rect 6377 2152 6435 2164
rect 6465 2224 6523 2236
rect 6465 2164 6477 2224
rect 6511 2164 6523 2224
rect 6465 2152 6523 2164
rect 13066 2224 13124 2236
rect 13066 2164 13078 2224
rect 13112 2164 13124 2224
rect 13066 2152 13124 2164
rect 13154 2224 13212 2236
rect 13154 2164 13166 2224
rect 13200 2164 13212 2224
rect 13154 2152 13212 2164
rect 1234 2083 1292 2095
rect 1234 2023 1246 2083
rect 1280 2023 1292 2083
rect 1234 2011 1292 2023
rect 1322 2083 1380 2095
rect 1322 2023 1334 2083
rect 1368 2023 1380 2083
rect 1322 2011 1380 2023
rect 1966 2083 2024 2095
rect 1966 2023 1978 2083
rect 2012 2023 2024 2083
rect 1966 2011 2024 2023
rect 2054 2083 2150 2095
rect 2054 2023 2083 2083
rect 2117 2023 2150 2083
rect 2054 2011 2150 2023
rect 2180 2083 2238 2095
rect 2180 2023 2192 2083
rect 2226 2023 2238 2083
rect 2180 2011 2238 2023
rect 3178 2083 3236 2095
rect 3178 2023 3190 2083
rect 3224 2023 3236 2083
rect 3178 2011 3236 2023
rect 3266 2083 3362 2095
rect 3266 2023 3294 2083
rect 3328 2023 3362 2083
rect 3266 2011 3362 2023
rect 3392 2083 3450 2095
rect 3392 2023 3404 2083
rect 3438 2023 3450 2083
rect 3392 2011 3450 2023
rect 4390 2083 4448 2095
rect 4390 2023 4402 2083
rect 4436 2023 4448 2083
rect 4390 2011 4448 2023
rect 4478 2083 4574 2095
rect 4478 2023 4507 2083
rect 4541 2023 4574 2083
rect 4478 2011 4574 2023
rect 4604 2083 4662 2095
rect 4604 2023 4616 2083
rect 4650 2023 4662 2083
rect 4604 2011 4662 2023
rect 5602 2083 5660 2095
rect 5602 2023 5614 2083
rect 5648 2023 5660 2083
rect 5602 2011 5660 2023
rect 5690 2083 5786 2095
rect 5690 2023 5721 2083
rect 5755 2023 5786 2083
rect 5690 2011 5786 2023
rect 5816 2083 5874 2095
rect 5816 2023 5828 2083
rect 5862 2023 5874 2083
rect 5816 2011 5874 2023
rect 6377 2086 6435 2098
rect 6377 2026 6389 2086
rect 6423 2026 6435 2086
rect 6377 2014 6435 2026
rect 6465 2086 6527 2098
rect 6465 2026 6477 2086
rect 6511 2026 6527 2086
rect 6465 2014 6527 2026
rect 6557 2086 6623 2098
rect 6557 2026 6573 2086
rect 6607 2026 6623 2086
rect 6557 2014 6623 2026
rect 6653 2086 6715 2098
rect 6653 2026 6669 2086
rect 6703 2026 6715 2086
rect 6653 2014 6715 2026
rect 7923 2083 7981 2095
rect 7923 2023 7935 2083
rect 7969 2023 7981 2083
rect 7923 2011 7981 2023
rect 8011 2083 8069 2095
rect 8011 2023 8023 2083
rect 8057 2023 8069 2083
rect 8011 2011 8069 2023
rect 8655 2083 8713 2095
rect 8655 2023 8667 2083
rect 8701 2023 8713 2083
rect 8655 2011 8713 2023
rect 8743 2083 8839 2095
rect 8743 2023 8772 2083
rect 8806 2023 8839 2083
rect 8743 2011 8839 2023
rect 8869 2083 8927 2095
rect 8869 2023 8881 2083
rect 8915 2023 8927 2083
rect 8869 2011 8927 2023
rect 9867 2083 9925 2095
rect 9867 2023 9879 2083
rect 9913 2023 9925 2083
rect 9867 2011 9925 2023
rect 9955 2083 10051 2095
rect 9955 2023 9983 2083
rect 10017 2023 10051 2083
rect 9955 2011 10051 2023
rect 10081 2083 10139 2095
rect 10081 2023 10093 2083
rect 10127 2023 10139 2083
rect 10081 2011 10139 2023
rect 11079 2083 11137 2095
rect 11079 2023 11091 2083
rect 11125 2023 11137 2083
rect 11079 2011 11137 2023
rect 11167 2083 11263 2095
rect 11167 2023 11196 2083
rect 11230 2023 11263 2083
rect 11167 2011 11263 2023
rect 11293 2083 11351 2095
rect 11293 2023 11305 2083
rect 11339 2023 11351 2083
rect 11293 2011 11351 2023
rect 12291 2083 12349 2095
rect 12291 2023 12303 2083
rect 12337 2023 12349 2083
rect 12291 2011 12349 2023
rect 12379 2083 12475 2095
rect 12379 2023 12410 2083
rect 12444 2023 12475 2083
rect 12379 2011 12475 2023
rect 12505 2083 12563 2095
rect 12505 2023 12517 2083
rect 12551 2023 12563 2083
rect 12505 2011 12563 2023
rect 13066 2086 13124 2098
rect 13066 2026 13078 2086
rect 13112 2026 13124 2086
rect 13066 2014 13124 2026
rect 13154 2086 13216 2098
rect 13154 2026 13166 2086
rect 13200 2026 13216 2086
rect 13154 2014 13216 2026
rect 13246 2086 13312 2098
rect 13246 2026 13262 2086
rect 13296 2026 13312 2086
rect 13246 2014 13312 2026
rect 13342 2086 13404 2098
rect 13342 2026 13358 2086
rect 13392 2026 13404 2086
rect 13342 2014 13404 2026
rect 134 -1078 196 -1066
rect 134 -1138 146 -1078
rect 180 -1138 196 -1078
rect 134 -1150 196 -1138
rect 226 -1078 292 -1066
rect 226 -1138 242 -1078
rect 276 -1138 292 -1078
rect 226 -1150 292 -1138
rect 322 -1078 384 -1066
rect 322 -1138 338 -1078
rect 372 -1138 384 -1078
rect 322 -1150 384 -1138
rect 414 -1078 472 -1066
rect 414 -1138 426 -1078
rect 460 -1138 472 -1078
rect 414 -1150 472 -1138
rect 975 -1075 1033 -1063
rect 975 -1135 987 -1075
rect 1021 -1135 1033 -1075
rect 975 -1147 1033 -1135
rect 1063 -1075 1159 -1063
rect 1063 -1135 1094 -1075
rect 1128 -1135 1159 -1075
rect 1063 -1147 1159 -1135
rect 1189 -1075 1247 -1063
rect 1189 -1135 1201 -1075
rect 1235 -1135 1247 -1075
rect 1189 -1147 1247 -1135
rect 2187 -1075 2245 -1063
rect 2187 -1135 2199 -1075
rect 2233 -1135 2245 -1075
rect 2187 -1147 2245 -1135
rect 2275 -1075 2371 -1063
rect 2275 -1135 2308 -1075
rect 2342 -1135 2371 -1075
rect 2275 -1147 2371 -1135
rect 2401 -1075 2459 -1063
rect 2401 -1135 2413 -1075
rect 2447 -1135 2459 -1075
rect 2401 -1147 2459 -1135
rect 3399 -1075 3457 -1063
rect 3399 -1135 3411 -1075
rect 3445 -1135 3457 -1075
rect 3399 -1147 3457 -1135
rect 3487 -1075 3583 -1063
rect 3487 -1135 3521 -1075
rect 3555 -1135 3583 -1075
rect 3487 -1147 3583 -1135
rect 3613 -1075 3671 -1063
rect 3613 -1135 3625 -1075
rect 3659 -1135 3671 -1075
rect 3613 -1147 3671 -1135
rect 4611 -1075 4669 -1063
rect 4611 -1135 4623 -1075
rect 4657 -1135 4669 -1075
rect 4611 -1147 4669 -1135
rect 4699 -1075 4795 -1063
rect 4699 -1135 4732 -1075
rect 4766 -1135 4795 -1075
rect 4699 -1147 4795 -1135
rect 4825 -1075 4883 -1063
rect 4825 -1135 4837 -1075
rect 4871 -1135 4883 -1075
rect 4825 -1147 4883 -1135
rect 5469 -1075 5527 -1063
rect 5469 -1135 5481 -1075
rect 5515 -1135 5527 -1075
rect 5469 -1147 5527 -1135
rect 5557 -1075 5615 -1063
rect 5557 -1135 5569 -1075
rect 5603 -1135 5615 -1075
rect 5557 -1147 5615 -1135
rect 6889 -1078 6951 -1066
rect 6889 -1138 6901 -1078
rect 6935 -1138 6951 -1078
rect 6889 -1150 6951 -1138
rect 6981 -1078 7047 -1066
rect 6981 -1138 6997 -1078
rect 7031 -1138 7047 -1078
rect 6981 -1150 7047 -1138
rect 7077 -1078 7139 -1066
rect 7077 -1138 7093 -1078
rect 7127 -1138 7139 -1078
rect 7077 -1150 7139 -1138
rect 7169 -1078 7227 -1066
rect 7169 -1138 7181 -1078
rect 7215 -1138 7227 -1078
rect 7169 -1150 7227 -1138
rect 7730 -1075 7788 -1063
rect 7730 -1135 7742 -1075
rect 7776 -1135 7788 -1075
rect 7730 -1147 7788 -1135
rect 7818 -1075 7914 -1063
rect 7818 -1135 7849 -1075
rect 7883 -1135 7914 -1075
rect 7818 -1147 7914 -1135
rect 7944 -1075 8002 -1063
rect 7944 -1135 7956 -1075
rect 7990 -1135 8002 -1075
rect 7944 -1147 8002 -1135
rect 8942 -1075 9000 -1063
rect 8942 -1135 8954 -1075
rect 8988 -1135 9000 -1075
rect 8942 -1147 9000 -1135
rect 9030 -1075 9126 -1063
rect 9030 -1135 9063 -1075
rect 9097 -1135 9126 -1075
rect 9030 -1147 9126 -1135
rect 9156 -1075 9214 -1063
rect 9156 -1135 9168 -1075
rect 9202 -1135 9214 -1075
rect 9156 -1147 9214 -1135
rect 10154 -1075 10212 -1063
rect 10154 -1135 10166 -1075
rect 10200 -1135 10212 -1075
rect 10154 -1147 10212 -1135
rect 10242 -1075 10338 -1063
rect 10242 -1135 10276 -1075
rect 10310 -1135 10338 -1075
rect 10242 -1147 10338 -1135
rect 10368 -1075 10426 -1063
rect 10368 -1135 10380 -1075
rect 10414 -1135 10426 -1075
rect 10368 -1147 10426 -1135
rect 11366 -1075 11424 -1063
rect 11366 -1135 11378 -1075
rect 11412 -1135 11424 -1075
rect 11366 -1147 11424 -1135
rect 11454 -1075 11550 -1063
rect 11454 -1135 11487 -1075
rect 11521 -1135 11550 -1075
rect 11454 -1147 11550 -1135
rect 11580 -1075 11638 -1063
rect 11580 -1135 11592 -1075
rect 11626 -1135 11638 -1075
rect 11580 -1147 11638 -1135
rect 12224 -1075 12282 -1063
rect 12224 -1135 12236 -1075
rect 12270 -1135 12282 -1075
rect 12224 -1147 12282 -1135
rect 12312 -1075 12370 -1063
rect 12312 -1135 12324 -1075
rect 12358 -1135 12370 -1075
rect 12312 -1147 12370 -1135
rect 326 -1216 384 -1204
rect 326 -1276 338 -1216
rect 372 -1276 384 -1216
rect 326 -1288 384 -1276
rect 414 -1216 472 -1204
rect 414 -1276 426 -1216
rect 460 -1276 472 -1216
rect 414 -1288 472 -1276
rect 7081 -1216 7139 -1204
rect 7081 -1276 7093 -1216
rect 7127 -1276 7139 -1216
rect 7081 -1288 7139 -1276
rect 7169 -1216 7227 -1204
rect 7169 -1276 7181 -1216
rect 7215 -1276 7227 -1216
rect 7169 -1288 7227 -1276
rect 6395 -1460 6447 -1442
rect 6395 -1494 6403 -1460
rect 6437 -1494 6447 -1460
rect 6090 -1527 6148 -1515
rect 6090 -1587 6102 -1527
rect 6136 -1587 6148 -1527
rect 6090 -1599 6148 -1587
rect 6178 -1527 6236 -1515
rect 6178 -1587 6190 -1527
rect 6224 -1587 6236 -1527
rect 6178 -1599 6236 -1587
rect 6395 -1528 6447 -1494
rect 6395 -1562 6403 -1528
rect 6437 -1562 6447 -1528
rect 6395 -1596 6447 -1562
rect 6395 -1630 6403 -1596
rect 6437 -1630 6447 -1596
rect 6395 -1642 6447 -1630
rect 6477 -1460 6529 -1442
rect 6477 -1494 6487 -1460
rect 6521 -1494 6529 -1460
rect 6477 -1528 6529 -1494
rect 6477 -1562 6487 -1528
rect 6521 -1562 6529 -1528
rect 6477 -1596 6529 -1562
rect 6477 -1630 6487 -1596
rect 6521 -1630 6529 -1596
rect 6477 -1642 6529 -1630
rect 6585 -1460 6637 -1442
rect 6585 -1494 6593 -1460
rect 6627 -1494 6637 -1460
rect 6585 -1528 6637 -1494
rect 6585 -1562 6593 -1528
rect 6627 -1562 6637 -1528
rect 6585 -1596 6637 -1562
rect 6585 -1630 6593 -1596
rect 6627 -1630 6637 -1596
rect 6585 -1642 6637 -1630
rect 6667 -1460 6719 -1442
rect 6667 -1494 6677 -1460
rect 6711 -1494 6719 -1460
rect 13150 -1460 13202 -1442
rect 6667 -1528 6719 -1494
rect 13150 -1494 13158 -1460
rect 13192 -1494 13202 -1460
rect 6667 -1562 6677 -1528
rect 6711 -1562 6719 -1528
rect 6667 -1596 6719 -1562
rect 6667 -1630 6677 -1596
rect 6711 -1630 6719 -1596
rect 12845 -1527 12903 -1515
rect 12845 -1587 12857 -1527
rect 12891 -1587 12903 -1527
rect 12845 -1599 12903 -1587
rect 12933 -1527 12991 -1515
rect 12933 -1587 12945 -1527
rect 12979 -1587 12991 -1527
rect 12933 -1599 12991 -1587
rect 13150 -1528 13202 -1494
rect 13150 -1562 13158 -1528
rect 13192 -1562 13202 -1528
rect 13150 -1596 13202 -1562
rect 6667 -1642 6719 -1630
rect 6090 -1665 6148 -1653
rect 6090 -1725 6102 -1665
rect 6136 -1725 6148 -1665
rect 6090 -1737 6148 -1725
rect 6178 -1665 6236 -1653
rect 6178 -1725 6190 -1665
rect 6224 -1725 6236 -1665
rect 13150 -1630 13158 -1596
rect 13192 -1630 13202 -1596
rect 13150 -1642 13202 -1630
rect 13232 -1460 13284 -1442
rect 13232 -1494 13242 -1460
rect 13276 -1494 13284 -1460
rect 13232 -1528 13284 -1494
rect 13232 -1562 13242 -1528
rect 13276 -1562 13284 -1528
rect 13232 -1596 13284 -1562
rect 13232 -1630 13242 -1596
rect 13276 -1630 13284 -1596
rect 13232 -1642 13284 -1630
rect 13340 -1460 13392 -1442
rect 13340 -1494 13348 -1460
rect 13382 -1494 13392 -1460
rect 13340 -1528 13392 -1494
rect 13340 -1562 13348 -1528
rect 13382 -1562 13392 -1528
rect 13340 -1596 13392 -1562
rect 13340 -1630 13348 -1596
rect 13382 -1630 13392 -1596
rect 13340 -1642 13392 -1630
rect 13422 -1460 13474 -1442
rect 13422 -1494 13432 -1460
rect 13466 -1494 13474 -1460
rect 13422 -1528 13474 -1494
rect 13422 -1562 13432 -1528
rect 13466 -1562 13474 -1528
rect 13422 -1596 13474 -1562
rect 13422 -1630 13432 -1596
rect 13466 -1630 13474 -1596
rect 13422 -1642 13474 -1630
rect 12845 -1665 12903 -1653
rect 6178 -1737 6236 -1725
rect 12845 -1725 12857 -1665
rect 12891 -1725 12903 -1665
rect 12845 -1737 12903 -1725
rect 12933 -1665 12991 -1653
rect 12933 -1725 12945 -1665
rect 12979 -1725 12991 -1665
rect 12933 -1737 12991 -1725
rect 6090 -1803 6148 -1791
rect 6090 -1863 6102 -1803
rect 6136 -1863 6148 -1803
rect 6090 -1875 6148 -1863
rect 6178 -1803 6236 -1791
rect 6178 -1863 6190 -1803
rect 6224 -1863 6236 -1803
rect 6178 -1875 6236 -1863
rect 12845 -1803 12903 -1791
rect 12845 -1863 12857 -1803
rect 12891 -1863 12903 -1803
rect 12845 -1875 12903 -1863
rect 12933 -1803 12991 -1791
rect 12933 -1863 12945 -1803
rect 12979 -1863 12991 -1803
rect 12933 -1875 12991 -1863
rect 6090 -1941 6148 -1929
rect 6090 -2001 6102 -1941
rect 6136 -2001 6148 -1941
rect 6090 -2013 6148 -2001
rect 6178 -1941 6236 -1929
rect 6178 -2001 6190 -1941
rect 6224 -2001 6236 -1941
rect 6178 -2013 6236 -2001
rect 12845 -1941 12903 -1929
rect 12845 -2001 12857 -1941
rect 12891 -2001 12903 -1941
rect 12845 -2013 12903 -2001
rect 12933 -1941 12991 -1929
rect 12933 -2001 12945 -1941
rect 12979 -2001 12991 -1941
rect 12933 -2013 12991 -2001
rect 6090 -2079 6148 -2067
rect 6090 -2139 6102 -2079
rect 6136 -2139 6148 -2079
rect 6090 -2151 6148 -2139
rect 6178 -2079 6236 -2067
rect 6178 -2139 6190 -2079
rect 6224 -2139 6236 -2079
rect 6178 -2151 6236 -2139
rect 12845 -2079 12903 -2067
rect 12845 -2139 12857 -2079
rect 12891 -2139 12903 -2079
rect 12845 -2151 12903 -2139
rect 12933 -2079 12991 -2067
rect 12933 -2139 12945 -2079
rect 12979 -2139 12991 -2079
rect 12933 -2151 12991 -2139
rect 6090 -2217 6148 -2205
rect 6090 -2277 6102 -2217
rect 6136 -2277 6148 -2217
rect 6090 -2289 6148 -2277
rect 6178 -2217 6236 -2205
rect 6178 -2277 6190 -2217
rect 6224 -2277 6236 -2217
rect 6178 -2289 6236 -2277
rect 12845 -2217 12903 -2205
rect 12845 -2277 12857 -2217
rect 12891 -2277 12903 -2217
rect 12845 -2289 12903 -2277
rect 12933 -2217 12991 -2205
rect 12933 -2277 12945 -2217
rect 12979 -2277 12991 -2217
rect 12933 -2289 12991 -2277
<< ndiffc >>
rect 138 2224 172 2258
rect 138 2156 172 2190
rect 222 2224 256 2258
rect 222 2156 256 2190
rect 328 2224 362 2258
rect 328 2156 362 2190
rect 412 2224 446 2258
rect 412 2156 446 2190
rect 6827 2224 6861 2258
rect 6827 2156 6861 2190
rect 6911 2224 6945 2258
rect 6911 2156 6945 2190
rect 7017 2224 7051 2258
rect 7017 2156 7051 2190
rect 7101 2224 7135 2258
rect 7101 2156 7135 2190
rect 1601 1822 1635 1882
rect 1689 1822 1723 1882
rect 2333 1822 2367 1882
rect 2438 1822 2472 1882
rect 2545 1822 2579 1882
rect 3545 1822 3579 1882
rect 3649 1822 3683 1882
rect 3757 1822 3791 1882
rect 4883 1822 4917 1882
rect 4989 1822 5023 1882
rect 5095 1822 5129 1882
rect 5738 1822 5772 1882
rect 5827 1822 5861 1882
rect 6389 1823 6423 1883
rect 6477 1823 6511 1883
rect 6573 1823 6607 1883
rect 6669 1823 6703 1883
rect 8290 1822 8324 1882
rect 8378 1822 8412 1882
rect 9022 1822 9056 1882
rect 9127 1822 9161 1882
rect 9234 1822 9268 1882
rect 10234 1822 10268 1882
rect 10338 1822 10372 1882
rect 10446 1822 10480 1882
rect 11572 1822 11606 1882
rect 11678 1822 11712 1882
rect 11784 1822 11818 1882
rect 12427 1822 12461 1882
rect 12516 1822 12550 1882
rect 13078 1823 13112 1883
rect 13166 1823 13200 1883
rect 13262 1823 13296 1883
rect 13358 1823 13392 1883
rect 579 1638 613 1698
rect 739 1638 773 1698
rect 6389 1685 6423 1745
rect 6477 1685 6511 1745
rect 7268 1638 7302 1698
rect 7428 1638 7462 1698
rect 13078 1685 13112 1745
rect 13166 1685 13200 1745
rect 579 1500 613 1560
rect 739 1500 773 1560
rect 7268 1500 7302 1560
rect 7428 1500 7462 1560
rect 579 1362 613 1422
rect 739 1362 773 1422
rect 7268 1362 7302 1422
rect 7428 1362 7462 1422
rect 579 1224 613 1284
rect 739 1224 773 1284
rect 7268 1224 7302 1284
rect 7428 1224 7462 1284
rect 579 1086 613 1146
rect 739 1086 773 1146
rect 7268 1086 7302 1146
rect 7428 1086 7462 1146
rect 579 948 613 1008
rect 739 948 773 1008
rect 7268 948 7302 1008
rect 7428 948 7462 1008
rect 579 810 613 870
rect 739 810 773 870
rect 7268 810 7302 870
rect 7428 810 7462 870
rect 579 672 613 732
rect 739 672 773 732
rect 7268 672 7302 732
rect 7428 672 7462 732
rect 6076 216 6110 276
rect 6236 216 6270 276
rect 12831 216 12865 276
rect 12991 216 13025 276
rect 6076 78 6110 138
rect 6236 78 6270 138
rect 12831 78 12865 138
rect 12991 78 13025 138
rect 6076 -60 6110 0
rect 6236 -60 6270 0
rect 12831 -60 12865 0
rect 12991 -60 13025 0
rect 6076 -198 6110 -138
rect 6236 -198 6270 -138
rect 12831 -198 12865 -138
rect 12991 -198 13025 -138
rect 6076 -336 6110 -276
rect 6236 -336 6270 -276
rect 12831 -336 12865 -276
rect 12991 -336 13025 -276
rect 6076 -474 6110 -414
rect 6236 -474 6270 -414
rect 12831 -474 12865 -414
rect 12991 -474 13025 -414
rect 6076 -612 6110 -552
rect 6236 -612 6270 -552
rect 12831 -612 12865 -552
rect 12991 -612 13025 -552
rect 338 -797 372 -737
rect 426 -797 460 -737
rect 6076 -750 6110 -690
rect 6236 -750 6270 -690
rect 7093 -797 7127 -737
rect 7181 -797 7215 -737
rect 12831 -750 12865 -690
rect 12991 -750 13025 -690
rect 146 -935 180 -875
rect 242 -935 276 -875
rect 338 -935 372 -875
rect 426 -935 460 -875
rect 988 -934 1022 -874
rect 1077 -934 1111 -874
rect 1720 -934 1754 -874
rect 1826 -934 1860 -874
rect 1932 -934 1966 -874
rect 3058 -934 3092 -874
rect 3166 -934 3200 -874
rect 3270 -934 3304 -874
rect 4270 -934 4304 -874
rect 4377 -934 4411 -874
rect 4482 -934 4516 -874
rect 5126 -934 5160 -874
rect 5214 -934 5248 -874
rect 6901 -935 6935 -875
rect 6997 -935 7031 -875
rect 7093 -935 7127 -875
rect 7181 -935 7215 -875
rect 7743 -934 7777 -874
rect 7832 -934 7866 -874
rect 8475 -934 8509 -874
rect 8581 -934 8615 -874
rect 8687 -934 8721 -874
rect 9813 -934 9847 -874
rect 9921 -934 9955 -874
rect 10025 -934 10059 -874
rect 11025 -934 11059 -874
rect 11132 -934 11166 -874
rect 11237 -934 11271 -874
rect 11881 -934 11915 -874
rect 11969 -934 12003 -874
rect 6403 -1242 6437 -1208
rect 6403 -1310 6437 -1276
rect 6487 -1242 6521 -1208
rect 6487 -1310 6521 -1276
rect 6593 -1242 6627 -1208
rect 6593 -1310 6627 -1276
rect 6677 -1242 6711 -1208
rect 6677 -1310 6711 -1276
rect 13158 -1242 13192 -1208
rect 13158 -1310 13192 -1276
rect 13242 -1242 13276 -1208
rect 13242 -1310 13276 -1276
rect 13348 -1242 13382 -1208
rect 13348 -1310 13382 -1276
rect 13432 -1242 13466 -1208
rect 13432 -1310 13466 -1276
<< pdiffc >>
rect 625 3165 659 3225
rect 713 3165 747 3225
rect 7314 3165 7348 3225
rect 7402 3165 7436 3225
rect 625 3027 659 3087
rect 713 3027 747 3087
rect 7314 3027 7348 3087
rect 7402 3027 7436 3087
rect 625 2889 659 2949
rect 713 2889 747 2949
rect 7314 2889 7348 2949
rect 7402 2889 7436 2949
rect 625 2751 659 2811
rect 713 2751 747 2811
rect 7314 2751 7348 2811
rect 7402 2751 7436 2811
rect 625 2613 659 2673
rect 713 2613 747 2673
rect 138 2544 172 2578
rect 138 2476 172 2510
rect 138 2408 172 2442
rect 222 2544 256 2578
rect 222 2476 256 2510
rect 222 2408 256 2442
rect 328 2544 362 2578
rect 328 2476 362 2510
rect 328 2408 362 2442
rect 412 2544 446 2578
rect 7314 2613 7348 2673
rect 7402 2613 7436 2673
rect 412 2476 446 2510
rect 625 2475 659 2535
rect 713 2475 747 2535
rect 6827 2544 6861 2578
rect 6827 2476 6861 2510
rect 412 2408 446 2442
rect 6827 2408 6861 2442
rect 6911 2544 6945 2578
rect 6911 2476 6945 2510
rect 6911 2408 6945 2442
rect 7017 2544 7051 2578
rect 7017 2476 7051 2510
rect 7017 2408 7051 2442
rect 7101 2544 7135 2578
rect 7101 2476 7135 2510
rect 7314 2475 7348 2535
rect 7402 2475 7436 2535
rect 7101 2408 7135 2442
rect 6389 2164 6423 2224
rect 6477 2164 6511 2224
rect 13078 2164 13112 2224
rect 13166 2164 13200 2224
rect 1246 2023 1280 2083
rect 1334 2023 1368 2083
rect 1978 2023 2012 2083
rect 2083 2023 2117 2083
rect 2192 2023 2226 2083
rect 3190 2023 3224 2083
rect 3294 2023 3328 2083
rect 3404 2023 3438 2083
rect 4402 2023 4436 2083
rect 4507 2023 4541 2083
rect 4616 2023 4650 2083
rect 5614 2023 5648 2083
rect 5721 2023 5755 2083
rect 5828 2023 5862 2083
rect 6389 2026 6423 2086
rect 6477 2026 6511 2086
rect 6573 2026 6607 2086
rect 6669 2026 6703 2086
rect 7935 2023 7969 2083
rect 8023 2023 8057 2083
rect 8667 2023 8701 2083
rect 8772 2023 8806 2083
rect 8881 2023 8915 2083
rect 9879 2023 9913 2083
rect 9983 2023 10017 2083
rect 10093 2023 10127 2083
rect 11091 2023 11125 2083
rect 11196 2023 11230 2083
rect 11305 2023 11339 2083
rect 12303 2023 12337 2083
rect 12410 2023 12444 2083
rect 12517 2023 12551 2083
rect 13078 2026 13112 2086
rect 13166 2026 13200 2086
rect 13262 2026 13296 2086
rect 13358 2026 13392 2086
rect 146 -1138 180 -1078
rect 242 -1138 276 -1078
rect 338 -1138 372 -1078
rect 426 -1138 460 -1078
rect 987 -1135 1021 -1075
rect 1094 -1135 1128 -1075
rect 1201 -1135 1235 -1075
rect 2199 -1135 2233 -1075
rect 2308 -1135 2342 -1075
rect 2413 -1135 2447 -1075
rect 3411 -1135 3445 -1075
rect 3521 -1135 3555 -1075
rect 3625 -1135 3659 -1075
rect 4623 -1135 4657 -1075
rect 4732 -1135 4766 -1075
rect 4837 -1135 4871 -1075
rect 5481 -1135 5515 -1075
rect 5569 -1135 5603 -1075
rect 6901 -1138 6935 -1078
rect 6997 -1138 7031 -1078
rect 7093 -1138 7127 -1078
rect 7181 -1138 7215 -1078
rect 7742 -1135 7776 -1075
rect 7849 -1135 7883 -1075
rect 7956 -1135 7990 -1075
rect 8954 -1135 8988 -1075
rect 9063 -1135 9097 -1075
rect 9168 -1135 9202 -1075
rect 10166 -1135 10200 -1075
rect 10276 -1135 10310 -1075
rect 10380 -1135 10414 -1075
rect 11378 -1135 11412 -1075
rect 11487 -1135 11521 -1075
rect 11592 -1135 11626 -1075
rect 12236 -1135 12270 -1075
rect 12324 -1135 12358 -1075
rect 338 -1276 372 -1216
rect 426 -1276 460 -1216
rect 7093 -1276 7127 -1216
rect 7181 -1276 7215 -1216
rect 6403 -1494 6437 -1460
rect 6102 -1587 6136 -1527
rect 6190 -1587 6224 -1527
rect 6403 -1562 6437 -1528
rect 6403 -1630 6437 -1596
rect 6487 -1494 6521 -1460
rect 6487 -1562 6521 -1528
rect 6487 -1630 6521 -1596
rect 6593 -1494 6627 -1460
rect 6593 -1562 6627 -1528
rect 6593 -1630 6627 -1596
rect 6677 -1494 6711 -1460
rect 13158 -1494 13192 -1460
rect 6677 -1562 6711 -1528
rect 6677 -1630 6711 -1596
rect 12857 -1587 12891 -1527
rect 12945 -1587 12979 -1527
rect 13158 -1562 13192 -1528
rect 6102 -1725 6136 -1665
rect 6190 -1725 6224 -1665
rect 13158 -1630 13192 -1596
rect 13242 -1494 13276 -1460
rect 13242 -1562 13276 -1528
rect 13242 -1630 13276 -1596
rect 13348 -1494 13382 -1460
rect 13348 -1562 13382 -1528
rect 13348 -1630 13382 -1596
rect 13432 -1494 13466 -1460
rect 13432 -1562 13466 -1528
rect 13432 -1630 13466 -1596
rect 12857 -1725 12891 -1665
rect 12945 -1725 12979 -1665
rect 6102 -1863 6136 -1803
rect 6190 -1863 6224 -1803
rect 12857 -1863 12891 -1803
rect 12945 -1863 12979 -1803
rect 6102 -2001 6136 -1941
rect 6190 -2001 6224 -1941
rect 12857 -2001 12891 -1941
rect 12945 -2001 12979 -1941
rect 6102 -2139 6136 -2079
rect 6190 -2139 6224 -2079
rect 12857 -2139 12891 -2079
rect 12945 -2139 12979 -2079
rect 6102 -2277 6136 -2217
rect 6190 -2277 6224 -2217
rect 12857 -2277 12891 -2217
rect 12945 -2277 12979 -2217
<< poly >>
rect 671 3237 701 3267
rect 7360 3237 7390 3267
rect 671 3099 701 3153
rect 7360 3099 7390 3153
rect 671 2961 701 3015
rect 7360 2961 7390 3015
rect 671 2823 701 2877
rect 7360 2823 7390 2877
rect 671 2685 701 2739
rect 7360 2685 7390 2739
rect 182 2590 212 2616
rect 372 2590 402 2616
rect 671 2547 701 2601
rect 6871 2590 6901 2616
rect 7061 2590 7091 2616
rect 671 2432 701 2463
rect 653 2416 719 2432
rect 182 2358 212 2390
rect 126 2342 212 2358
rect 126 2308 142 2342
rect 176 2308 212 2342
rect 126 2292 212 2308
rect 182 2270 212 2292
rect 372 2358 402 2390
rect 653 2382 669 2416
rect 703 2382 719 2416
rect 7360 2547 7390 2601
rect 7360 2432 7390 2463
rect 7342 2416 7408 2432
rect 653 2366 719 2382
rect 6871 2358 6901 2390
rect 372 2342 458 2358
rect 372 2308 408 2342
rect 442 2308 458 2342
rect 372 2292 458 2308
rect 6815 2342 6901 2358
rect 6815 2308 6831 2342
rect 6865 2308 6901 2342
rect 6815 2292 6901 2308
rect 372 2270 402 2292
rect 6871 2270 6901 2292
rect 7061 2358 7091 2390
rect 7342 2382 7358 2416
rect 7392 2382 7408 2416
rect 7342 2366 7408 2382
rect 7061 2342 7147 2358
rect 7061 2308 7097 2342
rect 7131 2308 7147 2342
rect 7061 2292 7147 2308
rect 7061 2270 7091 2292
rect 6435 2236 6465 2267
rect 1274 2176 1340 2192
rect 1274 2142 1290 2176
rect 1324 2142 1340 2176
rect 182 2114 212 2140
rect 372 2114 402 2140
rect 1274 2126 1340 2142
rect 2006 2176 2072 2192
rect 2006 2142 2022 2176
rect 2056 2142 2072 2176
rect 2006 2126 2072 2142
rect 2132 2176 2198 2192
rect 2132 2142 2148 2176
rect 2182 2142 2198 2176
rect 2132 2126 2198 2142
rect 3218 2176 3284 2192
rect 3218 2142 3234 2176
rect 3268 2142 3284 2176
rect 3218 2126 3284 2142
rect 3344 2176 3410 2192
rect 3344 2142 3360 2176
rect 3394 2142 3410 2176
rect 3344 2126 3410 2142
rect 4430 2176 4496 2192
rect 4430 2142 4446 2176
rect 4480 2142 4496 2176
rect 4430 2126 4496 2142
rect 4556 2176 4622 2192
rect 4556 2142 4572 2176
rect 4606 2142 4622 2176
rect 4556 2126 4622 2142
rect 5642 2176 5708 2192
rect 5642 2142 5658 2176
rect 5692 2142 5708 2176
rect 5642 2126 5708 2142
rect 5768 2176 5834 2192
rect 5768 2142 5784 2176
rect 5818 2142 5834 2176
rect 5768 2126 5834 2142
rect 1292 2095 1322 2126
rect 2024 2095 2054 2126
rect 2150 2095 2180 2126
rect 3236 2095 3266 2126
rect 3362 2095 3392 2126
rect 4448 2095 4478 2126
rect 4574 2095 4604 2126
rect 5660 2095 5690 2126
rect 5786 2095 5816 2126
rect 6435 2098 6465 2152
rect 13124 2236 13154 2267
rect 7963 2176 8029 2192
rect 7963 2142 7979 2176
rect 8013 2142 8029 2176
rect 6527 2098 6557 2124
rect 6623 2098 6653 2129
rect 6871 2114 6901 2140
rect 7061 2114 7091 2140
rect 7963 2126 8029 2142
rect 8695 2176 8761 2192
rect 8695 2142 8711 2176
rect 8745 2142 8761 2176
rect 8695 2126 8761 2142
rect 8821 2176 8887 2192
rect 8821 2142 8837 2176
rect 8871 2142 8887 2176
rect 8821 2126 8887 2142
rect 9907 2176 9973 2192
rect 9907 2142 9923 2176
rect 9957 2142 9973 2176
rect 9907 2126 9973 2142
rect 10033 2176 10099 2192
rect 10033 2142 10049 2176
rect 10083 2142 10099 2176
rect 10033 2126 10099 2142
rect 11119 2176 11185 2192
rect 11119 2142 11135 2176
rect 11169 2142 11185 2176
rect 11119 2126 11185 2142
rect 11245 2176 11311 2192
rect 11245 2142 11261 2176
rect 11295 2142 11311 2176
rect 11245 2126 11311 2142
rect 12331 2176 12397 2192
rect 12331 2142 12347 2176
rect 12381 2142 12397 2176
rect 12331 2126 12397 2142
rect 12457 2176 12523 2192
rect 12457 2142 12473 2176
rect 12507 2142 12523 2176
rect 12457 2126 12523 2142
rect 7981 2095 8011 2126
rect 8713 2095 8743 2126
rect 8839 2095 8869 2126
rect 9925 2095 9955 2126
rect 10051 2095 10081 2126
rect 11137 2095 11167 2126
rect 11263 2095 11293 2126
rect 12349 2095 12379 2126
rect 12475 2095 12505 2126
rect 13124 2098 13154 2152
rect 13216 2098 13246 2124
rect 13312 2098 13342 2129
rect 1292 1983 1322 2011
rect 2024 1983 2054 2011
rect 2150 1983 2180 2011
rect 3236 1983 3266 2011
rect 3362 1983 3392 2011
rect 4448 1983 4478 2011
rect 4574 1983 4604 2011
rect 5660 1983 5690 2011
rect 5786 1983 5816 2011
rect 6435 1989 6465 2014
rect 6306 1969 6465 1989
rect 6527 1989 6557 2014
rect 6623 1989 6653 2014
rect 6527 1983 6653 1989
rect 7981 1983 8011 2011
rect 8713 1983 8743 2011
rect 8839 1983 8869 2011
rect 9925 1983 9955 2011
rect 10051 1983 10081 2011
rect 11137 1983 11167 2011
rect 11263 1983 11293 2011
rect 12349 1983 12379 2011
rect 12475 1983 12505 2011
rect 13124 1989 13154 2014
rect 6306 1935 6318 1969
rect 6352 1935 6465 1969
rect 1647 1894 1677 1920
rect 2379 1894 2409 1920
rect 2503 1894 2533 1920
rect 3591 1894 3621 1920
rect 3715 1894 3745 1920
rect 4929 1894 4959 1920
rect 5053 1894 5083 1920
rect 5785 1894 5815 1920
rect 6306 1916 6465 1935
rect 6509 1967 6653 1983
rect 6509 1933 6525 1967
rect 6559 1933 6653 1967
rect 6509 1917 6653 1933
rect 12995 1969 13154 1989
rect 13216 1989 13246 2014
rect 13312 1989 13342 2014
rect 13216 1983 13342 1989
rect 12995 1935 13007 1969
rect 13041 1935 13154 1969
rect 6435 1895 6465 1916
rect 6527 1910 6653 1917
rect 6527 1895 6557 1910
rect 6623 1895 6653 1910
rect 8336 1894 8366 1920
rect 9068 1894 9098 1920
rect 9192 1894 9222 1920
rect 10280 1894 10310 1920
rect 10404 1894 10434 1920
rect 11618 1894 11648 1920
rect 11742 1894 11772 1920
rect 12474 1894 12504 1920
rect 12995 1916 13154 1935
rect 13198 1967 13342 1983
rect 13198 1933 13214 1967
rect 13248 1933 13342 1967
rect 13198 1917 13342 1933
rect 13124 1895 13154 1916
rect 13216 1910 13342 1917
rect 13216 1895 13246 1910
rect 13312 1895 13342 1910
rect 643 1782 709 1798
rect 1647 1788 1677 1810
rect 2379 1788 2409 1810
rect 2503 1788 2533 1810
rect 3591 1788 3621 1810
rect 3715 1788 3745 1810
rect 4929 1788 4959 1810
rect 5053 1788 5083 1810
rect 5785 1788 5815 1810
rect 643 1755 659 1782
rect 625 1748 659 1755
rect 693 1755 709 1782
rect 1629 1772 1695 1788
rect 693 1748 727 1755
rect 625 1725 727 1748
rect 625 1710 655 1725
rect 697 1710 727 1725
rect 1629 1738 1645 1772
rect 1679 1738 1695 1772
rect 1629 1722 1695 1738
rect 2361 1772 2427 1788
rect 2361 1738 2377 1772
rect 2411 1738 2427 1772
rect 2361 1722 2427 1738
rect 2485 1772 2551 1788
rect 2485 1738 2501 1772
rect 2535 1738 2551 1772
rect 2485 1722 2551 1738
rect 3573 1772 3639 1788
rect 3573 1738 3589 1772
rect 3623 1738 3639 1772
rect 3573 1722 3639 1738
rect 3697 1772 3763 1788
rect 3697 1738 3713 1772
rect 3747 1738 3763 1772
rect 3697 1722 3763 1738
rect 4911 1772 4977 1788
rect 4911 1738 4927 1772
rect 4961 1738 4977 1772
rect 4911 1722 4977 1738
rect 5035 1772 5101 1788
rect 5035 1738 5051 1772
rect 5085 1738 5101 1772
rect 5035 1722 5101 1738
rect 5767 1772 5833 1788
rect 5767 1738 5783 1772
rect 5817 1738 5833 1772
rect 6435 1757 6465 1811
rect 6527 1785 6557 1811
rect 6623 1785 6653 1811
rect 7332 1782 7398 1798
rect 8336 1788 8366 1810
rect 9068 1788 9098 1810
rect 9192 1788 9222 1810
rect 10280 1788 10310 1810
rect 10404 1788 10434 1810
rect 11618 1788 11648 1810
rect 11742 1788 11772 1810
rect 12474 1788 12504 1810
rect 5767 1722 5833 1738
rect 7332 1755 7348 1782
rect 7314 1748 7348 1755
rect 7382 1755 7398 1782
rect 8318 1772 8384 1788
rect 7382 1748 7416 1755
rect 7314 1725 7416 1748
rect 7314 1710 7344 1725
rect 7386 1710 7416 1725
rect 8318 1738 8334 1772
rect 8368 1738 8384 1772
rect 8318 1722 8384 1738
rect 9050 1772 9116 1788
rect 9050 1738 9066 1772
rect 9100 1738 9116 1772
rect 9050 1722 9116 1738
rect 9174 1772 9240 1788
rect 9174 1738 9190 1772
rect 9224 1738 9240 1772
rect 9174 1722 9240 1738
rect 10262 1772 10328 1788
rect 10262 1738 10278 1772
rect 10312 1738 10328 1772
rect 10262 1722 10328 1738
rect 10386 1772 10452 1788
rect 10386 1738 10402 1772
rect 10436 1738 10452 1772
rect 10386 1722 10452 1738
rect 11600 1772 11666 1788
rect 11600 1738 11616 1772
rect 11650 1738 11666 1772
rect 11600 1722 11666 1738
rect 11724 1772 11790 1788
rect 11724 1738 11740 1772
rect 11774 1738 11790 1772
rect 11724 1722 11790 1738
rect 12456 1772 12522 1788
rect 12456 1738 12472 1772
rect 12506 1738 12522 1772
rect 13124 1757 13154 1811
rect 13216 1785 13246 1811
rect 13312 1785 13342 1811
rect 12456 1722 12522 1738
rect 6435 1646 6465 1673
rect 13124 1646 13154 1673
rect 625 1572 655 1626
rect 697 1572 727 1626
rect 7314 1572 7344 1626
rect 7386 1572 7416 1626
rect 625 1434 655 1488
rect 697 1434 727 1488
rect 7314 1434 7344 1488
rect 7386 1434 7416 1488
rect 625 1296 655 1350
rect 697 1296 727 1350
rect 7314 1296 7344 1350
rect 7386 1296 7416 1350
rect 625 1158 655 1212
rect 697 1158 727 1212
rect 7314 1158 7344 1212
rect 7386 1158 7416 1212
rect 625 1020 655 1074
rect 697 1020 727 1074
rect 7314 1020 7344 1074
rect 7386 1020 7416 1074
rect 625 882 655 936
rect 697 882 727 936
rect 7314 882 7344 936
rect 7386 882 7416 936
rect 625 744 655 798
rect 697 744 727 798
rect 7314 744 7344 798
rect 7386 744 7416 798
rect 625 634 655 660
rect 697 634 727 660
rect 7314 634 7344 660
rect 7386 634 7416 660
rect 6122 288 6152 314
rect 6194 288 6224 314
rect 12877 288 12907 314
rect 12949 288 12979 314
rect 6122 150 6152 204
rect 6194 150 6224 204
rect 12877 150 12907 204
rect 12949 150 12979 204
rect 6122 12 6152 66
rect 6194 12 6224 66
rect 12877 12 12907 66
rect 12949 12 12979 66
rect 6122 -126 6152 -72
rect 6194 -126 6224 -72
rect 12877 -126 12907 -72
rect 12949 -126 12979 -72
rect 6122 -264 6152 -210
rect 6194 -264 6224 -210
rect 12877 -264 12907 -210
rect 12949 -264 12979 -210
rect 6122 -402 6152 -348
rect 6194 -402 6224 -348
rect 12877 -402 12907 -348
rect 12949 -402 12979 -348
rect 6122 -540 6152 -486
rect 6194 -540 6224 -486
rect 12877 -540 12907 -486
rect 12949 -540 12979 -486
rect 6122 -678 6152 -624
rect 6194 -678 6224 -624
rect 12877 -678 12907 -624
rect 12949 -678 12979 -624
rect 384 -725 414 -698
rect 7139 -725 7169 -698
rect 1016 -790 1082 -774
rect 196 -863 226 -837
rect 292 -863 322 -837
rect 384 -863 414 -809
rect 1016 -824 1032 -790
rect 1066 -824 1082 -790
rect 1016 -840 1082 -824
rect 1748 -790 1814 -774
rect 1748 -824 1764 -790
rect 1798 -824 1814 -790
rect 1748 -840 1814 -824
rect 1872 -790 1938 -774
rect 1872 -824 1888 -790
rect 1922 -824 1938 -790
rect 1872 -840 1938 -824
rect 3086 -790 3152 -774
rect 3086 -824 3102 -790
rect 3136 -824 3152 -790
rect 3086 -840 3152 -824
rect 3210 -790 3276 -774
rect 3210 -824 3226 -790
rect 3260 -824 3276 -790
rect 3210 -840 3276 -824
rect 4298 -790 4364 -774
rect 4298 -824 4314 -790
rect 4348 -824 4364 -790
rect 4298 -840 4364 -824
rect 4422 -790 4488 -774
rect 4422 -824 4438 -790
rect 4472 -824 4488 -790
rect 4422 -840 4488 -824
rect 5154 -790 5220 -774
rect 5154 -824 5170 -790
rect 5204 -824 5220 -790
rect 6122 -777 6152 -762
rect 6194 -777 6224 -762
rect 6122 -800 6224 -777
rect 6122 -807 6156 -800
rect 5154 -840 5220 -824
rect 6140 -834 6156 -807
rect 6190 -807 6224 -800
rect 6190 -834 6206 -807
rect 7771 -790 7837 -774
rect 1034 -862 1064 -840
rect 1766 -862 1796 -840
rect 1890 -862 1920 -840
rect 3104 -862 3134 -840
rect 3228 -862 3258 -840
rect 4316 -862 4346 -840
rect 4440 -862 4470 -840
rect 5172 -862 5202 -840
rect 6140 -850 6206 -834
rect 6951 -863 6981 -837
rect 7047 -863 7077 -837
rect 7139 -863 7169 -809
rect 7771 -824 7787 -790
rect 7821 -824 7837 -790
rect 7771 -840 7837 -824
rect 8503 -790 8569 -774
rect 8503 -824 8519 -790
rect 8553 -824 8569 -790
rect 8503 -840 8569 -824
rect 8627 -790 8693 -774
rect 8627 -824 8643 -790
rect 8677 -824 8693 -790
rect 8627 -840 8693 -824
rect 9841 -790 9907 -774
rect 9841 -824 9857 -790
rect 9891 -824 9907 -790
rect 9841 -840 9907 -824
rect 9965 -790 10031 -774
rect 9965 -824 9981 -790
rect 10015 -824 10031 -790
rect 9965 -840 10031 -824
rect 11053 -790 11119 -774
rect 11053 -824 11069 -790
rect 11103 -824 11119 -790
rect 11053 -840 11119 -824
rect 11177 -790 11243 -774
rect 11177 -824 11193 -790
rect 11227 -824 11243 -790
rect 11177 -840 11243 -824
rect 11909 -790 11975 -774
rect 11909 -824 11925 -790
rect 11959 -824 11975 -790
rect 12877 -777 12907 -762
rect 12949 -777 12979 -762
rect 12877 -800 12979 -777
rect 12877 -807 12911 -800
rect 11909 -840 11975 -824
rect 12895 -834 12911 -807
rect 12945 -807 12979 -800
rect 12945 -834 12961 -807
rect 7789 -862 7819 -840
rect 8521 -862 8551 -840
rect 8645 -862 8675 -840
rect 9859 -862 9889 -840
rect 9983 -862 10013 -840
rect 11071 -862 11101 -840
rect 11195 -862 11225 -840
rect 11927 -862 11957 -840
rect 12895 -850 12961 -834
rect 196 -962 226 -947
rect 292 -962 322 -947
rect 196 -969 322 -962
rect 384 -968 414 -947
rect 196 -985 340 -969
rect 196 -1019 290 -985
rect 324 -1019 340 -985
rect 196 -1035 340 -1019
rect 384 -987 543 -968
rect 1034 -972 1064 -946
rect 1766 -972 1796 -946
rect 1890 -972 1920 -946
rect 3104 -972 3134 -946
rect 3228 -972 3258 -946
rect 4316 -972 4346 -946
rect 4440 -972 4470 -946
rect 5172 -972 5202 -946
rect 6951 -962 6981 -947
rect 7047 -962 7077 -947
rect 6951 -969 7077 -962
rect 7139 -968 7169 -947
rect 384 -1021 497 -987
rect 531 -1021 543 -987
rect 196 -1041 322 -1035
rect 196 -1066 226 -1041
rect 292 -1066 322 -1041
rect 384 -1041 543 -1021
rect 6951 -985 7095 -969
rect 6951 -1019 7045 -985
rect 7079 -1019 7095 -985
rect 6951 -1035 7095 -1019
rect 7139 -987 7298 -968
rect 7789 -972 7819 -946
rect 8521 -972 8551 -946
rect 8645 -972 8675 -946
rect 9859 -972 9889 -946
rect 9983 -972 10013 -946
rect 11071 -972 11101 -946
rect 11195 -972 11225 -946
rect 11927 -972 11957 -946
rect 7139 -1021 7252 -987
rect 7286 -1021 7298 -987
rect 384 -1066 414 -1041
rect 1033 -1063 1063 -1035
rect 1159 -1063 1189 -1035
rect 2245 -1063 2275 -1035
rect 2371 -1063 2401 -1035
rect 3457 -1063 3487 -1035
rect 3583 -1063 3613 -1035
rect 4669 -1063 4699 -1035
rect 4795 -1063 4825 -1035
rect 5527 -1063 5557 -1035
rect 6951 -1041 7077 -1035
rect 6951 -1066 6981 -1041
rect 7047 -1066 7077 -1041
rect 7139 -1041 7298 -1021
rect 7139 -1066 7169 -1041
rect 7788 -1063 7818 -1035
rect 7914 -1063 7944 -1035
rect 9000 -1063 9030 -1035
rect 9126 -1063 9156 -1035
rect 10212 -1063 10242 -1035
rect 10338 -1063 10368 -1035
rect 11424 -1063 11454 -1035
rect 11550 -1063 11580 -1035
rect 12282 -1063 12312 -1035
rect 196 -1181 226 -1150
rect 292 -1176 322 -1150
rect 384 -1204 414 -1150
rect 1033 -1178 1063 -1147
rect 1159 -1178 1189 -1147
rect 2245 -1178 2275 -1147
rect 2371 -1178 2401 -1147
rect 3457 -1178 3487 -1147
rect 3583 -1178 3613 -1147
rect 4669 -1178 4699 -1147
rect 4795 -1178 4825 -1147
rect 5527 -1178 5557 -1147
rect 1015 -1194 1081 -1178
rect 1015 -1228 1031 -1194
rect 1065 -1228 1081 -1194
rect 1015 -1244 1081 -1228
rect 1141 -1194 1207 -1178
rect 1141 -1228 1157 -1194
rect 1191 -1228 1207 -1194
rect 1141 -1244 1207 -1228
rect 2227 -1194 2293 -1178
rect 2227 -1228 2243 -1194
rect 2277 -1228 2293 -1194
rect 2227 -1244 2293 -1228
rect 2353 -1194 2419 -1178
rect 2353 -1228 2369 -1194
rect 2403 -1228 2419 -1194
rect 2353 -1244 2419 -1228
rect 3439 -1194 3505 -1178
rect 3439 -1228 3455 -1194
rect 3489 -1228 3505 -1194
rect 3439 -1244 3505 -1228
rect 3565 -1194 3631 -1178
rect 3565 -1228 3581 -1194
rect 3615 -1228 3631 -1194
rect 3565 -1244 3631 -1228
rect 4651 -1194 4717 -1178
rect 4651 -1228 4667 -1194
rect 4701 -1228 4717 -1194
rect 4651 -1244 4717 -1228
rect 4777 -1194 4843 -1178
rect 4777 -1228 4793 -1194
rect 4827 -1228 4843 -1194
rect 4777 -1244 4843 -1228
rect 5509 -1194 5575 -1178
rect 6447 -1192 6477 -1166
rect 6637 -1192 6667 -1166
rect 6951 -1181 6981 -1150
rect 7047 -1176 7077 -1150
rect 5509 -1228 5525 -1194
rect 5559 -1228 5575 -1194
rect 5509 -1244 5575 -1228
rect 384 -1319 414 -1288
rect 7139 -1204 7169 -1150
rect 7788 -1178 7818 -1147
rect 7914 -1178 7944 -1147
rect 9000 -1178 9030 -1147
rect 9126 -1178 9156 -1147
rect 10212 -1178 10242 -1147
rect 10338 -1178 10368 -1147
rect 11424 -1178 11454 -1147
rect 11550 -1178 11580 -1147
rect 12282 -1178 12312 -1147
rect 7770 -1194 7836 -1178
rect 7770 -1228 7786 -1194
rect 7820 -1228 7836 -1194
rect 7770 -1244 7836 -1228
rect 7896 -1194 7962 -1178
rect 7896 -1228 7912 -1194
rect 7946 -1228 7962 -1194
rect 7896 -1244 7962 -1228
rect 8982 -1194 9048 -1178
rect 8982 -1228 8998 -1194
rect 9032 -1228 9048 -1194
rect 8982 -1244 9048 -1228
rect 9108 -1194 9174 -1178
rect 9108 -1228 9124 -1194
rect 9158 -1228 9174 -1194
rect 9108 -1244 9174 -1228
rect 10194 -1194 10260 -1178
rect 10194 -1228 10210 -1194
rect 10244 -1228 10260 -1194
rect 10194 -1244 10260 -1228
rect 10320 -1194 10386 -1178
rect 10320 -1228 10336 -1194
rect 10370 -1228 10386 -1194
rect 10320 -1244 10386 -1228
rect 11406 -1194 11472 -1178
rect 11406 -1228 11422 -1194
rect 11456 -1228 11472 -1194
rect 11406 -1244 11472 -1228
rect 11532 -1194 11598 -1178
rect 11532 -1228 11548 -1194
rect 11582 -1228 11598 -1194
rect 11532 -1244 11598 -1228
rect 12264 -1194 12330 -1178
rect 13202 -1192 13232 -1166
rect 13392 -1192 13422 -1166
rect 12264 -1228 12280 -1194
rect 12314 -1228 12330 -1194
rect 12264 -1244 12330 -1228
rect 7139 -1319 7169 -1288
rect 6447 -1344 6477 -1322
rect 6391 -1360 6477 -1344
rect 6391 -1394 6407 -1360
rect 6441 -1394 6477 -1360
rect 6391 -1410 6477 -1394
rect 6130 -1434 6196 -1418
rect 6130 -1468 6146 -1434
rect 6180 -1468 6196 -1434
rect 6447 -1442 6477 -1410
rect 6637 -1344 6667 -1322
rect 13202 -1344 13232 -1322
rect 6637 -1360 6723 -1344
rect 6637 -1394 6673 -1360
rect 6707 -1394 6723 -1360
rect 6637 -1410 6723 -1394
rect 13146 -1360 13232 -1344
rect 13146 -1394 13162 -1360
rect 13196 -1394 13232 -1360
rect 13146 -1410 13232 -1394
rect 6637 -1442 6667 -1410
rect 12885 -1434 12951 -1418
rect 6130 -1484 6196 -1468
rect 6148 -1515 6178 -1484
rect 6148 -1653 6178 -1599
rect 12885 -1468 12901 -1434
rect 12935 -1468 12951 -1434
rect 13202 -1442 13232 -1410
rect 13392 -1344 13422 -1322
rect 13392 -1360 13478 -1344
rect 13392 -1394 13428 -1360
rect 13462 -1394 13478 -1360
rect 13392 -1410 13478 -1394
rect 13392 -1442 13422 -1410
rect 12885 -1484 12951 -1468
rect 12903 -1515 12933 -1484
rect 6447 -1668 6477 -1642
rect 6637 -1668 6667 -1642
rect 12903 -1653 12933 -1599
rect 13202 -1668 13232 -1642
rect 13392 -1668 13422 -1642
rect 6148 -1791 6178 -1737
rect 12903 -1791 12933 -1737
rect 6148 -1929 6178 -1875
rect 12903 -1929 12933 -1875
rect 6148 -2067 6178 -2013
rect 12903 -2067 12933 -2013
rect 6148 -2205 6178 -2151
rect 12903 -2205 12933 -2151
rect 6148 -2319 6178 -2289
rect 12903 -2319 12933 -2289
<< polycont >>
rect 142 2308 176 2342
rect 669 2382 703 2416
rect 408 2308 442 2342
rect 6831 2308 6865 2342
rect 7358 2382 7392 2416
rect 7097 2308 7131 2342
rect 1290 2142 1324 2176
rect 2022 2142 2056 2176
rect 2148 2142 2182 2176
rect 3234 2142 3268 2176
rect 3360 2142 3394 2176
rect 4446 2142 4480 2176
rect 4572 2142 4606 2176
rect 5658 2142 5692 2176
rect 5784 2142 5818 2176
rect 7979 2142 8013 2176
rect 8711 2142 8745 2176
rect 8837 2142 8871 2176
rect 9923 2142 9957 2176
rect 10049 2142 10083 2176
rect 11135 2142 11169 2176
rect 11261 2142 11295 2176
rect 12347 2142 12381 2176
rect 12473 2142 12507 2176
rect 6318 1935 6352 1969
rect 6525 1933 6559 1967
rect 13007 1935 13041 1969
rect 13214 1933 13248 1967
rect 659 1748 693 1782
rect 1645 1738 1679 1772
rect 2377 1738 2411 1772
rect 2501 1738 2535 1772
rect 3589 1738 3623 1772
rect 3713 1738 3747 1772
rect 4927 1738 4961 1772
rect 5051 1738 5085 1772
rect 5783 1738 5817 1772
rect 7348 1748 7382 1782
rect 8334 1738 8368 1772
rect 9066 1738 9100 1772
rect 9190 1738 9224 1772
rect 10278 1738 10312 1772
rect 10402 1738 10436 1772
rect 11616 1738 11650 1772
rect 11740 1738 11774 1772
rect 12472 1738 12506 1772
rect 1032 -824 1066 -790
rect 1764 -824 1798 -790
rect 1888 -824 1922 -790
rect 3102 -824 3136 -790
rect 3226 -824 3260 -790
rect 4314 -824 4348 -790
rect 4438 -824 4472 -790
rect 5170 -824 5204 -790
rect 6156 -834 6190 -800
rect 7787 -824 7821 -790
rect 8519 -824 8553 -790
rect 8643 -824 8677 -790
rect 9857 -824 9891 -790
rect 9981 -824 10015 -790
rect 11069 -824 11103 -790
rect 11193 -824 11227 -790
rect 11925 -824 11959 -790
rect 12911 -834 12945 -800
rect 290 -1019 324 -985
rect 497 -1021 531 -987
rect 7045 -1019 7079 -985
rect 7252 -1021 7286 -987
rect 1031 -1228 1065 -1194
rect 1157 -1228 1191 -1194
rect 2243 -1228 2277 -1194
rect 2369 -1228 2403 -1194
rect 3455 -1228 3489 -1194
rect 3581 -1228 3615 -1194
rect 4667 -1228 4701 -1194
rect 4793 -1228 4827 -1194
rect 5525 -1228 5559 -1194
rect 7786 -1228 7820 -1194
rect 7912 -1228 7946 -1194
rect 8998 -1228 9032 -1194
rect 9124 -1228 9158 -1194
rect 10210 -1228 10244 -1194
rect 10336 -1228 10370 -1194
rect 11422 -1228 11456 -1194
rect 11548 -1228 11582 -1194
rect 12280 -1228 12314 -1194
rect 6407 -1394 6441 -1360
rect 6146 -1468 6180 -1434
rect 6673 -1394 6707 -1360
rect 13162 -1394 13196 -1360
rect 12901 -1468 12935 -1434
rect 13428 -1394 13462 -1360
<< locali >>
rect 625 3225 659 3241
rect 625 3149 659 3165
rect 713 3225 747 3241
rect 713 3149 747 3165
rect 7314 3225 7348 3241
rect 7314 3149 7348 3165
rect 7402 3225 7436 3241
rect 7402 3149 7436 3165
rect 625 3087 659 3103
rect 625 3011 659 3027
rect 713 3087 747 3103
rect 713 3011 747 3027
rect 7314 3087 7348 3103
rect 7314 3011 7348 3027
rect 7402 3087 7436 3103
rect 7402 3011 7436 3027
rect 625 2949 659 2965
rect 625 2873 659 2889
rect 713 2949 747 2965
rect 713 2873 747 2889
rect 7314 2949 7348 2965
rect 7314 2873 7348 2889
rect 7402 2949 7436 2965
rect 7402 2873 7436 2889
rect 625 2811 659 2827
rect 625 2735 659 2751
rect 713 2811 747 2827
rect 713 2735 747 2751
rect 7314 2811 7348 2827
rect 7314 2735 7348 2751
rect 7402 2811 7436 2827
rect 7402 2735 7436 2751
rect 625 2673 659 2689
rect 62 2620 91 2654
rect 125 2620 183 2654
rect 217 2620 275 2654
rect 309 2620 367 2654
rect 401 2620 459 2654
rect 493 2620 522 2654
rect 130 2578 172 2620
rect 130 2544 138 2578
rect 130 2510 172 2544
rect 130 2476 138 2510
rect 130 2442 172 2476
rect 130 2408 138 2442
rect 130 2392 172 2408
rect 206 2578 272 2586
rect 206 2544 222 2578
rect 256 2544 272 2578
rect 206 2511 272 2544
rect 206 2477 219 2511
rect 253 2510 272 2511
rect 206 2476 222 2477
rect 256 2476 272 2510
rect 206 2442 272 2476
rect 206 2408 222 2442
rect 256 2408 272 2442
rect 206 2390 272 2408
rect 126 2346 192 2356
rect 126 2312 138 2346
rect 172 2342 192 2346
rect 126 2308 142 2312
rect 176 2308 192 2342
rect 126 2258 172 2274
rect 226 2270 272 2390
rect 126 2224 138 2258
rect 126 2190 172 2224
rect 126 2156 138 2190
rect 126 2110 172 2156
rect 206 2258 272 2270
rect 206 2224 222 2258
rect 256 2224 272 2258
rect 206 2190 272 2224
rect 206 2156 222 2190
rect 256 2156 272 2190
rect 206 2144 272 2156
rect 312 2578 378 2586
rect 312 2544 328 2578
rect 362 2544 378 2578
rect 312 2510 378 2544
rect 312 2476 328 2510
rect 362 2476 378 2510
rect 312 2456 378 2476
rect 312 2408 328 2456
rect 362 2408 378 2456
rect 312 2390 378 2408
rect 412 2578 454 2620
rect 625 2597 659 2613
rect 713 2673 747 2689
rect 7314 2673 7348 2689
rect 6751 2620 6780 2654
rect 6814 2620 6872 2654
rect 6906 2620 6964 2654
rect 6998 2620 7056 2654
rect 7090 2620 7148 2654
rect 7182 2620 7211 2654
rect 713 2597 747 2613
rect 446 2544 454 2578
rect 6819 2578 6861 2620
rect 412 2510 454 2544
rect 446 2476 454 2510
rect 412 2442 454 2476
rect 625 2535 659 2551
rect 625 2459 659 2475
rect 713 2535 747 2551
rect 713 2459 747 2475
rect 6819 2544 6827 2578
rect 6819 2510 6861 2544
rect 6819 2476 6827 2510
rect 446 2408 454 2442
rect 6819 2442 6861 2476
rect 412 2392 454 2408
rect 312 2270 358 2390
rect 653 2382 669 2416
rect 703 2382 719 2416
rect 6819 2408 6827 2442
rect 6819 2392 6861 2408
rect 6895 2578 6961 2586
rect 6895 2544 6911 2578
rect 6945 2544 6961 2578
rect 6895 2511 6961 2544
rect 6895 2477 6908 2511
rect 6942 2510 6961 2511
rect 6895 2476 6911 2477
rect 6945 2476 6961 2510
rect 6895 2442 6961 2476
rect 6895 2408 6911 2442
rect 6945 2408 6961 2442
rect 6895 2390 6961 2408
rect 392 2345 458 2356
rect 392 2342 412 2345
rect 392 2308 408 2342
rect 446 2311 458 2345
rect 442 2308 458 2311
rect 579 2346 628 2358
rect 579 2312 588 2346
rect 622 2341 628 2346
rect 6815 2346 6881 2356
rect 622 2312 874 2341
rect 579 2306 874 2312
rect 6815 2312 6827 2346
rect 6861 2342 6881 2346
rect 6815 2308 6831 2312
rect 6865 2308 6881 2342
rect 579 2299 628 2306
rect 839 2283 874 2306
rect 312 2258 378 2270
rect 312 2224 328 2258
rect 362 2224 378 2258
rect 312 2190 378 2224
rect 312 2156 328 2190
rect 362 2156 378 2190
rect 312 2144 378 2156
rect 412 2258 458 2274
rect 839 2271 888 2283
rect 446 2224 458 2258
rect 412 2190 458 2224
rect 580 2253 629 2265
rect 580 2219 589 2253
rect 623 2219 790 2253
rect 839 2237 848 2271
rect 882 2237 888 2271
rect 6815 2258 6861 2274
rect 6915 2270 6961 2390
rect 839 2224 888 2237
rect 6389 2224 6423 2240
rect 580 2206 629 2219
rect 446 2156 458 2190
rect 412 2110 458 2156
rect 749 2177 790 2219
rect 840 2178 889 2190
rect 840 2177 849 2178
rect 749 2144 849 2177
rect 883 2144 889 2178
rect 749 2143 889 2144
rect 840 2131 889 2143
rect 1274 2142 1290 2176
rect 1324 2142 1340 2176
rect 2006 2142 2022 2176
rect 2056 2142 2072 2176
rect 2132 2142 2148 2176
rect 2182 2142 2198 2176
rect 3218 2142 3234 2176
rect 3268 2142 3284 2176
rect 3344 2142 3360 2176
rect 3394 2142 3410 2176
rect 4430 2142 4446 2176
rect 4480 2142 4496 2176
rect 4556 2142 4572 2176
rect 4606 2142 4622 2176
rect 5642 2142 5658 2176
rect 5692 2142 5708 2176
rect 5768 2142 5784 2176
rect 5818 2142 5834 2176
rect 6389 2148 6423 2164
rect 6477 2224 6511 2240
rect 6477 2148 6511 2164
rect 6815 2224 6827 2258
rect 6815 2190 6861 2224
rect 6815 2156 6827 2190
rect 6815 2110 6861 2156
rect 6895 2258 6961 2270
rect 6895 2224 6911 2258
rect 6945 2224 6961 2258
rect 6895 2190 6961 2224
rect 6895 2156 6911 2190
rect 6945 2156 6961 2190
rect 6895 2144 6961 2156
rect 7001 2578 7067 2586
rect 7001 2544 7017 2578
rect 7051 2544 7067 2578
rect 7001 2510 7067 2544
rect 7001 2476 7017 2510
rect 7051 2476 7067 2510
rect 7001 2456 7067 2476
rect 7001 2408 7017 2456
rect 7051 2408 7067 2456
rect 7001 2390 7067 2408
rect 7101 2578 7143 2620
rect 7314 2597 7348 2613
rect 7402 2673 7436 2689
rect 7402 2597 7436 2613
rect 7135 2544 7143 2578
rect 7101 2510 7143 2544
rect 7135 2476 7143 2510
rect 7101 2442 7143 2476
rect 7314 2535 7348 2551
rect 7314 2459 7348 2475
rect 7402 2535 7436 2551
rect 7402 2459 7436 2475
rect 7135 2408 7143 2442
rect 7101 2392 7143 2408
rect 7001 2270 7047 2390
rect 7342 2382 7358 2416
rect 7392 2382 7408 2416
rect 7081 2345 7147 2356
rect 7081 2342 7101 2345
rect 7081 2308 7097 2342
rect 7135 2311 7147 2345
rect 7131 2308 7147 2311
rect 7268 2346 7317 2358
rect 7268 2312 7277 2346
rect 7311 2341 7317 2346
rect 7311 2312 7563 2341
rect 7268 2306 7563 2312
rect 7268 2299 7317 2306
rect 7528 2283 7563 2306
rect 7001 2258 7067 2270
rect 7001 2224 7017 2258
rect 7051 2224 7067 2258
rect 7001 2190 7067 2224
rect 7001 2156 7017 2190
rect 7051 2156 7067 2190
rect 7001 2144 7067 2156
rect 7101 2258 7147 2274
rect 7528 2271 7577 2283
rect 7135 2224 7147 2258
rect 7101 2190 7147 2224
rect 7269 2253 7318 2265
rect 7269 2219 7278 2253
rect 7312 2219 7479 2253
rect 7528 2237 7537 2271
rect 7571 2237 7577 2271
rect 7528 2224 7577 2237
rect 13078 2224 13112 2240
rect 7269 2206 7318 2219
rect 7135 2156 7147 2190
rect 7101 2110 7147 2156
rect 7438 2177 7479 2219
rect 7529 2178 7578 2190
rect 7529 2177 7538 2178
rect 7438 2144 7538 2177
rect 7572 2144 7578 2178
rect 7438 2143 7578 2144
rect 7529 2131 7578 2143
rect 7963 2142 7979 2176
rect 8013 2142 8029 2176
rect 8695 2142 8711 2176
rect 8745 2142 8761 2176
rect 8821 2142 8837 2176
rect 8871 2142 8887 2176
rect 9907 2142 9923 2176
rect 9957 2142 9973 2176
rect 10033 2142 10049 2176
rect 10083 2142 10099 2176
rect 11119 2142 11135 2176
rect 11169 2142 11185 2176
rect 11245 2142 11261 2176
rect 11295 2142 11311 2176
rect 12331 2142 12347 2176
rect 12381 2142 12397 2176
rect 12457 2142 12473 2176
rect 12507 2142 12523 2176
rect 13078 2148 13112 2164
rect 13166 2224 13200 2240
rect 13166 2148 13200 2164
rect 62 2076 91 2110
rect 125 2076 183 2110
rect 217 2076 275 2110
rect 309 2076 367 2110
rect 401 2076 459 2110
rect 493 2076 522 2110
rect 1246 2083 1280 2099
rect 1246 2007 1280 2023
rect 1334 2083 1368 2099
rect 1334 2007 1368 2023
rect 1978 2083 2012 2099
rect 1978 2007 2012 2023
rect 2083 2083 2117 2099
rect 2083 2007 2117 2023
rect 2192 2083 2226 2099
rect 2192 2007 2226 2023
rect 3190 2083 3224 2099
rect 3190 2007 3224 2023
rect 3294 2083 3328 2099
rect 3294 2007 3328 2023
rect 3404 2083 3438 2099
rect 3404 2007 3438 2023
rect 4402 2083 4436 2099
rect 4402 2007 4436 2023
rect 4507 2083 4541 2099
rect 4507 2007 4541 2023
rect 4616 2083 4650 2099
rect 4616 2007 4650 2023
rect 5614 2083 5648 2099
rect 5614 2007 5648 2023
rect 5721 2083 5755 2099
rect 5721 2007 5755 2023
rect 5828 2083 5862 2099
rect 5828 2007 5862 2023
rect 6389 2086 6423 2102
rect 6389 2010 6423 2026
rect 6477 2086 6511 2102
rect 6477 2010 6511 2026
rect 6573 2086 6607 2102
rect 6573 2010 6607 2026
rect 6669 2086 6703 2102
rect 6751 2076 6780 2110
rect 6814 2076 6872 2110
rect 6906 2076 6964 2110
rect 6998 2076 7056 2110
rect 7090 2076 7148 2110
rect 7182 2076 7211 2110
rect 7935 2083 7969 2099
rect 6669 2010 6703 2026
rect 7935 2007 7969 2023
rect 8023 2083 8057 2099
rect 8023 2007 8057 2023
rect 8667 2083 8701 2099
rect 8667 2007 8701 2023
rect 8772 2083 8806 2099
rect 8772 2007 8806 2023
rect 8881 2083 8915 2099
rect 8881 2007 8915 2023
rect 9879 2083 9913 2099
rect 9879 2007 9913 2023
rect 9983 2083 10017 2099
rect 9983 2007 10017 2023
rect 10093 2083 10127 2099
rect 10093 2007 10127 2023
rect 11091 2083 11125 2099
rect 11091 2007 11125 2023
rect 11196 2083 11230 2099
rect 11196 2007 11230 2023
rect 11305 2083 11339 2099
rect 11305 2007 11339 2023
rect 12303 2083 12337 2099
rect 12303 2007 12337 2023
rect 12410 2083 12444 2099
rect 12410 2007 12444 2023
rect 12517 2083 12551 2099
rect 12517 2007 12551 2023
rect 13078 2086 13112 2102
rect 13078 2010 13112 2026
rect 13166 2086 13200 2102
rect 13166 2010 13200 2026
rect 13262 2086 13296 2102
rect 13262 2010 13296 2026
rect 13358 2086 13392 2102
rect 13358 2010 13392 2026
rect 6302 1935 6318 1969
rect 6352 1935 6368 1969
rect 6509 1933 6525 1967
rect 6559 1933 6575 1967
rect 12991 1935 13007 1969
rect 13041 1935 13057 1969
rect 13198 1933 13214 1967
rect 13248 1933 13264 1967
rect 1601 1882 1635 1898
rect 1601 1806 1635 1822
rect 1689 1882 1723 1898
rect 1689 1806 1723 1822
rect 2333 1882 2367 1898
rect 2333 1806 2367 1822
rect 2438 1882 2472 1898
rect 2438 1806 2472 1822
rect 2545 1882 2579 1898
rect 2545 1806 2579 1822
rect 3545 1882 3579 1898
rect 3545 1806 3579 1822
rect 3649 1882 3683 1898
rect 3649 1806 3683 1822
rect 3757 1882 3791 1898
rect 3757 1806 3791 1822
rect 4883 1882 4917 1898
rect 4883 1806 4917 1822
rect 4989 1882 5023 1898
rect 4989 1806 5023 1822
rect 5095 1882 5129 1898
rect 5095 1806 5129 1822
rect 5738 1882 5772 1898
rect 5738 1806 5772 1822
rect 5827 1882 5861 1898
rect 5827 1806 5861 1822
rect 6389 1883 6423 1899
rect 6389 1807 6423 1823
rect 6477 1883 6511 1899
rect 6477 1807 6511 1823
rect 6573 1883 6607 1899
rect 6573 1807 6607 1823
rect 6669 1883 6703 1899
rect 6669 1807 6703 1823
rect 8290 1882 8324 1898
rect 8290 1806 8324 1822
rect 8378 1882 8412 1898
rect 8378 1806 8412 1822
rect 9022 1882 9056 1898
rect 9022 1806 9056 1822
rect 9127 1882 9161 1898
rect 9127 1806 9161 1822
rect 9234 1882 9268 1898
rect 9234 1806 9268 1822
rect 10234 1882 10268 1898
rect 10234 1806 10268 1822
rect 10338 1882 10372 1898
rect 10338 1806 10372 1822
rect 10446 1882 10480 1898
rect 10446 1806 10480 1822
rect 11572 1882 11606 1898
rect 11572 1806 11606 1822
rect 11678 1882 11712 1898
rect 11678 1806 11712 1822
rect 11784 1882 11818 1898
rect 11784 1806 11818 1822
rect 12427 1882 12461 1898
rect 12427 1806 12461 1822
rect 12516 1882 12550 1898
rect 12516 1806 12550 1822
rect 13078 1883 13112 1899
rect 13078 1807 13112 1823
rect 13166 1883 13200 1899
rect 13166 1807 13200 1823
rect 13262 1883 13296 1899
rect 13262 1807 13296 1823
rect 13358 1883 13392 1899
rect 13358 1807 13392 1823
rect 643 1748 659 1782
rect 693 1748 709 1782
rect 1629 1738 1645 1772
rect 1679 1738 1695 1772
rect 2361 1738 2377 1772
rect 2411 1738 2427 1772
rect 2485 1738 2501 1772
rect 2535 1738 2551 1772
rect 3573 1738 3589 1772
rect 3623 1738 3639 1772
rect 3697 1738 3713 1772
rect 3747 1738 3763 1772
rect 4911 1738 4927 1772
rect 4961 1738 4977 1772
rect 5035 1738 5051 1772
rect 5085 1738 5101 1772
rect 5767 1738 5783 1772
rect 5817 1738 5833 1772
rect 6389 1745 6423 1761
rect 579 1698 613 1714
rect 579 1622 613 1638
rect 739 1698 773 1714
rect 6389 1669 6423 1685
rect 6477 1745 6511 1761
rect 7332 1748 7348 1782
rect 7382 1748 7398 1782
rect 8318 1738 8334 1772
rect 8368 1738 8384 1772
rect 9050 1738 9066 1772
rect 9100 1738 9116 1772
rect 9174 1738 9190 1772
rect 9224 1738 9240 1772
rect 10262 1738 10278 1772
rect 10312 1738 10328 1772
rect 10386 1738 10402 1772
rect 10436 1738 10452 1772
rect 11600 1738 11616 1772
rect 11650 1738 11666 1772
rect 11724 1738 11740 1772
rect 11774 1738 11790 1772
rect 12456 1738 12472 1772
rect 12506 1738 12522 1772
rect 13078 1745 13112 1761
rect 6477 1669 6511 1685
rect 7268 1698 7302 1714
rect 739 1622 773 1638
rect 7268 1622 7302 1638
rect 7428 1698 7462 1714
rect 13078 1669 13112 1685
rect 13166 1745 13200 1761
rect 13166 1669 13200 1685
rect 7428 1622 7462 1638
rect 579 1560 613 1576
rect 579 1484 613 1500
rect 739 1560 773 1576
rect 739 1484 773 1500
rect 7268 1560 7302 1576
rect 7268 1484 7302 1500
rect 7428 1560 7462 1576
rect 7428 1484 7462 1500
rect 579 1422 613 1438
rect 579 1346 613 1362
rect 739 1422 773 1438
rect 739 1346 773 1362
rect 7268 1422 7302 1438
rect 7268 1346 7302 1362
rect 7428 1422 7462 1438
rect 7428 1346 7462 1362
rect 579 1284 613 1300
rect 579 1208 613 1224
rect 739 1284 773 1300
rect 739 1208 773 1224
rect 7268 1284 7302 1300
rect 7268 1208 7302 1224
rect 7428 1284 7462 1300
rect 7428 1208 7462 1224
rect 579 1146 613 1162
rect 579 1070 613 1086
rect 739 1146 773 1162
rect 739 1070 773 1086
rect 7268 1146 7302 1162
rect 7268 1070 7302 1086
rect 7428 1146 7462 1162
rect 7428 1070 7462 1086
rect 579 1008 613 1024
rect 579 932 613 948
rect 739 1008 773 1024
rect 739 932 773 948
rect 7268 1008 7302 1024
rect 7268 932 7302 948
rect 7428 1008 7462 1024
rect 7428 932 7462 948
rect 579 870 613 886
rect 579 794 613 810
rect 739 870 773 886
rect 739 794 773 810
rect 7268 870 7302 886
rect 7268 794 7302 810
rect 7428 870 7462 886
rect 7428 794 7462 810
rect 579 732 613 748
rect 579 656 613 672
rect 739 732 773 748
rect 739 656 773 672
rect 7268 732 7302 748
rect 7268 656 7302 672
rect 7428 732 7462 748
rect 7428 656 7462 672
rect 6076 276 6110 292
rect 6076 200 6110 216
rect 6236 276 6270 292
rect 6236 200 6270 216
rect 12831 276 12865 292
rect 12831 200 12865 216
rect 12991 276 13025 292
rect 12991 200 13025 216
rect 6076 138 6110 154
rect 6076 62 6110 78
rect 6236 138 6270 154
rect 6236 62 6270 78
rect 12831 138 12865 154
rect 12831 62 12865 78
rect 12991 138 13025 154
rect 12991 62 13025 78
rect 6076 0 6110 16
rect 6076 -76 6110 -60
rect 6236 0 6270 16
rect 6236 -76 6270 -60
rect 12831 0 12865 16
rect 12831 -76 12865 -60
rect 12991 0 13025 16
rect 12991 -76 13025 -60
rect 6076 -138 6110 -122
rect 6076 -214 6110 -198
rect 6236 -138 6270 -122
rect 6236 -214 6270 -198
rect 12831 -138 12865 -122
rect 12831 -214 12865 -198
rect 12991 -138 13025 -122
rect 12991 -214 13025 -198
rect 6076 -276 6110 -260
rect 6076 -352 6110 -336
rect 6236 -276 6270 -260
rect 6236 -352 6270 -336
rect 12831 -276 12865 -260
rect 12831 -352 12865 -336
rect 12991 -276 13025 -260
rect 12991 -352 13025 -336
rect 6076 -414 6110 -398
rect 6076 -490 6110 -474
rect 6236 -414 6270 -398
rect 6236 -490 6270 -474
rect 12831 -414 12865 -398
rect 12831 -490 12865 -474
rect 12991 -414 13025 -398
rect 12991 -490 13025 -474
rect 6076 -552 6110 -536
rect 6076 -628 6110 -612
rect 6236 -552 6270 -536
rect 6236 -628 6270 -612
rect 12831 -552 12865 -536
rect 12831 -628 12865 -612
rect 12991 -552 13025 -536
rect 12991 -628 13025 -612
rect 6076 -690 6110 -674
rect 338 -737 372 -721
rect 338 -813 372 -797
rect 426 -737 460 -721
rect 6076 -766 6110 -750
rect 6236 -690 6270 -674
rect 12831 -690 12865 -674
rect 6236 -766 6270 -750
rect 7093 -737 7127 -721
rect 426 -813 460 -797
rect 1016 -824 1032 -790
rect 1066 -824 1082 -790
rect 1748 -824 1764 -790
rect 1798 -824 1814 -790
rect 1872 -824 1888 -790
rect 1922 -824 1938 -790
rect 3086 -824 3102 -790
rect 3136 -824 3152 -790
rect 3210 -824 3226 -790
rect 3260 -824 3276 -790
rect 4298 -824 4314 -790
rect 4348 -824 4364 -790
rect 4422 -824 4438 -790
rect 4472 -824 4488 -790
rect 5154 -824 5170 -790
rect 5204 -824 5220 -790
rect 6140 -834 6156 -800
rect 6190 -834 6206 -800
rect 7093 -813 7127 -797
rect 7181 -737 7215 -721
rect 12831 -766 12865 -750
rect 12991 -690 13025 -674
rect 12991 -766 13025 -750
rect 7181 -813 7215 -797
rect 7771 -824 7787 -790
rect 7821 -824 7837 -790
rect 8503 -824 8519 -790
rect 8553 -824 8569 -790
rect 8627 -824 8643 -790
rect 8677 -824 8693 -790
rect 9841 -824 9857 -790
rect 9891 -824 9907 -790
rect 9965 -824 9981 -790
rect 10015 -824 10031 -790
rect 11053 -824 11069 -790
rect 11103 -824 11119 -790
rect 11177 -824 11193 -790
rect 11227 -824 11243 -790
rect 11909 -824 11925 -790
rect 11959 -824 11975 -790
rect 12895 -834 12911 -800
rect 12945 -834 12961 -800
rect 146 -875 180 -859
rect 146 -951 180 -935
rect 242 -875 276 -859
rect 242 -951 276 -935
rect 338 -875 372 -859
rect 338 -951 372 -935
rect 426 -875 460 -859
rect 426 -951 460 -935
rect 988 -874 1022 -858
rect 988 -950 1022 -934
rect 1077 -874 1111 -858
rect 1077 -950 1111 -934
rect 1720 -874 1754 -858
rect 1720 -950 1754 -934
rect 1826 -874 1860 -858
rect 1826 -950 1860 -934
rect 1932 -874 1966 -858
rect 1932 -950 1966 -934
rect 3058 -874 3092 -858
rect 3058 -950 3092 -934
rect 3166 -874 3200 -858
rect 3166 -950 3200 -934
rect 3270 -874 3304 -858
rect 3270 -950 3304 -934
rect 4270 -874 4304 -858
rect 4270 -950 4304 -934
rect 4377 -874 4411 -858
rect 4377 -950 4411 -934
rect 4482 -874 4516 -858
rect 4482 -950 4516 -934
rect 5126 -874 5160 -858
rect 5126 -950 5160 -934
rect 5214 -874 5248 -858
rect 5214 -950 5248 -934
rect 6901 -875 6935 -859
rect 6901 -951 6935 -935
rect 6997 -875 7031 -859
rect 6997 -951 7031 -935
rect 7093 -875 7127 -859
rect 7093 -951 7127 -935
rect 7181 -875 7215 -859
rect 7181 -951 7215 -935
rect 7743 -874 7777 -858
rect 7743 -950 7777 -934
rect 7832 -874 7866 -858
rect 7832 -950 7866 -934
rect 8475 -874 8509 -858
rect 8475 -950 8509 -934
rect 8581 -874 8615 -858
rect 8581 -950 8615 -934
rect 8687 -874 8721 -858
rect 8687 -950 8721 -934
rect 9813 -874 9847 -858
rect 9813 -950 9847 -934
rect 9921 -874 9955 -858
rect 9921 -950 9955 -934
rect 10025 -874 10059 -858
rect 10025 -950 10059 -934
rect 11025 -874 11059 -858
rect 11025 -950 11059 -934
rect 11132 -874 11166 -858
rect 11132 -950 11166 -934
rect 11237 -874 11271 -858
rect 11237 -950 11271 -934
rect 11881 -874 11915 -858
rect 11881 -950 11915 -934
rect 11969 -874 12003 -858
rect 11969 -950 12003 -934
rect 274 -1019 290 -985
rect 324 -1019 340 -985
rect 481 -1021 497 -987
rect 531 -1021 547 -987
rect 7029 -1019 7045 -985
rect 7079 -1019 7095 -985
rect 7236 -1021 7252 -987
rect 7286 -1021 7302 -987
rect 146 -1078 180 -1062
rect 146 -1154 180 -1138
rect 242 -1078 276 -1062
rect 242 -1154 276 -1138
rect 338 -1078 372 -1062
rect 338 -1154 372 -1138
rect 426 -1078 460 -1062
rect 426 -1154 460 -1138
rect 987 -1075 1021 -1059
rect 987 -1151 1021 -1135
rect 1094 -1075 1128 -1059
rect 1094 -1151 1128 -1135
rect 1201 -1075 1235 -1059
rect 1201 -1151 1235 -1135
rect 2199 -1075 2233 -1059
rect 2199 -1151 2233 -1135
rect 2308 -1075 2342 -1059
rect 2308 -1151 2342 -1135
rect 2413 -1075 2447 -1059
rect 2413 -1151 2447 -1135
rect 3411 -1075 3445 -1059
rect 3411 -1151 3445 -1135
rect 3521 -1075 3555 -1059
rect 3521 -1151 3555 -1135
rect 3625 -1075 3659 -1059
rect 3625 -1151 3659 -1135
rect 4623 -1075 4657 -1059
rect 4623 -1151 4657 -1135
rect 4732 -1075 4766 -1059
rect 4732 -1151 4766 -1135
rect 4837 -1075 4871 -1059
rect 4837 -1151 4871 -1135
rect 5481 -1075 5515 -1059
rect 5481 -1151 5515 -1135
rect 5569 -1075 5603 -1059
rect 6901 -1078 6935 -1062
rect 5569 -1151 5603 -1135
rect 6327 -1162 6356 -1128
rect 6390 -1162 6448 -1128
rect 6482 -1162 6540 -1128
rect 6574 -1162 6632 -1128
rect 6666 -1162 6724 -1128
rect 6758 -1162 6787 -1128
rect 6901 -1154 6935 -1138
rect 6997 -1078 7031 -1062
rect 6997 -1154 7031 -1138
rect 7093 -1078 7127 -1062
rect 7093 -1154 7127 -1138
rect 7181 -1078 7215 -1062
rect 7181 -1154 7215 -1138
rect 7742 -1075 7776 -1059
rect 7742 -1151 7776 -1135
rect 7849 -1075 7883 -1059
rect 7849 -1151 7883 -1135
rect 7956 -1075 7990 -1059
rect 7956 -1151 7990 -1135
rect 8954 -1075 8988 -1059
rect 8954 -1151 8988 -1135
rect 9063 -1075 9097 -1059
rect 9063 -1151 9097 -1135
rect 9168 -1075 9202 -1059
rect 9168 -1151 9202 -1135
rect 10166 -1075 10200 -1059
rect 10166 -1151 10200 -1135
rect 10276 -1075 10310 -1059
rect 10276 -1151 10310 -1135
rect 10380 -1075 10414 -1059
rect 10380 -1151 10414 -1135
rect 11378 -1075 11412 -1059
rect 11378 -1151 11412 -1135
rect 11487 -1075 11521 -1059
rect 11487 -1151 11521 -1135
rect 11592 -1075 11626 -1059
rect 11592 -1151 11626 -1135
rect 12236 -1075 12270 -1059
rect 12236 -1151 12270 -1135
rect 12324 -1075 12358 -1059
rect 12324 -1151 12358 -1135
rect 13082 -1162 13111 -1128
rect 13145 -1162 13203 -1128
rect 13237 -1162 13295 -1128
rect 13329 -1162 13387 -1128
rect 13421 -1162 13479 -1128
rect 13513 -1162 13542 -1128
rect 338 -1216 372 -1200
rect 338 -1292 372 -1276
rect 426 -1216 460 -1200
rect 1015 -1228 1031 -1194
rect 1065 -1228 1081 -1194
rect 1141 -1228 1157 -1194
rect 1191 -1228 1207 -1194
rect 2227 -1228 2243 -1194
rect 2277 -1228 2293 -1194
rect 2353 -1228 2369 -1194
rect 2403 -1228 2419 -1194
rect 3439 -1228 3455 -1194
rect 3489 -1228 3505 -1194
rect 3565 -1228 3581 -1194
rect 3615 -1228 3631 -1194
rect 4651 -1228 4667 -1194
rect 4701 -1228 4717 -1194
rect 4777 -1228 4793 -1194
rect 4827 -1228 4843 -1194
rect 5509 -1228 5525 -1194
rect 5559 -1228 5575 -1194
rect 5960 -1195 6009 -1183
rect 5960 -1196 6100 -1195
rect 5960 -1230 5966 -1196
rect 6000 -1229 6100 -1196
rect 6000 -1230 6009 -1229
rect 5960 -1242 6009 -1230
rect 6059 -1271 6100 -1229
rect 6391 -1208 6437 -1162
rect 6391 -1242 6403 -1208
rect 6220 -1271 6269 -1258
rect 426 -1292 460 -1276
rect 5961 -1289 6010 -1276
rect 5961 -1323 5967 -1289
rect 6001 -1323 6010 -1289
rect 6059 -1305 6226 -1271
rect 6260 -1305 6269 -1271
rect 6220 -1317 6269 -1305
rect 6391 -1276 6437 -1242
rect 6391 -1310 6403 -1276
rect 5961 -1335 6010 -1323
rect 6391 -1326 6437 -1310
rect 6471 -1208 6537 -1196
rect 6471 -1242 6487 -1208
rect 6521 -1242 6537 -1208
rect 6471 -1276 6537 -1242
rect 6471 -1310 6487 -1276
rect 6521 -1310 6537 -1276
rect 6471 -1322 6537 -1310
rect 5975 -1358 6010 -1335
rect 6221 -1358 6270 -1351
rect 5975 -1364 6270 -1358
rect 5975 -1393 6227 -1364
rect 6221 -1398 6227 -1393
rect 6261 -1398 6270 -1364
rect 6221 -1410 6270 -1398
rect 6391 -1363 6407 -1360
rect 6391 -1397 6403 -1363
rect 6441 -1394 6457 -1360
rect 6437 -1397 6457 -1394
rect 6391 -1408 6457 -1397
rect 6130 -1468 6146 -1434
rect 6180 -1468 6196 -1434
rect 6491 -1442 6537 -1322
rect 6395 -1460 6437 -1444
rect 6395 -1494 6403 -1460
rect 6102 -1527 6136 -1511
rect 6102 -1603 6136 -1587
rect 6190 -1527 6224 -1511
rect 6190 -1603 6224 -1587
rect 6395 -1528 6437 -1494
rect 6395 -1562 6403 -1528
rect 6395 -1596 6437 -1562
rect 6395 -1630 6403 -1596
rect 6102 -1665 6136 -1649
rect 6102 -1741 6136 -1725
rect 6190 -1665 6224 -1649
rect 6395 -1672 6437 -1630
rect 6471 -1460 6537 -1442
rect 6471 -1508 6487 -1460
rect 6521 -1508 6537 -1460
rect 6471 -1528 6537 -1508
rect 6471 -1562 6487 -1528
rect 6521 -1562 6537 -1528
rect 6471 -1596 6537 -1562
rect 6471 -1630 6487 -1596
rect 6521 -1630 6537 -1596
rect 6471 -1638 6537 -1630
rect 6577 -1208 6643 -1196
rect 6577 -1242 6593 -1208
rect 6627 -1242 6643 -1208
rect 6577 -1276 6643 -1242
rect 6577 -1310 6593 -1276
rect 6627 -1310 6643 -1276
rect 6577 -1322 6643 -1310
rect 6677 -1208 6723 -1162
rect 6711 -1242 6723 -1208
rect 6677 -1276 6723 -1242
rect 6711 -1310 6723 -1276
rect 7093 -1216 7127 -1200
rect 7093 -1292 7127 -1276
rect 7181 -1216 7215 -1200
rect 7770 -1228 7786 -1194
rect 7820 -1228 7836 -1194
rect 7896 -1228 7912 -1194
rect 7946 -1228 7962 -1194
rect 8982 -1228 8998 -1194
rect 9032 -1228 9048 -1194
rect 9108 -1228 9124 -1194
rect 9158 -1228 9174 -1194
rect 10194 -1228 10210 -1194
rect 10244 -1228 10260 -1194
rect 10320 -1228 10336 -1194
rect 10370 -1228 10386 -1194
rect 11406 -1228 11422 -1194
rect 11456 -1228 11472 -1194
rect 11532 -1228 11548 -1194
rect 11582 -1228 11598 -1194
rect 12264 -1228 12280 -1194
rect 12314 -1228 12330 -1194
rect 12715 -1195 12764 -1183
rect 12715 -1196 12855 -1195
rect 12715 -1230 12721 -1196
rect 12755 -1229 12855 -1196
rect 12755 -1230 12764 -1229
rect 12715 -1242 12764 -1230
rect 12814 -1271 12855 -1229
rect 13146 -1208 13192 -1162
rect 13146 -1242 13158 -1208
rect 12975 -1271 13024 -1258
rect 7181 -1292 7215 -1276
rect 12716 -1289 12765 -1276
rect 6577 -1442 6623 -1322
rect 6677 -1326 6723 -1310
rect 12716 -1323 12722 -1289
rect 12756 -1323 12765 -1289
rect 12814 -1305 12981 -1271
rect 13015 -1305 13024 -1271
rect 12975 -1317 13024 -1305
rect 13146 -1276 13192 -1242
rect 13146 -1310 13158 -1276
rect 12716 -1335 12765 -1323
rect 13146 -1326 13192 -1310
rect 13226 -1208 13292 -1196
rect 13226 -1242 13242 -1208
rect 13276 -1242 13292 -1208
rect 13226 -1276 13292 -1242
rect 13226 -1310 13242 -1276
rect 13276 -1310 13292 -1276
rect 13226 -1322 13292 -1310
rect 12730 -1358 12765 -1335
rect 12976 -1358 13025 -1351
rect 6657 -1394 6673 -1360
rect 6707 -1364 6723 -1360
rect 6657 -1398 6677 -1394
rect 6711 -1398 6723 -1364
rect 12730 -1364 13025 -1358
rect 12730 -1393 12982 -1364
rect 6657 -1408 6723 -1398
rect 12976 -1398 12982 -1393
rect 13016 -1398 13025 -1364
rect 12976 -1410 13025 -1398
rect 13146 -1363 13162 -1360
rect 13146 -1397 13158 -1363
rect 13196 -1394 13212 -1360
rect 13192 -1397 13212 -1394
rect 13146 -1408 13212 -1397
rect 6577 -1460 6643 -1442
rect 6577 -1494 6593 -1460
rect 6627 -1494 6643 -1460
rect 6577 -1528 6643 -1494
rect 6577 -1562 6593 -1528
rect 6627 -1529 6643 -1528
rect 6577 -1563 6596 -1562
rect 6630 -1563 6643 -1529
rect 6577 -1596 6643 -1563
rect 6577 -1630 6593 -1596
rect 6627 -1630 6643 -1596
rect 6577 -1638 6643 -1630
rect 6677 -1460 6719 -1444
rect 6711 -1494 6719 -1460
rect 12885 -1468 12901 -1434
rect 12935 -1468 12951 -1434
rect 13246 -1442 13292 -1322
rect 13150 -1460 13192 -1444
rect 6677 -1528 6719 -1494
rect 13150 -1494 13158 -1460
rect 6711 -1562 6719 -1528
rect 6677 -1596 6719 -1562
rect 6711 -1630 6719 -1596
rect 12857 -1527 12891 -1511
rect 12857 -1603 12891 -1587
rect 12945 -1527 12979 -1511
rect 12945 -1603 12979 -1587
rect 13150 -1528 13192 -1494
rect 13150 -1562 13158 -1528
rect 13150 -1596 13192 -1562
rect 6677 -1672 6719 -1630
rect 13150 -1630 13158 -1596
rect 12857 -1665 12891 -1649
rect 6327 -1706 6356 -1672
rect 6390 -1706 6448 -1672
rect 6482 -1706 6540 -1672
rect 6574 -1706 6632 -1672
rect 6666 -1706 6724 -1672
rect 6758 -1706 6787 -1672
rect 6190 -1741 6224 -1725
rect 12857 -1741 12891 -1725
rect 12945 -1665 12979 -1649
rect 13150 -1672 13192 -1630
rect 13226 -1460 13292 -1442
rect 13226 -1508 13242 -1460
rect 13276 -1508 13292 -1460
rect 13226 -1528 13292 -1508
rect 13226 -1562 13242 -1528
rect 13276 -1562 13292 -1528
rect 13226 -1596 13292 -1562
rect 13226 -1630 13242 -1596
rect 13276 -1630 13292 -1596
rect 13226 -1638 13292 -1630
rect 13332 -1208 13398 -1196
rect 13332 -1242 13348 -1208
rect 13382 -1242 13398 -1208
rect 13332 -1276 13398 -1242
rect 13332 -1310 13348 -1276
rect 13382 -1310 13398 -1276
rect 13332 -1322 13398 -1310
rect 13432 -1208 13478 -1162
rect 13466 -1242 13478 -1208
rect 13432 -1276 13478 -1242
rect 13466 -1310 13478 -1276
rect 13332 -1442 13378 -1322
rect 13432 -1326 13478 -1310
rect 13412 -1394 13428 -1360
rect 13462 -1364 13478 -1360
rect 13412 -1398 13432 -1394
rect 13466 -1398 13478 -1364
rect 13412 -1408 13478 -1398
rect 13332 -1460 13398 -1442
rect 13332 -1494 13348 -1460
rect 13382 -1494 13398 -1460
rect 13332 -1528 13398 -1494
rect 13332 -1562 13348 -1528
rect 13382 -1529 13398 -1528
rect 13332 -1563 13351 -1562
rect 13385 -1563 13398 -1529
rect 13332 -1596 13398 -1563
rect 13332 -1630 13348 -1596
rect 13382 -1630 13398 -1596
rect 13332 -1638 13398 -1630
rect 13432 -1460 13474 -1444
rect 13466 -1494 13474 -1460
rect 13432 -1528 13474 -1494
rect 13466 -1562 13474 -1528
rect 13432 -1596 13474 -1562
rect 13466 -1630 13474 -1596
rect 13432 -1672 13474 -1630
rect 13082 -1706 13111 -1672
rect 13145 -1706 13203 -1672
rect 13237 -1706 13295 -1672
rect 13329 -1706 13387 -1672
rect 13421 -1706 13479 -1672
rect 13513 -1706 13542 -1672
rect 12945 -1741 12979 -1725
rect 6102 -1803 6136 -1787
rect 6102 -1879 6136 -1863
rect 6190 -1803 6224 -1787
rect 6190 -1879 6224 -1863
rect 12857 -1803 12891 -1787
rect 12857 -1879 12891 -1863
rect 12945 -1803 12979 -1787
rect 12945 -1879 12979 -1863
rect 6102 -1941 6136 -1925
rect 6102 -2017 6136 -2001
rect 6190 -1941 6224 -1925
rect 6190 -2017 6224 -2001
rect 12857 -1941 12891 -1925
rect 12857 -2017 12891 -2001
rect 12945 -1941 12979 -1925
rect 12945 -2017 12979 -2001
rect 6102 -2079 6136 -2063
rect 6102 -2155 6136 -2139
rect 6190 -2079 6224 -2063
rect 6190 -2155 6224 -2139
rect 12857 -2079 12891 -2063
rect 12857 -2155 12891 -2139
rect 12945 -2079 12979 -2063
rect 12945 -2155 12979 -2139
rect 6102 -2217 6136 -2201
rect 6102 -2293 6136 -2277
rect 6190 -2217 6224 -2201
rect 6190 -2293 6224 -2277
rect 12857 -2217 12891 -2201
rect 12857 -2293 12891 -2277
rect 12945 -2217 12979 -2201
rect 12945 -2293 12979 -2277
<< viali >>
rect 625 3165 659 3225
rect 713 3165 747 3225
rect 7314 3165 7348 3225
rect 7402 3165 7436 3225
rect 625 3027 659 3087
rect 713 3027 747 3087
rect 7314 3027 7348 3087
rect 7402 3027 7436 3087
rect 625 2889 659 2949
rect 713 2889 747 2949
rect 7314 2889 7348 2949
rect 7402 2889 7436 2949
rect 625 2751 659 2811
rect 713 2751 747 2811
rect 7314 2751 7348 2811
rect 7402 2751 7436 2811
rect 91 2620 125 2654
rect 183 2620 217 2654
rect 275 2620 309 2654
rect 367 2620 401 2654
rect 459 2620 493 2654
rect 219 2510 253 2511
rect 219 2477 222 2510
rect 222 2477 253 2510
rect 138 2342 172 2346
rect 138 2312 142 2342
rect 142 2312 172 2342
rect 328 2442 362 2456
rect 328 2422 362 2442
rect 625 2613 659 2673
rect 713 2613 747 2673
rect 6780 2620 6814 2654
rect 6872 2620 6906 2654
rect 6964 2620 6998 2654
rect 7056 2620 7090 2654
rect 7148 2620 7182 2654
rect 625 2475 659 2535
rect 713 2475 747 2535
rect 669 2382 703 2416
rect 6908 2510 6942 2511
rect 6908 2477 6911 2510
rect 6911 2477 6942 2510
rect 412 2342 446 2345
rect 412 2311 442 2342
rect 442 2311 446 2342
rect 588 2312 622 2346
rect 6827 2342 6861 2346
rect 6827 2312 6831 2342
rect 6831 2312 6861 2342
rect 589 2219 623 2253
rect 848 2237 882 2271
rect 849 2144 883 2178
rect 1290 2142 1324 2176
rect 2022 2142 2056 2176
rect 2148 2142 2182 2176
rect 3234 2142 3268 2176
rect 3360 2142 3394 2176
rect 4446 2142 4480 2176
rect 4572 2142 4606 2176
rect 5658 2142 5692 2176
rect 5784 2142 5818 2176
rect 6389 2164 6423 2224
rect 6477 2164 6511 2224
rect 7017 2442 7051 2456
rect 7017 2422 7051 2442
rect 7314 2613 7348 2673
rect 7402 2613 7436 2673
rect 7314 2475 7348 2535
rect 7402 2475 7436 2535
rect 7358 2382 7392 2416
rect 7101 2342 7135 2345
rect 7101 2311 7131 2342
rect 7131 2311 7135 2342
rect 7277 2312 7311 2346
rect 7278 2219 7312 2253
rect 7537 2237 7571 2271
rect 7538 2144 7572 2178
rect 7979 2142 8013 2176
rect 8711 2142 8745 2176
rect 8837 2142 8871 2176
rect 9923 2142 9957 2176
rect 10049 2142 10083 2176
rect 11135 2142 11169 2176
rect 11261 2142 11295 2176
rect 12347 2142 12381 2176
rect 12473 2142 12507 2176
rect 13078 2164 13112 2224
rect 13166 2164 13200 2224
rect 91 2076 125 2110
rect 183 2076 217 2110
rect 275 2076 309 2110
rect 367 2076 401 2110
rect 459 2076 493 2110
rect 1246 2023 1280 2083
rect 1334 2023 1368 2083
rect 1978 2023 2012 2083
rect 2083 2023 2117 2083
rect 2192 2023 2226 2083
rect 3190 2023 3224 2083
rect 3294 2023 3328 2083
rect 3404 2023 3438 2083
rect 4402 2023 4436 2083
rect 4507 2023 4541 2083
rect 4616 2023 4650 2083
rect 5614 2023 5648 2083
rect 5721 2023 5755 2083
rect 5828 2023 5862 2083
rect 6389 2026 6423 2086
rect 6477 2026 6511 2086
rect 6573 2026 6607 2086
rect 6669 2026 6703 2086
rect 6780 2076 6814 2110
rect 6872 2076 6906 2110
rect 6964 2076 6998 2110
rect 7056 2076 7090 2110
rect 7148 2076 7182 2110
rect 7935 2023 7969 2083
rect 8023 2023 8057 2083
rect 8667 2023 8701 2083
rect 8772 2023 8806 2083
rect 8881 2023 8915 2083
rect 9879 2023 9913 2083
rect 9983 2023 10017 2083
rect 10093 2023 10127 2083
rect 11091 2023 11125 2083
rect 11196 2023 11230 2083
rect 11305 2023 11339 2083
rect 12303 2023 12337 2083
rect 12410 2023 12444 2083
rect 12517 2023 12551 2083
rect 13078 2026 13112 2086
rect 13166 2026 13200 2086
rect 13262 2026 13296 2086
rect 13358 2026 13392 2086
rect 6318 1935 6352 1969
rect 6525 1933 6559 1967
rect 13007 1935 13041 1969
rect 13214 1933 13248 1967
rect 1601 1822 1635 1882
rect 1689 1822 1723 1882
rect 2333 1822 2367 1882
rect 2438 1822 2472 1882
rect 2545 1822 2579 1882
rect 3545 1822 3579 1882
rect 3649 1822 3683 1882
rect 3757 1822 3791 1882
rect 4883 1822 4917 1882
rect 4989 1822 5023 1882
rect 5095 1822 5129 1882
rect 5738 1822 5772 1882
rect 5827 1822 5861 1882
rect 6389 1823 6423 1883
rect 6477 1823 6511 1883
rect 6573 1823 6607 1883
rect 6669 1823 6703 1883
rect 8290 1822 8324 1882
rect 8378 1822 8412 1882
rect 9022 1822 9056 1882
rect 9127 1822 9161 1882
rect 9234 1822 9268 1882
rect 10234 1822 10268 1882
rect 10338 1822 10372 1882
rect 10446 1822 10480 1882
rect 11572 1822 11606 1882
rect 11678 1822 11712 1882
rect 11784 1822 11818 1882
rect 12427 1822 12461 1882
rect 12516 1822 12550 1882
rect 13078 1823 13112 1883
rect 13166 1823 13200 1883
rect 13262 1823 13296 1883
rect 13358 1823 13392 1883
rect 659 1748 693 1782
rect 1645 1738 1679 1772
rect 2377 1738 2411 1772
rect 2501 1738 2535 1772
rect 3589 1738 3623 1772
rect 3713 1738 3747 1772
rect 4927 1738 4961 1772
rect 5051 1738 5085 1772
rect 5783 1738 5817 1772
rect 579 1638 613 1698
rect 739 1638 773 1698
rect 6389 1685 6423 1745
rect 7348 1748 7382 1782
rect 6477 1685 6511 1745
rect 8334 1738 8368 1772
rect 9066 1738 9100 1772
rect 9190 1738 9224 1772
rect 10278 1738 10312 1772
rect 10402 1738 10436 1772
rect 11616 1738 11650 1772
rect 11740 1738 11774 1772
rect 12472 1738 12506 1772
rect 7268 1638 7302 1698
rect 7428 1638 7462 1698
rect 13078 1685 13112 1745
rect 13166 1685 13200 1745
rect 579 1500 613 1560
rect 739 1500 773 1560
rect 7268 1500 7302 1560
rect 7428 1500 7462 1560
rect 579 1362 613 1422
rect 739 1362 773 1422
rect 7268 1362 7302 1422
rect 7428 1362 7462 1422
rect 579 1224 613 1284
rect 739 1224 773 1284
rect 7268 1224 7302 1284
rect 7428 1224 7462 1284
rect 579 1086 613 1146
rect 739 1086 773 1146
rect 7268 1086 7302 1146
rect 7428 1086 7462 1146
rect 579 948 613 1008
rect 739 948 773 1008
rect 7268 948 7302 1008
rect 7428 948 7462 1008
rect 579 810 613 870
rect 739 810 773 870
rect 7268 810 7302 870
rect 7428 810 7462 870
rect 579 672 613 732
rect 739 672 773 732
rect 7268 672 7302 732
rect 7428 672 7462 732
rect 6076 216 6110 276
rect 6236 216 6270 276
rect 12831 216 12865 276
rect 12991 216 13025 276
rect 6076 78 6110 138
rect 6236 78 6270 138
rect 12831 78 12865 138
rect 12991 78 13025 138
rect 6076 -60 6110 0
rect 6236 -60 6270 0
rect 12831 -60 12865 0
rect 12991 -60 13025 0
rect 6076 -198 6110 -138
rect 6236 -198 6270 -138
rect 12831 -198 12865 -138
rect 12991 -198 13025 -138
rect 6076 -336 6110 -276
rect 6236 -336 6270 -276
rect 12831 -336 12865 -276
rect 12991 -336 13025 -276
rect 6076 -474 6110 -414
rect 6236 -474 6270 -414
rect 12831 -474 12865 -414
rect 12991 -474 13025 -414
rect 6076 -612 6110 -552
rect 6236 -612 6270 -552
rect 12831 -612 12865 -552
rect 12991 -612 13025 -552
rect 338 -797 372 -737
rect 426 -797 460 -737
rect 6076 -750 6110 -690
rect 6236 -750 6270 -690
rect 1032 -824 1066 -790
rect 1764 -824 1798 -790
rect 1888 -824 1922 -790
rect 3102 -824 3136 -790
rect 3226 -824 3260 -790
rect 4314 -824 4348 -790
rect 4438 -824 4472 -790
rect 5170 -824 5204 -790
rect 7093 -797 7127 -737
rect 6156 -834 6190 -800
rect 7181 -797 7215 -737
rect 12831 -750 12865 -690
rect 12991 -750 13025 -690
rect 7787 -824 7821 -790
rect 8519 -824 8553 -790
rect 8643 -824 8677 -790
rect 9857 -824 9891 -790
rect 9981 -824 10015 -790
rect 11069 -824 11103 -790
rect 11193 -824 11227 -790
rect 11925 -824 11959 -790
rect 12911 -834 12945 -800
rect 146 -935 180 -875
rect 242 -935 276 -875
rect 338 -935 372 -875
rect 426 -935 460 -875
rect 988 -934 1022 -874
rect 1077 -934 1111 -874
rect 1720 -934 1754 -874
rect 1826 -934 1860 -874
rect 1932 -934 1966 -874
rect 3058 -934 3092 -874
rect 3166 -934 3200 -874
rect 3270 -934 3304 -874
rect 4270 -934 4304 -874
rect 4377 -934 4411 -874
rect 4482 -934 4516 -874
rect 5126 -934 5160 -874
rect 5214 -934 5248 -874
rect 6901 -935 6935 -875
rect 6997 -935 7031 -875
rect 7093 -935 7127 -875
rect 7181 -935 7215 -875
rect 7743 -934 7777 -874
rect 7832 -934 7866 -874
rect 8475 -934 8509 -874
rect 8581 -934 8615 -874
rect 8687 -934 8721 -874
rect 9813 -934 9847 -874
rect 9921 -934 9955 -874
rect 10025 -934 10059 -874
rect 11025 -934 11059 -874
rect 11132 -934 11166 -874
rect 11237 -934 11271 -874
rect 11881 -934 11915 -874
rect 11969 -934 12003 -874
rect 290 -1019 324 -985
rect 497 -1021 531 -987
rect 7045 -1019 7079 -985
rect 7252 -1021 7286 -987
rect 146 -1138 180 -1078
rect 242 -1138 276 -1078
rect 338 -1138 372 -1078
rect 426 -1138 460 -1078
rect 987 -1135 1021 -1075
rect 1094 -1135 1128 -1075
rect 1201 -1135 1235 -1075
rect 2199 -1135 2233 -1075
rect 2308 -1135 2342 -1075
rect 2413 -1135 2447 -1075
rect 3411 -1135 3445 -1075
rect 3521 -1135 3555 -1075
rect 3625 -1135 3659 -1075
rect 4623 -1135 4657 -1075
rect 4732 -1135 4766 -1075
rect 4837 -1135 4871 -1075
rect 5481 -1135 5515 -1075
rect 5569 -1135 5603 -1075
rect 6356 -1162 6390 -1128
rect 6448 -1162 6482 -1128
rect 6540 -1162 6574 -1128
rect 6632 -1162 6666 -1128
rect 6724 -1162 6758 -1128
rect 6901 -1138 6935 -1078
rect 6997 -1138 7031 -1078
rect 7093 -1138 7127 -1078
rect 7181 -1138 7215 -1078
rect 7742 -1135 7776 -1075
rect 7849 -1135 7883 -1075
rect 7956 -1135 7990 -1075
rect 8954 -1135 8988 -1075
rect 9063 -1135 9097 -1075
rect 9168 -1135 9202 -1075
rect 10166 -1135 10200 -1075
rect 10276 -1135 10310 -1075
rect 10380 -1135 10414 -1075
rect 11378 -1135 11412 -1075
rect 11487 -1135 11521 -1075
rect 11592 -1135 11626 -1075
rect 12236 -1135 12270 -1075
rect 12324 -1135 12358 -1075
rect 13111 -1162 13145 -1128
rect 13203 -1162 13237 -1128
rect 13295 -1162 13329 -1128
rect 13387 -1162 13421 -1128
rect 13479 -1162 13513 -1128
rect 338 -1276 372 -1216
rect 426 -1276 460 -1216
rect 1031 -1228 1065 -1194
rect 1157 -1228 1191 -1194
rect 2243 -1228 2277 -1194
rect 2369 -1228 2403 -1194
rect 3455 -1228 3489 -1194
rect 3581 -1228 3615 -1194
rect 4667 -1228 4701 -1194
rect 4793 -1228 4827 -1194
rect 5525 -1228 5559 -1194
rect 5966 -1230 6000 -1196
rect 5967 -1323 6001 -1289
rect 6226 -1305 6260 -1271
rect 6227 -1398 6261 -1364
rect 6403 -1394 6407 -1363
rect 6407 -1394 6437 -1363
rect 6403 -1397 6437 -1394
rect 6146 -1468 6180 -1434
rect 6102 -1587 6136 -1527
rect 6190 -1587 6224 -1527
rect 6102 -1725 6136 -1665
rect 6190 -1725 6224 -1665
rect 6487 -1494 6521 -1474
rect 6487 -1508 6521 -1494
rect 7093 -1276 7127 -1216
rect 7181 -1276 7215 -1216
rect 7786 -1228 7820 -1194
rect 7912 -1228 7946 -1194
rect 8998 -1228 9032 -1194
rect 9124 -1228 9158 -1194
rect 10210 -1228 10244 -1194
rect 10336 -1228 10370 -1194
rect 11422 -1228 11456 -1194
rect 11548 -1228 11582 -1194
rect 12280 -1228 12314 -1194
rect 12721 -1230 12755 -1196
rect 12722 -1323 12756 -1289
rect 12981 -1305 13015 -1271
rect 6677 -1394 6707 -1364
rect 6707 -1394 6711 -1364
rect 6677 -1398 6711 -1394
rect 12982 -1398 13016 -1364
rect 13158 -1394 13162 -1363
rect 13162 -1394 13192 -1363
rect 13158 -1397 13192 -1394
rect 6596 -1562 6627 -1529
rect 6627 -1562 6630 -1529
rect 6596 -1563 6630 -1562
rect 12901 -1468 12935 -1434
rect 12857 -1587 12891 -1527
rect 12945 -1587 12979 -1527
rect 6356 -1706 6390 -1672
rect 6448 -1706 6482 -1672
rect 6540 -1706 6574 -1672
rect 6632 -1706 6666 -1672
rect 6724 -1706 6758 -1672
rect 12857 -1725 12891 -1665
rect 12945 -1725 12979 -1665
rect 13242 -1494 13276 -1474
rect 13242 -1508 13276 -1494
rect 13432 -1394 13462 -1364
rect 13462 -1394 13466 -1364
rect 13432 -1398 13466 -1394
rect 13351 -1562 13382 -1529
rect 13382 -1562 13385 -1529
rect 13351 -1563 13385 -1562
rect 13111 -1706 13145 -1672
rect 13203 -1706 13237 -1672
rect 13295 -1706 13329 -1672
rect 13387 -1706 13421 -1672
rect 13479 -1706 13513 -1672
rect 6102 -1863 6136 -1803
rect 6190 -1863 6224 -1803
rect 12857 -1863 12891 -1803
rect 12945 -1863 12979 -1803
rect 6102 -2001 6136 -1941
rect 6190 -2001 6224 -1941
rect 12857 -2001 12891 -1941
rect 12945 -2001 12979 -1941
rect 6102 -2139 6136 -2079
rect 6190 -2139 6224 -2079
rect 12857 -2139 12891 -2079
rect 12945 -2139 12979 -2079
rect 6102 -2277 6136 -2217
rect 6190 -2277 6224 -2217
rect 12857 -2277 12891 -2217
rect 12945 -2277 12979 -2217
<< metal1 >>
rect 725 3270 815 3286
rect 725 3259 744 3270
rect 619 3225 665 3237
rect 619 3165 625 3225
rect 659 3165 665 3225
rect 619 3087 665 3165
rect 707 3225 744 3259
rect 707 3165 713 3225
rect 796 3218 815 3270
rect 7414 3270 7504 3286
rect 7414 3259 7433 3270
rect 747 3203 815 3218
rect 7308 3225 7354 3237
rect 747 3165 753 3203
rect 707 3153 753 3165
rect 7308 3165 7314 3225
rect 7348 3165 7354 3225
rect 619 3027 625 3087
rect 659 3027 665 3087
rect 619 3015 665 3027
rect 707 3087 753 3099
rect 707 3027 713 3087
rect 747 3027 753 3087
rect 619 2949 665 2961
rect 619 2889 625 2949
rect 659 2889 665 2949
rect 619 2811 665 2889
rect 707 2949 753 3027
rect 7308 3087 7354 3165
rect 7396 3225 7433 3259
rect 7396 3165 7402 3225
rect 7485 3218 7504 3270
rect 7436 3203 7504 3218
rect 7436 3165 7442 3203
rect 7396 3153 7442 3165
rect 7308 3027 7314 3087
rect 7348 3027 7354 3087
rect 7308 3015 7354 3027
rect 7396 3087 7442 3099
rect 7396 3027 7402 3087
rect 7436 3027 7442 3087
rect 707 2889 713 2949
rect 747 2889 753 2949
rect 707 2877 753 2889
rect 7308 2949 7354 2961
rect 7308 2889 7314 2949
rect 7348 2889 7354 2949
rect 619 2751 625 2811
rect 659 2751 665 2811
rect 619 2739 665 2751
rect 707 2811 753 2823
rect 707 2751 713 2811
rect 747 2751 753 2811
rect 62 2665 522 2685
rect 62 2654 127 2665
rect 62 2620 91 2654
rect 125 2620 127 2654
rect 62 2613 127 2620
rect 179 2664 402 2665
rect 179 2654 258 2664
rect 310 2654 402 2664
rect 179 2620 183 2654
rect 217 2620 258 2654
rect 310 2620 367 2654
rect 401 2620 402 2654
rect 179 2613 258 2620
rect 62 2612 258 2613
rect 310 2613 402 2620
rect 454 2654 522 2665
rect 454 2620 459 2654
rect 493 2620 522 2654
rect 454 2613 522 2620
rect 310 2612 522 2613
rect 62 2589 522 2612
rect 619 2673 665 2685
rect 619 2613 625 2673
rect 659 2613 665 2673
rect 619 2535 665 2613
rect 707 2673 753 2751
rect 7308 2811 7354 2889
rect 7396 2949 7442 3027
rect 7396 2889 7402 2949
rect 7436 2889 7442 2949
rect 7396 2877 7442 2889
rect 7308 2751 7314 2811
rect 7348 2751 7354 2811
rect 7308 2739 7354 2751
rect 7396 2811 7442 2823
rect 7396 2751 7402 2811
rect 7436 2751 7442 2811
rect 707 2613 713 2673
rect 747 2613 753 2673
rect 707 2601 753 2613
rect 6751 2665 7211 2685
rect 6751 2654 6816 2665
rect 6751 2620 6780 2654
rect 6814 2620 6816 2654
rect 6751 2613 6816 2620
rect 6868 2664 7091 2665
rect 6868 2654 6947 2664
rect 6999 2654 7091 2664
rect 6868 2620 6872 2654
rect 6906 2620 6947 2654
rect 6999 2620 7056 2654
rect 7090 2620 7091 2654
rect 6868 2613 6947 2620
rect 6751 2612 6947 2613
rect 6999 2613 7091 2620
rect 7143 2654 7211 2665
rect 7143 2620 7148 2654
rect 7182 2620 7211 2654
rect 7143 2613 7211 2620
rect 6999 2612 7211 2613
rect 6751 2589 7211 2612
rect 7308 2673 7354 2685
rect 7308 2613 7314 2673
rect 7348 2613 7354 2673
rect 207 2511 579 2518
rect 207 2477 219 2511
rect 253 2490 579 2511
rect 253 2477 265 2490
rect 207 2470 265 2477
rect 312 2456 379 2462
rect 312 2422 328 2456
rect 362 2443 379 2456
rect 362 2422 523 2443
rect 312 2415 523 2422
rect 392 2354 458 2356
rect 130 2349 184 2353
rect 129 2346 184 2349
rect 0 2312 138 2346
rect 172 2312 184 2346
rect 129 2309 184 2312
rect 129 2305 183 2309
rect 392 2302 400 2354
rect 452 2302 458 2354
rect 392 2301 458 2302
rect 495 2271 523 2415
rect 551 2358 579 2490
rect 619 2475 625 2535
rect 659 2475 665 2535
rect 619 2463 665 2475
rect 707 2535 789 2547
rect 707 2475 713 2535
rect 747 2475 789 2535
rect 7308 2535 7354 2613
rect 7396 2673 7442 2751
rect 7396 2613 7402 2673
rect 7436 2613 7442 2673
rect 7396 2601 7442 2613
rect 707 2463 789 2475
rect 6896 2511 7268 2518
rect 6896 2477 6908 2511
rect 6942 2490 7268 2511
rect 6942 2477 6954 2490
rect 6896 2470 6954 2477
rect 657 2416 715 2422
rect 657 2382 669 2416
rect 703 2382 715 2416
rect 657 2376 715 2382
rect 551 2346 628 2358
rect 551 2312 588 2346
rect 622 2312 628 2346
rect 579 2299 628 2312
rect 495 2253 629 2271
rect 495 2243 589 2253
rect 580 2219 589 2243
rect 623 2219 629 2253
rect 580 2206 629 2219
rect 62 2119 522 2141
rect 62 2110 145 2119
rect 197 2110 265 2119
rect 317 2110 408 2119
rect 460 2110 522 2119
rect 62 2076 91 2110
rect 125 2076 145 2110
rect 217 2076 265 2110
rect 317 2076 367 2110
rect 401 2076 408 2110
rect 493 2076 522 2110
rect 62 2067 145 2076
rect 197 2067 265 2076
rect 317 2067 408 2076
rect 460 2067 522 2076
rect 62 2045 522 2067
rect 657 1976 705 2376
rect 37 1929 705 1976
rect 657 1788 705 1929
rect 647 1782 705 1788
rect 406 1776 471 1777
rect 406 1773 412 1776
rect 18 1726 412 1773
rect 406 1724 412 1726
rect 464 1724 471 1776
rect 647 1748 659 1782
rect 693 1748 705 1782
rect 647 1742 705 1748
rect 743 1973 789 2463
rect 7001 2456 7068 2462
rect 7001 2422 7017 2456
rect 7051 2443 7068 2456
rect 7051 2422 7212 2443
rect 7001 2415 7212 2422
rect 6457 2343 6547 2359
rect 7081 2354 7147 2356
rect 6819 2349 6873 2353
rect 6818 2346 6873 2349
rect 6457 2332 6476 2343
rect 6382 2291 6476 2332
rect 6528 2291 6547 2343
rect 6689 2312 6827 2346
rect 6861 2312 6873 2346
rect 6818 2309 6873 2312
rect 6818 2305 6872 2309
rect 7081 2302 7089 2354
rect 7141 2302 7147 2354
rect 7081 2301 7147 2302
rect 839 2276 888 2283
rect 839 2271 1458 2276
rect 839 2237 848 2271
rect 882 2237 1458 2271
rect 839 2229 1458 2237
rect 839 2224 888 2229
rect 840 2182 889 2190
rect 1409 2182 1458 2229
rect 6382 2273 6547 2291
rect 6382 2227 6429 2273
rect 7184 2271 7212 2415
rect 7240 2358 7268 2490
rect 7308 2475 7314 2535
rect 7348 2475 7354 2535
rect 7308 2463 7354 2475
rect 7396 2535 7478 2547
rect 7396 2475 7402 2535
rect 7436 2475 7478 2535
rect 7396 2463 7478 2475
rect 7346 2416 7404 2422
rect 7346 2382 7358 2416
rect 7392 2382 7404 2416
rect 7346 2376 7404 2382
rect 7240 2346 7317 2358
rect 7240 2312 7277 2346
rect 7311 2312 7317 2346
rect 7268 2299 7317 2312
rect 7184 2253 7318 2271
rect 7184 2243 7278 2253
rect 6383 2224 6429 2227
rect 840 2178 1341 2182
rect 840 2144 849 2178
rect 883 2176 1341 2178
rect 883 2144 1290 2176
rect 840 2142 1290 2144
rect 1324 2142 1341 2176
rect 840 2136 1341 2142
rect 1409 2176 5830 2182
rect 1409 2142 2022 2176
rect 2056 2142 2148 2176
rect 2182 2142 3234 2176
rect 3268 2142 3360 2176
rect 3394 2142 4446 2176
rect 4480 2142 4572 2176
rect 4606 2142 5658 2176
rect 5692 2142 5784 2176
rect 5818 2142 5830 2176
rect 6383 2164 6389 2224
rect 6423 2164 6429 2224
rect 6383 2152 6429 2164
rect 6471 2224 6517 2236
rect 6471 2164 6477 2224
rect 6511 2164 6517 2224
rect 7269 2219 7278 2243
rect 7312 2219 7318 2253
rect 7269 2206 7318 2219
rect 6471 2155 6517 2164
rect 1409 2136 5830 2142
rect 840 2135 1329 2136
rect 1409 2135 1855 2136
rect 840 2131 889 2135
rect 6471 2126 6709 2155
rect 1240 2087 1286 2095
rect 1217 2086 1296 2087
rect 1217 2022 1224 2086
rect 1288 2022 1296 2086
rect 1328 2083 1374 2095
rect 1972 2087 2018 2095
rect 1328 2023 1334 2083
rect 1368 2023 1374 2083
rect 1240 2011 1286 2022
rect 1328 1973 1374 2023
rect 1949 2086 2028 2087
rect 1949 2022 1956 2086
rect 2020 2022 2028 2086
rect 2077 2083 2123 2095
rect 2186 2087 2232 2095
rect 3184 2087 3230 2095
rect 2077 2023 2083 2083
rect 2117 2023 2123 2083
rect 1972 2011 2018 2022
rect 2077 1973 2123 2023
rect 2176 2086 2255 2087
rect 2176 2022 2184 2086
rect 2248 2022 2255 2086
rect 3161 2086 3240 2087
rect 3161 2022 3168 2086
rect 3232 2022 3240 2086
rect 3288 2083 3334 2095
rect 3398 2087 3444 2095
rect 4396 2087 4442 2095
rect 3288 2023 3294 2083
rect 3328 2023 3334 2083
rect 2186 2011 2232 2022
rect 3184 2011 3230 2022
rect 3288 1973 3334 2023
rect 3388 2086 3467 2087
rect 3388 2022 3396 2086
rect 3460 2022 3467 2086
rect 4373 2086 4452 2087
rect 4373 2022 4380 2086
rect 4444 2022 4452 2086
rect 4501 2083 4547 2095
rect 4610 2087 4656 2095
rect 5608 2087 5654 2095
rect 4501 2023 4507 2083
rect 4541 2023 4547 2083
rect 3398 2011 3444 2022
rect 4396 2011 4442 2022
rect 4501 1973 4547 2023
rect 4600 2086 4679 2087
rect 4600 2022 4608 2086
rect 4672 2022 4679 2086
rect 5585 2086 5664 2087
rect 5585 2022 5592 2086
rect 5656 2022 5664 2086
rect 5715 2083 5761 2095
rect 5822 2087 5868 2095
rect 5715 2023 5721 2083
rect 5755 2023 5761 2083
rect 4610 2011 4656 2022
rect 5608 2011 5654 2022
rect 5715 1973 5761 2023
rect 5812 2086 5891 2087
rect 5812 2022 5820 2086
rect 5884 2022 5891 2086
rect 6383 2086 6429 2098
rect 6383 2026 6389 2086
rect 6423 2026 6429 2086
rect 5822 2011 5868 2022
rect 6383 2014 6429 2026
rect 6471 2086 6517 2126
rect 6471 2026 6477 2086
rect 6511 2026 6517 2086
rect 6471 2014 6517 2026
rect 6545 2086 6635 2098
rect 6545 2082 6573 2086
rect 6607 2082 6635 2086
rect 6545 2030 6564 2082
rect 6616 2030 6635 2082
rect 6545 2026 6573 2030
rect 6607 2026 6635 2030
rect 6545 2014 6635 2026
rect 6663 2086 6709 2126
rect 6663 2026 6669 2086
rect 6703 2026 6709 2086
rect 6751 2119 7211 2141
rect 6751 2110 6834 2119
rect 6886 2110 6954 2119
rect 7006 2110 7097 2119
rect 7149 2110 7211 2119
rect 6751 2076 6780 2110
rect 6814 2076 6834 2110
rect 6906 2076 6954 2110
rect 7006 2076 7056 2110
rect 7090 2076 7097 2110
rect 7182 2076 7211 2110
rect 6751 2067 6834 2076
rect 6886 2067 6954 2076
rect 7006 2067 7097 2076
rect 7149 2067 7211 2076
rect 6751 2045 7211 2067
rect 6663 2014 6709 2026
rect 6302 1973 6368 1975
rect 743 1969 6368 1973
rect 743 1935 6318 1969
rect 6352 1935 6368 1969
rect 743 1931 6368 1935
rect 743 1710 789 1931
rect 1595 1884 1641 1894
rect 1573 1820 1582 1884
rect 1646 1820 1655 1884
rect 1573 1819 1655 1820
rect 1683 1882 1729 1931
rect 2327 1884 2373 1894
rect 1683 1822 1689 1882
rect 1723 1822 1729 1882
rect 1595 1810 1641 1819
rect 1683 1810 1729 1822
rect 2305 1820 2314 1884
rect 2378 1820 2387 1884
rect 2305 1819 2387 1820
rect 2432 1882 2478 1931
rect 2539 1884 2585 1894
rect 3539 1884 3585 1894
rect 2432 1822 2438 1882
rect 2472 1822 2478 1882
rect 2327 1810 2373 1819
rect 2432 1810 2478 1822
rect 2525 1820 2534 1884
rect 2598 1820 2607 1884
rect 2525 1819 2607 1820
rect 3517 1820 3526 1884
rect 3590 1820 3599 1884
rect 3517 1819 3599 1820
rect 3643 1882 3689 1931
rect 3751 1884 3797 1894
rect 4877 1884 4923 1894
rect 3643 1822 3649 1882
rect 3683 1822 3689 1882
rect 2539 1810 2585 1819
rect 3539 1810 3585 1819
rect 3643 1810 3689 1822
rect 3737 1820 3746 1884
rect 3810 1820 3819 1884
rect 3737 1819 3819 1820
rect 4855 1820 4864 1884
rect 4928 1820 4937 1884
rect 4855 1819 4937 1820
rect 4983 1882 5029 1931
rect 5089 1884 5135 1894
rect 4983 1822 4989 1882
rect 5023 1822 5029 1882
rect 3751 1810 3797 1819
rect 4877 1810 4923 1819
rect 4983 1810 5029 1822
rect 5075 1820 5084 1884
rect 5148 1820 5157 1884
rect 5075 1819 5157 1820
rect 5732 1882 5778 1931
rect 6306 1929 6368 1931
rect 6401 1966 6429 2014
rect 7346 1976 7394 2376
rect 6726 1974 7394 1976
rect 6674 1973 7394 1974
rect 6513 1967 7394 1973
rect 6513 1966 6525 1967
rect 6401 1937 6525 1966
rect 6401 1895 6429 1937
rect 6513 1933 6525 1937
rect 6559 1933 7394 1967
rect 6513 1930 7394 1933
rect 6513 1927 6695 1930
rect 6726 1929 7394 1930
rect 5821 1884 5867 1894
rect 5732 1822 5738 1882
rect 5772 1822 5778 1882
rect 5089 1810 5135 1819
rect 5732 1810 5778 1822
rect 5807 1820 5816 1884
rect 5880 1820 5889 1884
rect 5807 1819 5889 1820
rect 6383 1883 6429 1895
rect 6383 1823 6389 1883
rect 6423 1823 6429 1883
rect 5821 1810 5867 1819
rect 6383 1811 6429 1823
rect 6471 1883 6517 1895
rect 6471 1823 6477 1883
rect 6511 1823 6517 1883
rect 6471 1783 6517 1823
rect 6545 1883 6635 1895
rect 6545 1879 6573 1883
rect 6607 1879 6635 1883
rect 6545 1827 6564 1879
rect 6616 1827 6635 1879
rect 6545 1823 6573 1827
rect 6607 1823 6635 1827
rect 6545 1811 6635 1823
rect 6663 1883 6709 1895
rect 6663 1823 6669 1883
rect 6703 1823 6709 1883
rect 6663 1783 6709 1823
rect 7346 1788 7394 1929
rect 893 1724 900 1776
rect 952 1774 958 1776
rect 1633 1774 1691 1778
rect 952 1772 1691 1774
rect 952 1738 1645 1772
rect 1679 1738 1691 1772
rect 952 1727 1691 1738
rect 2365 1772 3759 1778
rect 2365 1738 2377 1772
rect 2411 1738 2501 1772
rect 2535 1738 3589 1772
rect 3623 1738 3713 1772
rect 3747 1738 3759 1772
rect 2365 1732 3759 1738
rect 4915 1772 5097 1778
rect 4915 1738 4927 1772
rect 4961 1738 5051 1772
rect 5085 1738 5097 1772
rect 4915 1732 5097 1738
rect 5771 1772 5829 1778
rect 5771 1738 5783 1772
rect 5817 1738 5829 1772
rect 6471 1773 6709 1783
rect 7336 1782 7394 1788
rect 7095 1776 7160 1777
rect 7095 1773 7101 1776
rect 952 1724 958 1727
rect 893 1723 958 1724
rect 1633 1722 1691 1727
rect 573 1698 619 1710
rect 573 1638 579 1698
rect 613 1638 619 1698
rect 573 1560 619 1638
rect 733 1698 789 1710
rect 733 1638 739 1698
rect 773 1638 789 1698
rect 733 1626 789 1638
rect 573 1500 579 1560
rect 613 1500 619 1560
rect 573 1488 619 1500
rect 733 1560 779 1572
rect 733 1500 739 1560
rect 773 1500 779 1560
rect 573 1422 619 1434
rect 573 1362 579 1422
rect 613 1362 619 1422
rect 573 1284 619 1362
rect 733 1422 779 1500
rect 733 1362 739 1422
rect 773 1362 779 1422
rect 733 1350 779 1362
rect 573 1224 579 1284
rect 613 1224 619 1284
rect 573 1212 619 1224
rect 733 1284 779 1296
rect 733 1224 739 1284
rect 773 1224 779 1284
rect 573 1146 619 1158
rect 573 1086 579 1146
rect 613 1086 619 1146
rect 573 1008 619 1086
rect 733 1146 779 1224
rect 733 1086 739 1146
rect 773 1086 779 1146
rect 733 1074 779 1086
rect 573 948 579 1008
rect 613 948 619 1008
rect 573 936 619 948
rect 733 1008 779 1020
rect 733 948 739 1008
rect 773 948 779 1008
rect 573 870 619 882
rect 573 810 579 870
rect 613 810 619 870
rect 573 732 619 810
rect 733 870 779 948
rect 733 810 739 870
rect 773 810 779 870
rect 733 798 779 810
rect 573 672 579 732
rect 613 672 619 732
rect 733 732 779 744
rect 733 708 739 732
rect 573 660 619 672
rect 694 692 739 708
rect 773 708 779 732
rect 773 692 801 708
rect 694 640 730 692
rect 782 640 801 692
rect 694 624 801 640
rect 2489 601 2547 1732
rect 4915 601 4973 1732
rect 5771 600 5829 1738
rect 6383 1745 6429 1757
rect 6383 1685 6389 1745
rect 6423 1685 6429 1745
rect 6383 1633 6429 1685
rect 6471 1754 7101 1773
rect 6471 1745 6517 1754
rect 6471 1685 6477 1745
rect 6511 1685 6517 1745
rect 6707 1726 7101 1754
rect 7095 1724 7101 1726
rect 7153 1724 7160 1776
rect 7336 1748 7348 1782
rect 7382 1748 7394 1782
rect 7336 1742 7394 1748
rect 7432 1973 7478 2463
rect 13146 2343 13236 2359
rect 13146 2332 13165 2343
rect 13071 2291 13165 2332
rect 13217 2291 13236 2343
rect 7528 2276 7577 2283
rect 7528 2271 8147 2276
rect 7528 2237 7537 2271
rect 7571 2237 8147 2271
rect 7528 2229 8147 2237
rect 7528 2224 7577 2229
rect 7529 2182 7578 2190
rect 8098 2182 8147 2229
rect 13071 2273 13236 2291
rect 13071 2227 13118 2273
rect 13072 2224 13118 2227
rect 7529 2178 8030 2182
rect 7529 2144 7538 2178
rect 7572 2176 8030 2178
rect 7572 2144 7979 2176
rect 7529 2142 7979 2144
rect 8013 2142 8030 2176
rect 7529 2136 8030 2142
rect 8098 2176 12519 2182
rect 8098 2142 8711 2176
rect 8745 2142 8837 2176
rect 8871 2142 9923 2176
rect 9957 2142 10049 2176
rect 10083 2142 11135 2176
rect 11169 2142 11261 2176
rect 11295 2142 12347 2176
rect 12381 2142 12473 2176
rect 12507 2142 12519 2176
rect 13072 2164 13078 2224
rect 13112 2164 13118 2224
rect 13072 2152 13118 2164
rect 13160 2224 13206 2236
rect 13160 2164 13166 2224
rect 13200 2164 13206 2224
rect 13160 2155 13206 2164
rect 8098 2136 12519 2142
rect 7529 2135 8018 2136
rect 8098 2135 8544 2136
rect 7529 2131 7578 2135
rect 13160 2126 13398 2155
rect 7929 2087 7975 2095
rect 7906 2086 7985 2087
rect 7906 2022 7913 2086
rect 7977 2022 7985 2086
rect 8017 2083 8063 2095
rect 8661 2087 8707 2095
rect 8017 2023 8023 2083
rect 8057 2023 8063 2083
rect 7929 2011 7975 2022
rect 8017 1973 8063 2023
rect 8638 2086 8717 2087
rect 8638 2022 8645 2086
rect 8709 2022 8717 2086
rect 8766 2083 8812 2095
rect 8875 2087 8921 2095
rect 9873 2087 9919 2095
rect 8766 2023 8772 2083
rect 8806 2023 8812 2083
rect 8661 2011 8707 2022
rect 8766 1973 8812 2023
rect 8865 2086 8944 2087
rect 8865 2022 8873 2086
rect 8937 2022 8944 2086
rect 9850 2086 9929 2087
rect 9850 2022 9857 2086
rect 9921 2022 9929 2086
rect 9977 2083 10023 2095
rect 10087 2087 10133 2095
rect 11085 2087 11131 2095
rect 9977 2023 9983 2083
rect 10017 2023 10023 2083
rect 8875 2011 8921 2022
rect 9873 2011 9919 2022
rect 9977 1973 10023 2023
rect 10077 2086 10156 2087
rect 10077 2022 10085 2086
rect 10149 2022 10156 2086
rect 11062 2086 11141 2087
rect 11062 2022 11069 2086
rect 11133 2022 11141 2086
rect 11190 2083 11236 2095
rect 11299 2087 11345 2095
rect 12297 2087 12343 2095
rect 11190 2023 11196 2083
rect 11230 2023 11236 2083
rect 10087 2011 10133 2022
rect 11085 2011 11131 2022
rect 11190 1973 11236 2023
rect 11289 2086 11368 2087
rect 11289 2022 11297 2086
rect 11361 2022 11368 2086
rect 12274 2086 12353 2087
rect 12274 2022 12281 2086
rect 12345 2022 12353 2086
rect 12404 2083 12450 2095
rect 12511 2087 12557 2095
rect 12404 2023 12410 2083
rect 12444 2023 12450 2083
rect 11299 2011 11345 2022
rect 12297 2011 12343 2022
rect 12404 1973 12450 2023
rect 12501 2086 12580 2087
rect 12501 2022 12509 2086
rect 12573 2022 12580 2086
rect 13072 2086 13118 2098
rect 13072 2026 13078 2086
rect 13112 2026 13118 2086
rect 12511 2011 12557 2022
rect 13072 2014 13118 2026
rect 13160 2086 13206 2126
rect 13160 2026 13166 2086
rect 13200 2026 13206 2086
rect 13160 2014 13206 2026
rect 13234 2086 13324 2098
rect 13234 2082 13262 2086
rect 13296 2082 13324 2086
rect 13234 2030 13253 2082
rect 13305 2030 13324 2082
rect 13234 2026 13262 2030
rect 13296 2026 13324 2030
rect 13234 2014 13324 2026
rect 13352 2086 13398 2126
rect 13352 2026 13358 2086
rect 13392 2026 13398 2086
rect 13352 2014 13398 2026
rect 12991 1973 13057 1975
rect 7432 1969 13057 1973
rect 7432 1935 13007 1969
rect 13041 1935 13057 1969
rect 7432 1931 13057 1935
rect 7432 1710 7478 1931
rect 8284 1884 8330 1894
rect 8262 1820 8271 1884
rect 8335 1820 8344 1884
rect 8262 1819 8344 1820
rect 8372 1882 8418 1931
rect 9016 1884 9062 1894
rect 8372 1822 8378 1882
rect 8412 1822 8418 1882
rect 8284 1810 8330 1819
rect 8372 1810 8418 1822
rect 8994 1820 9003 1884
rect 9067 1820 9076 1884
rect 8994 1819 9076 1820
rect 9121 1882 9167 1931
rect 9228 1884 9274 1894
rect 10228 1884 10274 1894
rect 9121 1822 9127 1882
rect 9161 1822 9167 1882
rect 9016 1810 9062 1819
rect 9121 1810 9167 1822
rect 9214 1820 9223 1884
rect 9287 1820 9296 1884
rect 9214 1819 9296 1820
rect 10206 1820 10215 1884
rect 10279 1820 10288 1884
rect 10206 1819 10288 1820
rect 10332 1882 10378 1931
rect 10440 1884 10486 1894
rect 11566 1884 11612 1894
rect 10332 1822 10338 1882
rect 10372 1822 10378 1882
rect 9228 1810 9274 1819
rect 10228 1810 10274 1819
rect 10332 1810 10378 1822
rect 10426 1820 10435 1884
rect 10499 1820 10508 1884
rect 10426 1819 10508 1820
rect 11544 1820 11553 1884
rect 11617 1820 11626 1884
rect 11544 1819 11626 1820
rect 11672 1882 11718 1931
rect 11778 1884 11824 1894
rect 11672 1822 11678 1882
rect 11712 1822 11718 1882
rect 10440 1810 10486 1819
rect 11566 1810 11612 1819
rect 11672 1810 11718 1822
rect 11764 1820 11773 1884
rect 11837 1820 11846 1884
rect 11764 1819 11846 1820
rect 12421 1882 12467 1931
rect 12995 1929 13057 1931
rect 13090 1966 13118 2014
rect 13202 1967 13384 1973
rect 13202 1966 13214 1967
rect 13090 1937 13214 1966
rect 13090 1895 13118 1937
rect 13202 1933 13214 1937
rect 13248 1933 13384 1967
rect 13202 1927 13384 1933
rect 12510 1884 12556 1894
rect 12421 1822 12427 1882
rect 12461 1822 12467 1882
rect 11778 1810 11824 1819
rect 12421 1810 12467 1822
rect 12496 1820 12505 1884
rect 12569 1820 12578 1884
rect 12496 1819 12578 1820
rect 13072 1883 13118 1895
rect 13072 1823 13078 1883
rect 13112 1823 13118 1883
rect 12510 1810 12556 1819
rect 13072 1811 13118 1823
rect 13160 1883 13206 1895
rect 13160 1823 13166 1883
rect 13200 1823 13206 1883
rect 13160 1783 13206 1823
rect 13234 1883 13324 1895
rect 13234 1879 13262 1883
rect 13296 1879 13324 1883
rect 13234 1827 13253 1879
rect 13305 1827 13324 1879
rect 13234 1823 13262 1827
rect 13296 1823 13324 1827
rect 13234 1811 13324 1823
rect 13352 1883 13398 1895
rect 13352 1823 13358 1883
rect 13392 1823 13398 1883
rect 13352 1783 13398 1823
rect 7582 1724 7589 1776
rect 7641 1774 7647 1776
rect 8322 1774 8380 1778
rect 7641 1772 8380 1774
rect 7641 1738 8334 1772
rect 8368 1738 8380 1772
rect 7641 1727 8380 1738
rect 9054 1772 10448 1778
rect 9054 1738 9066 1772
rect 9100 1738 9190 1772
rect 9224 1738 10278 1772
rect 10312 1738 10402 1772
rect 10436 1738 10448 1772
rect 9054 1732 10448 1738
rect 11604 1772 11786 1778
rect 11604 1738 11616 1772
rect 11650 1738 11740 1772
rect 11774 1738 11786 1772
rect 11604 1732 11786 1738
rect 12460 1772 12518 1778
rect 12460 1738 12472 1772
rect 12506 1738 12518 1772
rect 7641 1724 7647 1727
rect 7582 1723 7647 1724
rect 8322 1722 8380 1727
rect 6471 1673 6517 1685
rect 7262 1698 7308 1710
rect 7262 1638 7268 1698
rect 7302 1638 7308 1698
rect 6383 1617 6544 1633
rect 6383 1565 6473 1617
rect 6525 1565 6544 1617
rect 6383 1549 6544 1565
rect 7262 1560 7308 1638
rect 7422 1698 7478 1710
rect 7422 1638 7428 1698
rect 7462 1638 7478 1698
rect 7422 1626 7478 1638
rect 7262 1500 7268 1560
rect 7302 1500 7308 1560
rect 7262 1488 7308 1500
rect 7422 1560 7468 1572
rect 7422 1500 7428 1560
rect 7462 1500 7468 1560
rect 7262 1422 7308 1434
rect 7262 1362 7268 1422
rect 7302 1362 7308 1422
rect 7262 1284 7308 1362
rect 7422 1422 7468 1500
rect 7422 1362 7428 1422
rect 7462 1362 7468 1422
rect 7422 1350 7468 1362
rect 7262 1224 7268 1284
rect 7302 1224 7308 1284
rect 7262 1212 7308 1224
rect 7422 1284 7468 1296
rect 7422 1224 7428 1284
rect 7462 1224 7468 1284
rect 7262 1146 7308 1158
rect 7262 1086 7268 1146
rect 7302 1086 7308 1146
rect 7262 1008 7308 1086
rect 7422 1146 7468 1224
rect 7422 1086 7428 1146
rect 7462 1086 7468 1146
rect 7422 1074 7468 1086
rect 7262 948 7268 1008
rect 7302 948 7308 1008
rect 7262 936 7308 948
rect 7422 1008 7468 1020
rect 7422 948 7428 1008
rect 7462 948 7468 1008
rect 7262 870 7308 882
rect 7262 810 7268 870
rect 7302 810 7308 870
rect 7262 732 7308 810
rect 7422 870 7468 948
rect 7422 810 7428 870
rect 7462 810 7468 870
rect 7422 798 7468 810
rect 7262 672 7268 732
rect 7302 672 7308 732
rect 7422 732 7468 744
rect 7422 708 7428 732
rect 7262 660 7308 672
rect 7383 692 7428 708
rect 7462 708 7468 732
rect 7462 692 7490 708
rect 7383 640 7419 692
rect 7471 640 7490 692
rect 7383 624 7490 640
rect 9178 601 9236 1732
rect 11604 601 11662 1732
rect 12460 600 12518 1738
rect 13072 1745 13118 1757
rect 13072 1685 13078 1745
rect 13112 1685 13118 1745
rect 13072 1633 13118 1685
rect 13160 1754 13398 1783
rect 13160 1745 13206 1754
rect 13160 1685 13166 1745
rect 13200 1685 13206 1745
rect 13160 1673 13206 1685
rect 13072 1617 13233 1633
rect 13072 1565 13162 1617
rect 13214 1565 13233 1617
rect 13072 1549 13233 1565
rect 305 -617 466 -601
rect 305 -669 324 -617
rect 376 -669 466 -617
rect 305 -685 466 -669
rect 332 -737 378 -725
rect 332 -797 338 -737
rect 372 -797 378 -737
rect 332 -806 378 -797
rect 140 -835 378 -806
rect 420 -737 466 -685
rect 420 -797 426 -737
rect 460 -797 466 -737
rect 420 -809 466 -797
rect 1020 -790 1078 348
rect 1876 -784 1934 347
rect 4302 -784 4360 347
rect 6048 308 6155 324
rect 6048 256 6067 308
rect 6119 256 6155 308
rect 6048 240 6076 256
rect 6070 216 6076 240
rect 6110 240 6155 256
rect 6230 276 6276 288
rect 6110 216 6116 240
rect 6070 204 6116 216
rect 6230 216 6236 276
rect 6270 216 6276 276
rect 6070 138 6116 150
rect 6070 78 6076 138
rect 6110 78 6116 138
rect 6070 0 6116 78
rect 6230 138 6276 216
rect 6230 78 6236 138
rect 6270 78 6276 138
rect 6230 66 6276 78
rect 6070 -60 6076 0
rect 6110 -60 6116 0
rect 6070 -72 6116 -60
rect 6230 0 6276 12
rect 6230 -60 6236 0
rect 6270 -60 6276 0
rect 6070 -138 6116 -126
rect 6070 -198 6076 -138
rect 6110 -198 6116 -138
rect 6070 -276 6116 -198
rect 6230 -138 6276 -60
rect 6230 -198 6236 -138
rect 6270 -198 6276 -138
rect 6230 -210 6276 -198
rect 6070 -336 6076 -276
rect 6110 -336 6116 -276
rect 6070 -348 6116 -336
rect 6230 -276 6276 -264
rect 6230 -336 6236 -276
rect 6270 -336 6276 -276
rect 6070 -414 6116 -402
rect 6070 -474 6076 -414
rect 6110 -474 6116 -414
rect 6070 -552 6116 -474
rect 6230 -414 6276 -336
rect 6230 -474 6236 -414
rect 6270 -474 6276 -414
rect 6230 -486 6276 -474
rect 6070 -612 6076 -552
rect 6110 -612 6116 -552
rect 6070 -624 6116 -612
rect 6230 -552 6276 -540
rect 6230 -612 6236 -552
rect 6270 -612 6276 -552
rect 6060 -690 6116 -678
rect 6060 -750 6076 -690
rect 6110 -750 6116 -690
rect 6060 -762 6116 -750
rect 6230 -690 6276 -612
rect 7060 -617 7221 -601
rect 7060 -669 7079 -617
rect 7131 -669 7221 -617
rect 7060 -685 7221 -669
rect 6230 -750 6236 -690
rect 6270 -750 6276 -690
rect 6230 -762 6276 -750
rect 7087 -737 7133 -725
rect 5158 -779 5216 -774
rect 5891 -776 5956 -775
rect 5891 -779 5897 -776
rect 1020 -824 1032 -790
rect 1066 -824 1078 -790
rect 1020 -830 1078 -824
rect 1752 -790 1934 -784
rect 1752 -824 1764 -790
rect 1798 -824 1888 -790
rect 1922 -824 1934 -790
rect 1752 -830 1934 -824
rect 3090 -790 4484 -784
rect 3090 -824 3102 -790
rect 3136 -824 3226 -790
rect 3260 -824 4314 -790
rect 4348 -824 4438 -790
rect 4472 -824 4484 -790
rect 3090 -830 4484 -824
rect 5158 -790 5897 -779
rect 5158 -824 5170 -790
rect 5204 -824 5897 -790
rect 5158 -826 5897 -824
rect 5158 -830 5216 -826
rect 5891 -828 5897 -826
rect 5949 -828 5956 -776
rect 140 -875 186 -835
rect 140 -935 146 -875
rect 180 -935 186 -875
rect 140 -947 186 -935
rect 214 -875 304 -863
rect 214 -879 242 -875
rect 276 -879 304 -875
rect 214 -931 233 -879
rect 285 -931 304 -879
rect 214 -935 242 -931
rect 276 -935 304 -931
rect 214 -947 304 -935
rect 332 -875 378 -835
rect 332 -935 338 -875
rect 372 -935 378 -875
rect 332 -947 378 -935
rect 420 -875 466 -863
rect 982 -871 1028 -862
rect 420 -935 426 -875
rect 460 -935 466 -875
rect 420 -947 466 -935
rect 960 -872 1042 -871
rect 960 -936 969 -872
rect 1033 -936 1042 -872
rect 1071 -874 1117 -862
rect 1714 -871 1760 -862
rect 1071 -934 1077 -874
rect 1111 -934 1117 -874
rect 982 -946 1028 -936
rect 154 -985 336 -979
rect 154 -1019 290 -985
rect 324 -989 336 -985
rect 420 -989 448 -947
rect 324 -1018 448 -989
rect 324 -1019 336 -1018
rect 154 -1025 336 -1019
rect 420 -1066 448 -1018
rect 481 -983 543 -981
rect 1071 -983 1117 -934
rect 1692 -872 1774 -871
rect 1692 -936 1701 -872
rect 1765 -936 1774 -872
rect 1820 -874 1866 -862
rect 1926 -871 1972 -862
rect 3052 -871 3098 -862
rect 1820 -934 1826 -874
rect 1860 -934 1866 -874
rect 1714 -946 1760 -936
rect 1820 -983 1866 -934
rect 1912 -872 1994 -871
rect 1912 -936 1921 -872
rect 1985 -936 1994 -872
rect 3030 -872 3112 -871
rect 3030 -936 3039 -872
rect 3103 -936 3112 -872
rect 3160 -874 3206 -862
rect 3264 -871 3310 -862
rect 4264 -871 4310 -862
rect 3160 -934 3166 -874
rect 3200 -934 3206 -874
rect 1926 -946 1972 -936
rect 3052 -946 3098 -936
rect 3160 -983 3206 -934
rect 3250 -872 3332 -871
rect 3250 -936 3259 -872
rect 3323 -936 3332 -872
rect 4242 -872 4324 -871
rect 4242 -936 4251 -872
rect 4315 -936 4324 -872
rect 4371 -874 4417 -862
rect 4476 -871 4522 -862
rect 4371 -934 4377 -874
rect 4411 -934 4417 -874
rect 3264 -946 3310 -936
rect 4264 -946 4310 -936
rect 4371 -983 4417 -934
rect 4462 -872 4544 -871
rect 4462 -936 4471 -872
rect 4535 -936 4544 -872
rect 5120 -874 5166 -862
rect 5208 -871 5254 -862
rect 5120 -934 5126 -874
rect 5160 -934 5166 -874
rect 4476 -946 4522 -936
rect 5120 -983 5166 -934
rect 5194 -872 5276 -871
rect 5194 -936 5203 -872
rect 5267 -936 5276 -872
rect 5208 -946 5254 -936
rect 6060 -983 6106 -762
rect 481 -987 6106 -983
rect 481 -1021 497 -987
rect 531 -1021 6106 -987
rect 481 -1025 6106 -1021
rect 481 -1027 547 -1025
rect 140 -1078 186 -1066
rect 140 -1138 146 -1078
rect 180 -1138 186 -1078
rect 140 -1178 186 -1138
rect 214 -1078 304 -1066
rect 214 -1082 242 -1078
rect 276 -1082 304 -1078
rect 214 -1134 233 -1082
rect 285 -1134 304 -1082
rect 214 -1138 242 -1134
rect 276 -1138 304 -1134
rect 214 -1150 304 -1138
rect 332 -1078 378 -1066
rect 332 -1138 338 -1078
rect 372 -1138 378 -1078
rect 332 -1178 378 -1138
rect 420 -1078 466 -1066
rect 981 -1074 1027 -1063
rect 420 -1138 426 -1078
rect 460 -1138 466 -1078
rect 420 -1150 466 -1138
rect 958 -1138 965 -1074
rect 1029 -1138 1037 -1074
rect 958 -1139 1037 -1138
rect 1088 -1075 1134 -1025
rect 1195 -1074 1241 -1063
rect 2193 -1074 2239 -1063
rect 1088 -1135 1094 -1075
rect 1128 -1135 1134 -1075
rect 981 -1147 1027 -1139
rect 1088 -1147 1134 -1135
rect 1185 -1138 1193 -1074
rect 1257 -1138 1264 -1074
rect 1185 -1139 1264 -1138
rect 2170 -1138 2177 -1074
rect 2241 -1138 2249 -1074
rect 2170 -1139 2249 -1138
rect 2302 -1075 2348 -1025
rect 2407 -1074 2453 -1063
rect 3405 -1074 3451 -1063
rect 2302 -1135 2308 -1075
rect 2342 -1135 2348 -1075
rect 1195 -1147 1241 -1139
rect 2193 -1147 2239 -1139
rect 2302 -1147 2348 -1135
rect 2397 -1138 2405 -1074
rect 2469 -1138 2476 -1074
rect 2397 -1139 2476 -1138
rect 3382 -1138 3389 -1074
rect 3453 -1138 3461 -1074
rect 3382 -1139 3461 -1138
rect 3515 -1075 3561 -1025
rect 3619 -1074 3665 -1063
rect 4617 -1074 4663 -1063
rect 3515 -1135 3521 -1075
rect 3555 -1135 3561 -1075
rect 2407 -1147 2453 -1139
rect 3405 -1147 3451 -1139
rect 3515 -1147 3561 -1135
rect 3609 -1138 3617 -1074
rect 3681 -1138 3688 -1074
rect 3609 -1139 3688 -1138
rect 4594 -1138 4601 -1074
rect 4665 -1138 4673 -1074
rect 4594 -1139 4673 -1138
rect 4726 -1075 4772 -1025
rect 4831 -1074 4877 -1063
rect 4726 -1135 4732 -1075
rect 4766 -1135 4772 -1075
rect 3619 -1147 3665 -1139
rect 4617 -1147 4663 -1139
rect 4726 -1147 4772 -1135
rect 4821 -1138 4829 -1074
rect 4893 -1138 4900 -1074
rect 4821 -1139 4900 -1138
rect 5475 -1075 5521 -1025
rect 5563 -1074 5609 -1063
rect 5475 -1135 5481 -1075
rect 5515 -1135 5521 -1075
rect 4831 -1147 4877 -1139
rect 5475 -1147 5521 -1135
rect 5553 -1138 5561 -1074
rect 5625 -1138 5632 -1074
rect 5553 -1139 5632 -1138
rect 5563 -1147 5609 -1139
rect 140 -1207 378 -1178
rect 5960 -1187 6009 -1183
rect 4994 -1188 5440 -1187
rect 5520 -1188 6009 -1187
rect 1019 -1194 5440 -1188
rect 332 -1216 378 -1207
rect 332 -1276 338 -1216
rect 372 -1276 378 -1216
rect 332 -1288 378 -1276
rect 420 -1216 466 -1204
rect 420 -1276 426 -1216
rect 460 -1276 466 -1216
rect 1019 -1228 1031 -1194
rect 1065 -1228 1157 -1194
rect 1191 -1228 2243 -1194
rect 2277 -1228 2369 -1194
rect 2403 -1228 3455 -1194
rect 3489 -1228 3581 -1194
rect 3615 -1228 4667 -1194
rect 4701 -1228 4793 -1194
rect 4827 -1228 5440 -1194
rect 1019 -1234 5440 -1228
rect 5508 -1194 6009 -1188
rect 5508 -1228 5525 -1194
rect 5559 -1196 6009 -1194
rect 5559 -1228 5966 -1196
rect 5508 -1230 5966 -1228
rect 6000 -1230 6009 -1196
rect 5508 -1234 6009 -1230
rect 420 -1279 466 -1276
rect 420 -1325 467 -1279
rect 302 -1343 467 -1325
rect 5391 -1281 5440 -1234
rect 5960 -1242 6009 -1234
rect 5961 -1281 6010 -1276
rect 5391 -1289 6010 -1281
rect 5391 -1323 5967 -1289
rect 6001 -1323 6010 -1289
rect 5391 -1328 6010 -1323
rect 5961 -1335 6010 -1328
rect 302 -1395 321 -1343
rect 373 -1384 467 -1343
rect 373 -1395 392 -1384
rect 302 -1411 392 -1395
rect 6060 -1515 6106 -1025
rect 6144 -800 6202 -794
rect 6144 -834 6156 -800
rect 6190 -834 6202 -800
rect 6378 -828 6385 -776
rect 6437 -778 6443 -776
rect 6437 -825 6831 -778
rect 7087 -797 7093 -737
rect 7127 -797 7133 -737
rect 7087 -806 7133 -797
rect 6437 -828 6443 -825
rect 6378 -829 6443 -828
rect 6144 -840 6202 -834
rect 6895 -835 7133 -806
rect 7175 -737 7221 -685
rect 7175 -797 7181 -737
rect 7215 -797 7221 -737
rect 7175 -809 7221 -797
rect 7775 -790 7833 348
rect 8631 -784 8689 347
rect 11057 -784 11115 347
rect 12803 308 12910 324
rect 12803 256 12822 308
rect 12874 256 12910 308
rect 12803 240 12831 256
rect 12825 216 12831 240
rect 12865 240 12910 256
rect 12985 276 13031 288
rect 12865 216 12871 240
rect 12825 204 12871 216
rect 12985 216 12991 276
rect 13025 216 13031 276
rect 12825 138 12871 150
rect 12825 78 12831 138
rect 12865 78 12871 138
rect 12825 0 12871 78
rect 12985 138 13031 216
rect 12985 78 12991 138
rect 13025 78 13031 138
rect 12985 66 13031 78
rect 12825 -60 12831 0
rect 12865 -60 12871 0
rect 12825 -72 12871 -60
rect 12985 0 13031 12
rect 12985 -60 12991 0
rect 13025 -60 13031 0
rect 12825 -138 12871 -126
rect 12825 -198 12831 -138
rect 12865 -198 12871 -138
rect 12825 -276 12871 -198
rect 12985 -138 13031 -60
rect 12985 -198 12991 -138
rect 13025 -198 13031 -138
rect 12985 -210 13031 -198
rect 12825 -336 12831 -276
rect 12865 -336 12871 -276
rect 12825 -348 12871 -336
rect 12985 -276 13031 -264
rect 12985 -336 12991 -276
rect 13025 -336 13031 -276
rect 12825 -414 12871 -402
rect 12825 -474 12831 -414
rect 12865 -474 12871 -414
rect 12825 -552 12871 -474
rect 12985 -414 13031 -336
rect 12985 -474 12991 -414
rect 13025 -474 13031 -414
rect 12985 -486 13031 -474
rect 12825 -612 12831 -552
rect 12865 -612 12871 -552
rect 12825 -624 12871 -612
rect 12985 -552 13031 -540
rect 12985 -612 12991 -552
rect 13025 -612 13031 -552
rect 12815 -690 12871 -678
rect 12815 -750 12831 -690
rect 12865 -750 12871 -690
rect 12815 -762 12871 -750
rect 12985 -690 13031 -612
rect 12985 -750 12991 -690
rect 13025 -750 13031 -690
rect 12985 -762 13031 -750
rect 11913 -779 11971 -774
rect 12646 -776 12711 -775
rect 12646 -779 12652 -776
rect 7775 -824 7787 -790
rect 7821 -824 7833 -790
rect 7775 -830 7833 -824
rect 8507 -790 8689 -784
rect 8507 -824 8519 -790
rect 8553 -824 8643 -790
rect 8677 -824 8689 -790
rect 8507 -830 8689 -824
rect 9845 -790 11239 -784
rect 9845 -824 9857 -790
rect 9891 -824 9981 -790
rect 10015 -824 11069 -790
rect 11103 -824 11193 -790
rect 11227 -824 11239 -790
rect 9845 -830 11239 -824
rect 11913 -790 12652 -779
rect 11913 -824 11925 -790
rect 11959 -824 12652 -790
rect 11913 -826 12652 -824
rect 11913 -830 11971 -826
rect 12646 -828 12652 -826
rect 12704 -828 12711 -776
rect 6144 -981 6192 -840
rect 6895 -875 6941 -835
rect 6895 -935 6901 -875
rect 6935 -935 6941 -875
rect 6895 -947 6941 -935
rect 6969 -875 7059 -863
rect 6969 -879 6997 -875
rect 7031 -879 7059 -875
rect 6969 -931 6988 -879
rect 7040 -931 7059 -879
rect 6969 -935 6997 -931
rect 7031 -935 7059 -931
rect 6969 -947 7059 -935
rect 7087 -875 7133 -835
rect 7087 -935 7093 -875
rect 7127 -935 7133 -875
rect 7087 -947 7133 -935
rect 7175 -875 7221 -863
rect 7737 -871 7783 -862
rect 7175 -935 7181 -875
rect 7215 -935 7221 -875
rect 7175 -947 7221 -935
rect 7715 -872 7797 -871
rect 7715 -936 7724 -872
rect 7788 -936 7797 -872
rect 7826 -874 7872 -862
rect 8469 -871 8515 -862
rect 7826 -934 7832 -874
rect 7866 -934 7872 -874
rect 7737 -946 7783 -936
rect 6144 -1028 6812 -981
rect 6909 -985 7091 -979
rect 6909 -1019 7045 -985
rect 7079 -989 7091 -985
rect 7175 -989 7203 -947
rect 7079 -1018 7203 -989
rect 7079 -1019 7091 -1018
rect 6909 -1025 7091 -1019
rect 6144 -1428 6192 -1028
rect 7175 -1066 7203 -1018
rect 7236 -983 7298 -981
rect 7826 -983 7872 -934
rect 8447 -872 8529 -871
rect 8447 -936 8456 -872
rect 8520 -936 8529 -872
rect 8575 -874 8621 -862
rect 8681 -871 8727 -862
rect 9807 -871 9853 -862
rect 8575 -934 8581 -874
rect 8615 -934 8621 -874
rect 8469 -946 8515 -936
rect 8575 -983 8621 -934
rect 8667 -872 8749 -871
rect 8667 -936 8676 -872
rect 8740 -936 8749 -872
rect 9785 -872 9867 -871
rect 9785 -936 9794 -872
rect 9858 -936 9867 -872
rect 9915 -874 9961 -862
rect 10019 -871 10065 -862
rect 11019 -871 11065 -862
rect 9915 -934 9921 -874
rect 9955 -934 9961 -874
rect 8681 -946 8727 -936
rect 9807 -946 9853 -936
rect 9915 -983 9961 -934
rect 10005 -872 10087 -871
rect 10005 -936 10014 -872
rect 10078 -936 10087 -872
rect 10997 -872 11079 -871
rect 10997 -936 11006 -872
rect 11070 -936 11079 -872
rect 11126 -874 11172 -862
rect 11231 -871 11277 -862
rect 11126 -934 11132 -874
rect 11166 -934 11172 -874
rect 10019 -946 10065 -936
rect 11019 -946 11065 -936
rect 11126 -983 11172 -934
rect 11217 -872 11299 -871
rect 11217 -936 11226 -872
rect 11290 -936 11299 -872
rect 11875 -874 11921 -862
rect 11963 -871 12009 -862
rect 11875 -934 11881 -874
rect 11915 -934 11921 -874
rect 11231 -946 11277 -936
rect 11875 -983 11921 -934
rect 11949 -872 12031 -871
rect 11949 -936 11958 -872
rect 12022 -936 12031 -872
rect 11963 -946 12009 -936
rect 12815 -983 12861 -762
rect 7236 -987 12861 -983
rect 7236 -1021 7252 -987
rect 7286 -1021 12861 -987
rect 7236 -1025 12861 -1021
rect 7236 -1027 7302 -1025
rect 6895 -1078 6941 -1066
rect 6327 -1119 6787 -1097
rect 6327 -1128 6389 -1119
rect 6441 -1128 6532 -1119
rect 6584 -1128 6652 -1119
rect 6704 -1128 6787 -1119
rect 6327 -1162 6356 -1128
rect 6441 -1162 6448 -1128
rect 6482 -1162 6532 -1128
rect 6584 -1162 6632 -1128
rect 6704 -1162 6724 -1128
rect 6758 -1162 6787 -1128
rect 6327 -1171 6389 -1162
rect 6441 -1171 6532 -1162
rect 6584 -1171 6652 -1162
rect 6704 -1171 6787 -1162
rect 6327 -1193 6787 -1171
rect 6895 -1138 6901 -1078
rect 6935 -1138 6941 -1078
rect 6895 -1178 6941 -1138
rect 6969 -1078 7059 -1066
rect 6969 -1082 6997 -1078
rect 7031 -1082 7059 -1078
rect 6969 -1134 6988 -1082
rect 7040 -1134 7059 -1082
rect 6969 -1138 6997 -1134
rect 7031 -1138 7059 -1134
rect 6969 -1150 7059 -1138
rect 7087 -1078 7133 -1066
rect 7087 -1138 7093 -1078
rect 7127 -1138 7133 -1078
rect 7087 -1178 7133 -1138
rect 7175 -1078 7221 -1066
rect 7736 -1074 7782 -1063
rect 7175 -1138 7181 -1078
rect 7215 -1138 7221 -1078
rect 7175 -1150 7221 -1138
rect 7713 -1138 7720 -1074
rect 7784 -1138 7792 -1074
rect 7713 -1139 7792 -1138
rect 7843 -1075 7889 -1025
rect 7950 -1074 7996 -1063
rect 8948 -1074 8994 -1063
rect 7843 -1135 7849 -1075
rect 7883 -1135 7889 -1075
rect 7736 -1147 7782 -1139
rect 7843 -1147 7889 -1135
rect 7940 -1138 7948 -1074
rect 8012 -1138 8019 -1074
rect 7940 -1139 8019 -1138
rect 8925 -1138 8932 -1074
rect 8996 -1138 9004 -1074
rect 8925 -1139 9004 -1138
rect 9057 -1075 9103 -1025
rect 9162 -1074 9208 -1063
rect 10160 -1074 10206 -1063
rect 9057 -1135 9063 -1075
rect 9097 -1135 9103 -1075
rect 7950 -1147 7996 -1139
rect 8948 -1147 8994 -1139
rect 9057 -1147 9103 -1135
rect 9152 -1138 9160 -1074
rect 9224 -1138 9231 -1074
rect 9152 -1139 9231 -1138
rect 10137 -1138 10144 -1074
rect 10208 -1138 10216 -1074
rect 10137 -1139 10216 -1138
rect 10270 -1075 10316 -1025
rect 10374 -1074 10420 -1063
rect 11372 -1074 11418 -1063
rect 10270 -1135 10276 -1075
rect 10310 -1135 10316 -1075
rect 9162 -1147 9208 -1139
rect 10160 -1147 10206 -1139
rect 10270 -1147 10316 -1135
rect 10364 -1138 10372 -1074
rect 10436 -1138 10443 -1074
rect 10364 -1139 10443 -1138
rect 11349 -1138 11356 -1074
rect 11420 -1138 11428 -1074
rect 11349 -1139 11428 -1138
rect 11481 -1075 11527 -1025
rect 11586 -1074 11632 -1063
rect 11481 -1135 11487 -1075
rect 11521 -1135 11527 -1075
rect 10374 -1147 10420 -1139
rect 11372 -1147 11418 -1139
rect 11481 -1147 11527 -1135
rect 11576 -1138 11584 -1074
rect 11648 -1138 11655 -1074
rect 11576 -1139 11655 -1138
rect 12230 -1075 12276 -1025
rect 12318 -1074 12364 -1063
rect 12230 -1135 12236 -1075
rect 12270 -1135 12276 -1075
rect 11586 -1147 11632 -1139
rect 12230 -1147 12276 -1135
rect 12308 -1138 12316 -1074
rect 12380 -1138 12387 -1074
rect 12308 -1139 12387 -1138
rect 12318 -1147 12364 -1139
rect 6895 -1207 7133 -1178
rect 12715 -1187 12764 -1183
rect 11749 -1188 12195 -1187
rect 12275 -1188 12764 -1187
rect 7774 -1194 12195 -1188
rect 7087 -1216 7133 -1207
rect 6220 -1271 6269 -1258
rect 6220 -1305 6226 -1271
rect 6260 -1295 6269 -1271
rect 7087 -1276 7093 -1216
rect 7127 -1276 7133 -1216
rect 7087 -1288 7133 -1276
rect 7175 -1216 7221 -1204
rect 7175 -1276 7181 -1216
rect 7215 -1276 7221 -1216
rect 7774 -1228 7786 -1194
rect 7820 -1228 7912 -1194
rect 7946 -1228 8998 -1194
rect 9032 -1228 9124 -1194
rect 9158 -1228 10210 -1194
rect 10244 -1228 10336 -1194
rect 10370 -1228 11422 -1194
rect 11456 -1228 11548 -1194
rect 11582 -1228 12195 -1194
rect 7774 -1234 12195 -1228
rect 12263 -1194 12764 -1188
rect 12263 -1228 12280 -1194
rect 12314 -1196 12764 -1194
rect 12314 -1228 12721 -1196
rect 12263 -1230 12721 -1228
rect 12755 -1230 12764 -1196
rect 12263 -1234 12764 -1230
rect 7175 -1279 7221 -1276
rect 6260 -1305 6354 -1295
rect 6220 -1323 6354 -1305
rect 6221 -1364 6270 -1351
rect 6221 -1398 6227 -1364
rect 6261 -1398 6298 -1364
rect 6221 -1410 6298 -1398
rect 6134 -1434 6192 -1428
rect 6134 -1468 6146 -1434
rect 6180 -1468 6192 -1434
rect 6134 -1474 6192 -1468
rect 6060 -1527 6142 -1515
rect 6060 -1587 6102 -1527
rect 6136 -1587 6142 -1527
rect 6060 -1599 6142 -1587
rect 6184 -1527 6230 -1515
rect 6184 -1587 6190 -1527
rect 6224 -1587 6230 -1527
rect 6270 -1542 6298 -1410
rect 6326 -1467 6354 -1323
rect 7175 -1325 7222 -1279
rect 7057 -1343 7222 -1325
rect 12146 -1281 12195 -1234
rect 12715 -1242 12764 -1234
rect 12716 -1281 12765 -1276
rect 12146 -1289 12765 -1281
rect 12146 -1323 12722 -1289
rect 12756 -1323 12765 -1289
rect 12146 -1328 12765 -1323
rect 12716 -1335 12765 -1328
rect 6391 -1354 6457 -1353
rect 6391 -1406 6397 -1354
rect 6449 -1406 6457 -1354
rect 6666 -1361 6720 -1357
rect 6665 -1364 6720 -1361
rect 6665 -1398 6677 -1364
rect 6711 -1398 6849 -1364
rect 7057 -1395 7076 -1343
rect 7128 -1384 7222 -1343
rect 7128 -1395 7147 -1384
rect 6665 -1401 6720 -1398
rect 6665 -1405 6719 -1401
rect 6391 -1408 6457 -1406
rect 7057 -1411 7147 -1395
rect 6326 -1474 6537 -1467
rect 6326 -1495 6487 -1474
rect 6470 -1508 6487 -1495
rect 6521 -1508 6537 -1474
rect 6470 -1514 6537 -1508
rect 12815 -1515 12861 -1025
rect 12899 -800 12957 -794
rect 12899 -834 12911 -800
rect 12945 -834 12957 -800
rect 13133 -828 13140 -776
rect 13192 -778 13198 -776
rect 13192 -825 13586 -778
rect 13192 -828 13198 -825
rect 13133 -829 13198 -828
rect 12899 -840 12957 -834
rect 12899 -981 12947 -840
rect 12899 -1028 13567 -981
rect 12899 -1428 12947 -1028
rect 13082 -1119 13542 -1097
rect 13082 -1128 13144 -1119
rect 13196 -1128 13287 -1119
rect 13339 -1128 13407 -1119
rect 13459 -1128 13542 -1119
rect 13082 -1162 13111 -1128
rect 13196 -1162 13203 -1128
rect 13237 -1162 13287 -1128
rect 13339 -1162 13387 -1128
rect 13459 -1162 13479 -1128
rect 13513 -1162 13542 -1128
rect 13082 -1171 13144 -1162
rect 13196 -1171 13287 -1162
rect 13339 -1171 13407 -1162
rect 13459 -1171 13542 -1162
rect 13082 -1193 13542 -1171
rect 12975 -1271 13024 -1258
rect 12975 -1305 12981 -1271
rect 13015 -1295 13024 -1271
rect 13015 -1305 13109 -1295
rect 12975 -1323 13109 -1305
rect 12976 -1364 13025 -1351
rect 12976 -1398 12982 -1364
rect 13016 -1398 13053 -1364
rect 12976 -1410 13053 -1398
rect 12889 -1434 12947 -1428
rect 12889 -1468 12901 -1434
rect 12935 -1468 12947 -1434
rect 12889 -1474 12947 -1468
rect 6584 -1529 6642 -1522
rect 6584 -1542 6596 -1529
rect 6270 -1563 6596 -1542
rect 6630 -1563 6642 -1529
rect 6270 -1570 6642 -1563
rect 12815 -1527 12897 -1515
rect 6096 -1665 6142 -1653
rect 6096 -1725 6102 -1665
rect 6136 -1725 6142 -1665
rect 6096 -1803 6142 -1725
rect 6184 -1665 6230 -1587
rect 12815 -1587 12857 -1527
rect 12891 -1587 12897 -1527
rect 12815 -1599 12897 -1587
rect 12939 -1527 12985 -1515
rect 12939 -1587 12945 -1527
rect 12979 -1587 12985 -1527
rect 13025 -1542 13053 -1410
rect 13081 -1467 13109 -1323
rect 13146 -1354 13212 -1353
rect 13146 -1406 13152 -1354
rect 13204 -1406 13212 -1354
rect 13421 -1361 13475 -1357
rect 13420 -1364 13475 -1361
rect 13420 -1398 13432 -1364
rect 13466 -1398 13604 -1364
rect 13420 -1401 13475 -1398
rect 13420 -1405 13474 -1401
rect 13146 -1408 13212 -1406
rect 13081 -1474 13292 -1467
rect 13081 -1495 13242 -1474
rect 13225 -1508 13242 -1495
rect 13276 -1508 13292 -1474
rect 13225 -1514 13292 -1508
rect 13339 -1529 13397 -1522
rect 13339 -1542 13351 -1529
rect 13025 -1563 13351 -1542
rect 13385 -1563 13397 -1529
rect 13025 -1570 13397 -1563
rect 6184 -1725 6190 -1665
rect 6224 -1725 6230 -1665
rect 6184 -1737 6230 -1725
rect 6327 -1664 6787 -1641
rect 6327 -1665 6539 -1664
rect 6327 -1672 6395 -1665
rect 6327 -1706 6356 -1672
rect 6390 -1706 6395 -1672
rect 6327 -1717 6395 -1706
rect 6447 -1672 6539 -1665
rect 6591 -1665 6787 -1664
rect 6591 -1672 6670 -1665
rect 6447 -1706 6448 -1672
rect 6482 -1706 6539 -1672
rect 6591 -1706 6632 -1672
rect 6666 -1706 6670 -1672
rect 6447 -1716 6539 -1706
rect 6591 -1716 6670 -1706
rect 6447 -1717 6670 -1716
rect 6722 -1672 6787 -1665
rect 6722 -1706 6724 -1672
rect 6758 -1706 6787 -1672
rect 6722 -1717 6787 -1706
rect 6327 -1737 6787 -1717
rect 12851 -1665 12897 -1653
rect 12851 -1725 12857 -1665
rect 12891 -1725 12897 -1665
rect 6096 -1863 6102 -1803
rect 6136 -1863 6142 -1803
rect 6096 -1875 6142 -1863
rect 6184 -1803 6230 -1791
rect 6184 -1863 6190 -1803
rect 6224 -1863 6230 -1803
rect 6096 -1941 6142 -1929
rect 6096 -2001 6102 -1941
rect 6136 -2001 6142 -1941
rect 6096 -2079 6142 -2001
rect 6184 -1941 6230 -1863
rect 12851 -1803 12897 -1725
rect 12939 -1665 12985 -1587
rect 12939 -1725 12945 -1665
rect 12979 -1725 12985 -1665
rect 12939 -1737 12985 -1725
rect 13082 -1664 13542 -1641
rect 13082 -1665 13294 -1664
rect 13082 -1672 13150 -1665
rect 13082 -1706 13111 -1672
rect 13145 -1706 13150 -1672
rect 13082 -1717 13150 -1706
rect 13202 -1672 13294 -1665
rect 13346 -1665 13542 -1664
rect 13346 -1672 13425 -1665
rect 13202 -1706 13203 -1672
rect 13237 -1706 13294 -1672
rect 13346 -1706 13387 -1672
rect 13421 -1706 13425 -1672
rect 13202 -1716 13294 -1706
rect 13346 -1716 13425 -1706
rect 13202 -1717 13425 -1716
rect 13477 -1672 13542 -1665
rect 13477 -1706 13479 -1672
rect 13513 -1706 13542 -1672
rect 13477 -1717 13542 -1706
rect 13082 -1737 13542 -1717
rect 12851 -1863 12857 -1803
rect 12891 -1863 12897 -1803
rect 12851 -1875 12897 -1863
rect 12939 -1803 12985 -1791
rect 12939 -1863 12945 -1803
rect 12979 -1863 12985 -1803
rect 6184 -2001 6190 -1941
rect 6224 -2001 6230 -1941
rect 6184 -2013 6230 -2001
rect 12851 -1941 12897 -1929
rect 12851 -2001 12857 -1941
rect 12891 -2001 12897 -1941
rect 6096 -2139 6102 -2079
rect 6136 -2139 6142 -2079
rect 6096 -2151 6142 -2139
rect 6184 -2079 6230 -2067
rect 6184 -2139 6190 -2079
rect 6224 -2139 6230 -2079
rect 6096 -2217 6142 -2205
rect 6096 -2255 6102 -2217
rect 6034 -2270 6102 -2255
rect 6034 -2322 6053 -2270
rect 6136 -2277 6142 -2217
rect 6105 -2311 6142 -2277
rect 6184 -2217 6230 -2139
rect 12851 -2079 12897 -2001
rect 12939 -1941 12985 -1863
rect 12939 -2001 12945 -1941
rect 12979 -2001 12985 -1941
rect 12939 -2013 12985 -2001
rect 12851 -2139 12857 -2079
rect 12891 -2139 12897 -2079
rect 12851 -2151 12897 -2139
rect 12939 -2079 12985 -2067
rect 12939 -2139 12945 -2079
rect 12979 -2139 12985 -2079
rect 6184 -2277 6190 -2217
rect 6224 -2277 6230 -2217
rect 12851 -2217 12897 -2205
rect 12851 -2255 12857 -2217
rect 6184 -2289 6230 -2277
rect 12789 -2270 12857 -2255
rect 6105 -2322 6124 -2311
rect 6034 -2338 6124 -2322
rect 12789 -2322 12808 -2270
rect 12891 -2277 12897 -2217
rect 12860 -2311 12897 -2277
rect 12939 -2217 12985 -2139
rect 12939 -2277 12945 -2217
rect 12979 -2277 12985 -2217
rect 12939 -2289 12985 -2277
rect 12860 -2322 12879 -2311
rect 12789 -2338 12879 -2322
<< via1 >>
rect 744 3225 796 3270
rect 744 3218 747 3225
rect 747 3218 796 3225
rect 7433 3225 7485 3270
rect 7433 3218 7436 3225
rect 7436 3218 7485 3225
rect 127 2613 179 2665
rect 258 2654 310 2664
rect 258 2620 275 2654
rect 275 2620 309 2654
rect 309 2620 310 2654
rect 258 2612 310 2620
rect 402 2613 454 2665
rect 6816 2613 6868 2665
rect 6947 2654 6999 2664
rect 6947 2620 6964 2654
rect 6964 2620 6998 2654
rect 6998 2620 6999 2654
rect 6947 2612 6999 2620
rect 7091 2613 7143 2665
rect 400 2345 452 2354
rect 400 2311 412 2345
rect 412 2311 446 2345
rect 446 2311 452 2345
rect 400 2302 452 2311
rect 145 2110 197 2119
rect 265 2110 317 2119
rect 408 2110 460 2119
rect 145 2076 183 2110
rect 183 2076 197 2110
rect 265 2076 275 2110
rect 275 2076 309 2110
rect 309 2076 317 2110
rect 408 2076 459 2110
rect 459 2076 460 2110
rect 145 2067 197 2076
rect 265 2067 317 2076
rect 408 2067 460 2076
rect 412 1724 464 1776
rect 6476 2291 6528 2343
rect 7089 2345 7141 2354
rect 7089 2311 7101 2345
rect 7101 2311 7135 2345
rect 7135 2311 7141 2345
rect 7089 2302 7141 2311
rect 1224 2083 1288 2086
rect 1224 2023 1246 2083
rect 1246 2023 1280 2083
rect 1280 2023 1288 2083
rect 1224 2022 1288 2023
rect 1956 2083 2020 2086
rect 1956 2023 1978 2083
rect 1978 2023 2012 2083
rect 2012 2023 2020 2083
rect 1956 2022 2020 2023
rect 2184 2083 2248 2086
rect 2184 2023 2192 2083
rect 2192 2023 2226 2083
rect 2226 2023 2248 2083
rect 2184 2022 2248 2023
rect 3168 2083 3232 2086
rect 3168 2023 3190 2083
rect 3190 2023 3224 2083
rect 3224 2023 3232 2083
rect 3168 2022 3232 2023
rect 3396 2083 3460 2086
rect 3396 2023 3404 2083
rect 3404 2023 3438 2083
rect 3438 2023 3460 2083
rect 3396 2022 3460 2023
rect 4380 2083 4444 2086
rect 4380 2023 4402 2083
rect 4402 2023 4436 2083
rect 4436 2023 4444 2083
rect 4380 2022 4444 2023
rect 4608 2083 4672 2086
rect 4608 2023 4616 2083
rect 4616 2023 4650 2083
rect 4650 2023 4672 2083
rect 4608 2022 4672 2023
rect 5592 2083 5656 2086
rect 5592 2023 5614 2083
rect 5614 2023 5648 2083
rect 5648 2023 5656 2083
rect 5592 2022 5656 2023
rect 5820 2083 5884 2086
rect 5820 2023 5828 2083
rect 5828 2023 5862 2083
rect 5862 2023 5884 2083
rect 5820 2022 5884 2023
rect 6564 2030 6573 2082
rect 6573 2030 6607 2082
rect 6607 2030 6616 2082
rect 6834 2110 6886 2119
rect 6954 2110 7006 2119
rect 7097 2110 7149 2119
rect 6834 2076 6872 2110
rect 6872 2076 6886 2110
rect 6954 2076 6964 2110
rect 6964 2076 6998 2110
rect 6998 2076 7006 2110
rect 7097 2076 7148 2110
rect 7148 2076 7149 2110
rect 6834 2067 6886 2076
rect 6954 2067 7006 2076
rect 7097 2067 7149 2076
rect 1582 1882 1646 1884
rect 1582 1822 1601 1882
rect 1601 1822 1635 1882
rect 1635 1822 1646 1882
rect 1582 1820 1646 1822
rect 2314 1882 2378 1884
rect 2314 1822 2333 1882
rect 2333 1822 2367 1882
rect 2367 1822 2378 1882
rect 2314 1820 2378 1822
rect 2534 1882 2598 1884
rect 2534 1822 2545 1882
rect 2545 1822 2579 1882
rect 2579 1822 2598 1882
rect 2534 1820 2598 1822
rect 3526 1882 3590 1884
rect 3526 1822 3545 1882
rect 3545 1822 3579 1882
rect 3579 1822 3590 1882
rect 3526 1820 3590 1822
rect 3746 1882 3810 1884
rect 3746 1822 3757 1882
rect 3757 1822 3791 1882
rect 3791 1822 3810 1882
rect 3746 1820 3810 1822
rect 4864 1882 4928 1884
rect 4864 1822 4883 1882
rect 4883 1822 4917 1882
rect 4917 1822 4928 1882
rect 4864 1820 4928 1822
rect 5084 1882 5148 1884
rect 5084 1822 5095 1882
rect 5095 1822 5129 1882
rect 5129 1822 5148 1882
rect 5084 1820 5148 1822
rect 5816 1882 5880 1884
rect 5816 1822 5827 1882
rect 5827 1822 5861 1882
rect 5861 1822 5880 1882
rect 5816 1820 5880 1822
rect 6564 1827 6573 1879
rect 6573 1827 6607 1879
rect 6607 1827 6616 1879
rect 900 1724 952 1776
rect 730 672 739 692
rect 739 672 773 692
rect 773 672 782 692
rect 730 640 782 672
rect 7101 1724 7153 1776
rect 13165 2291 13217 2343
rect 7913 2083 7977 2086
rect 7913 2023 7935 2083
rect 7935 2023 7969 2083
rect 7969 2023 7977 2083
rect 7913 2022 7977 2023
rect 8645 2083 8709 2086
rect 8645 2023 8667 2083
rect 8667 2023 8701 2083
rect 8701 2023 8709 2083
rect 8645 2022 8709 2023
rect 8873 2083 8937 2086
rect 8873 2023 8881 2083
rect 8881 2023 8915 2083
rect 8915 2023 8937 2083
rect 8873 2022 8937 2023
rect 9857 2083 9921 2086
rect 9857 2023 9879 2083
rect 9879 2023 9913 2083
rect 9913 2023 9921 2083
rect 9857 2022 9921 2023
rect 10085 2083 10149 2086
rect 10085 2023 10093 2083
rect 10093 2023 10127 2083
rect 10127 2023 10149 2083
rect 10085 2022 10149 2023
rect 11069 2083 11133 2086
rect 11069 2023 11091 2083
rect 11091 2023 11125 2083
rect 11125 2023 11133 2083
rect 11069 2022 11133 2023
rect 11297 2083 11361 2086
rect 11297 2023 11305 2083
rect 11305 2023 11339 2083
rect 11339 2023 11361 2083
rect 11297 2022 11361 2023
rect 12281 2083 12345 2086
rect 12281 2023 12303 2083
rect 12303 2023 12337 2083
rect 12337 2023 12345 2083
rect 12281 2022 12345 2023
rect 12509 2083 12573 2086
rect 12509 2023 12517 2083
rect 12517 2023 12551 2083
rect 12551 2023 12573 2083
rect 12509 2022 12573 2023
rect 13253 2030 13262 2082
rect 13262 2030 13296 2082
rect 13296 2030 13305 2082
rect 8271 1882 8335 1884
rect 8271 1822 8290 1882
rect 8290 1822 8324 1882
rect 8324 1822 8335 1882
rect 8271 1820 8335 1822
rect 9003 1882 9067 1884
rect 9003 1822 9022 1882
rect 9022 1822 9056 1882
rect 9056 1822 9067 1882
rect 9003 1820 9067 1822
rect 9223 1882 9287 1884
rect 9223 1822 9234 1882
rect 9234 1822 9268 1882
rect 9268 1822 9287 1882
rect 9223 1820 9287 1822
rect 10215 1882 10279 1884
rect 10215 1822 10234 1882
rect 10234 1822 10268 1882
rect 10268 1822 10279 1882
rect 10215 1820 10279 1822
rect 10435 1882 10499 1884
rect 10435 1822 10446 1882
rect 10446 1822 10480 1882
rect 10480 1822 10499 1882
rect 10435 1820 10499 1822
rect 11553 1882 11617 1884
rect 11553 1822 11572 1882
rect 11572 1822 11606 1882
rect 11606 1822 11617 1882
rect 11553 1820 11617 1822
rect 11773 1882 11837 1884
rect 11773 1822 11784 1882
rect 11784 1822 11818 1882
rect 11818 1822 11837 1882
rect 11773 1820 11837 1822
rect 12505 1882 12569 1884
rect 12505 1822 12516 1882
rect 12516 1822 12550 1882
rect 12550 1822 12569 1882
rect 12505 1820 12569 1822
rect 13253 1827 13262 1879
rect 13262 1827 13296 1879
rect 13296 1827 13305 1879
rect 7589 1724 7641 1776
rect 6473 1565 6525 1617
rect 7419 672 7428 692
rect 7428 672 7462 692
rect 7462 672 7471 692
rect 7419 640 7471 672
rect 13162 1565 13214 1617
rect 324 -669 376 -617
rect 6067 276 6119 308
rect 6067 256 6076 276
rect 6076 256 6110 276
rect 6110 256 6119 276
rect 7079 -669 7131 -617
rect 5897 -828 5949 -776
rect 233 -931 242 -879
rect 242 -931 276 -879
rect 276 -931 285 -879
rect 969 -874 1033 -872
rect 969 -934 988 -874
rect 988 -934 1022 -874
rect 1022 -934 1033 -874
rect 969 -936 1033 -934
rect 1701 -874 1765 -872
rect 1701 -934 1720 -874
rect 1720 -934 1754 -874
rect 1754 -934 1765 -874
rect 1701 -936 1765 -934
rect 1921 -874 1985 -872
rect 1921 -934 1932 -874
rect 1932 -934 1966 -874
rect 1966 -934 1985 -874
rect 1921 -936 1985 -934
rect 3039 -874 3103 -872
rect 3039 -934 3058 -874
rect 3058 -934 3092 -874
rect 3092 -934 3103 -874
rect 3039 -936 3103 -934
rect 3259 -874 3323 -872
rect 3259 -934 3270 -874
rect 3270 -934 3304 -874
rect 3304 -934 3323 -874
rect 3259 -936 3323 -934
rect 4251 -874 4315 -872
rect 4251 -934 4270 -874
rect 4270 -934 4304 -874
rect 4304 -934 4315 -874
rect 4251 -936 4315 -934
rect 4471 -874 4535 -872
rect 4471 -934 4482 -874
rect 4482 -934 4516 -874
rect 4516 -934 4535 -874
rect 4471 -936 4535 -934
rect 5203 -874 5267 -872
rect 5203 -934 5214 -874
rect 5214 -934 5248 -874
rect 5248 -934 5267 -874
rect 5203 -936 5267 -934
rect 233 -1134 242 -1082
rect 242 -1134 276 -1082
rect 276 -1134 285 -1082
rect 965 -1075 1029 -1074
rect 965 -1135 987 -1075
rect 987 -1135 1021 -1075
rect 1021 -1135 1029 -1075
rect 965 -1138 1029 -1135
rect 1193 -1075 1257 -1074
rect 1193 -1135 1201 -1075
rect 1201 -1135 1235 -1075
rect 1235 -1135 1257 -1075
rect 1193 -1138 1257 -1135
rect 2177 -1075 2241 -1074
rect 2177 -1135 2199 -1075
rect 2199 -1135 2233 -1075
rect 2233 -1135 2241 -1075
rect 2177 -1138 2241 -1135
rect 2405 -1075 2469 -1074
rect 2405 -1135 2413 -1075
rect 2413 -1135 2447 -1075
rect 2447 -1135 2469 -1075
rect 2405 -1138 2469 -1135
rect 3389 -1075 3453 -1074
rect 3389 -1135 3411 -1075
rect 3411 -1135 3445 -1075
rect 3445 -1135 3453 -1075
rect 3389 -1138 3453 -1135
rect 3617 -1075 3681 -1074
rect 3617 -1135 3625 -1075
rect 3625 -1135 3659 -1075
rect 3659 -1135 3681 -1075
rect 3617 -1138 3681 -1135
rect 4601 -1075 4665 -1074
rect 4601 -1135 4623 -1075
rect 4623 -1135 4657 -1075
rect 4657 -1135 4665 -1075
rect 4601 -1138 4665 -1135
rect 4829 -1075 4893 -1074
rect 4829 -1135 4837 -1075
rect 4837 -1135 4871 -1075
rect 4871 -1135 4893 -1075
rect 4829 -1138 4893 -1135
rect 5561 -1075 5625 -1074
rect 5561 -1135 5569 -1075
rect 5569 -1135 5603 -1075
rect 5603 -1135 5625 -1075
rect 5561 -1138 5625 -1135
rect 321 -1395 373 -1343
rect 6385 -828 6437 -776
rect 12822 276 12874 308
rect 12822 256 12831 276
rect 12831 256 12865 276
rect 12865 256 12874 276
rect 12652 -828 12704 -776
rect 6988 -931 6997 -879
rect 6997 -931 7031 -879
rect 7031 -931 7040 -879
rect 7724 -874 7788 -872
rect 7724 -934 7743 -874
rect 7743 -934 7777 -874
rect 7777 -934 7788 -874
rect 7724 -936 7788 -934
rect 8456 -874 8520 -872
rect 8456 -934 8475 -874
rect 8475 -934 8509 -874
rect 8509 -934 8520 -874
rect 8456 -936 8520 -934
rect 8676 -874 8740 -872
rect 8676 -934 8687 -874
rect 8687 -934 8721 -874
rect 8721 -934 8740 -874
rect 8676 -936 8740 -934
rect 9794 -874 9858 -872
rect 9794 -934 9813 -874
rect 9813 -934 9847 -874
rect 9847 -934 9858 -874
rect 9794 -936 9858 -934
rect 10014 -874 10078 -872
rect 10014 -934 10025 -874
rect 10025 -934 10059 -874
rect 10059 -934 10078 -874
rect 10014 -936 10078 -934
rect 11006 -874 11070 -872
rect 11006 -934 11025 -874
rect 11025 -934 11059 -874
rect 11059 -934 11070 -874
rect 11006 -936 11070 -934
rect 11226 -874 11290 -872
rect 11226 -934 11237 -874
rect 11237 -934 11271 -874
rect 11271 -934 11290 -874
rect 11226 -936 11290 -934
rect 11958 -874 12022 -872
rect 11958 -934 11969 -874
rect 11969 -934 12003 -874
rect 12003 -934 12022 -874
rect 11958 -936 12022 -934
rect 6389 -1128 6441 -1119
rect 6532 -1128 6584 -1119
rect 6652 -1128 6704 -1119
rect 6389 -1162 6390 -1128
rect 6390 -1162 6441 -1128
rect 6532 -1162 6540 -1128
rect 6540 -1162 6574 -1128
rect 6574 -1162 6584 -1128
rect 6652 -1162 6666 -1128
rect 6666 -1162 6704 -1128
rect 6389 -1171 6441 -1162
rect 6532 -1171 6584 -1162
rect 6652 -1171 6704 -1162
rect 6988 -1134 6997 -1082
rect 6997 -1134 7031 -1082
rect 7031 -1134 7040 -1082
rect 7720 -1075 7784 -1074
rect 7720 -1135 7742 -1075
rect 7742 -1135 7776 -1075
rect 7776 -1135 7784 -1075
rect 7720 -1138 7784 -1135
rect 7948 -1075 8012 -1074
rect 7948 -1135 7956 -1075
rect 7956 -1135 7990 -1075
rect 7990 -1135 8012 -1075
rect 7948 -1138 8012 -1135
rect 8932 -1075 8996 -1074
rect 8932 -1135 8954 -1075
rect 8954 -1135 8988 -1075
rect 8988 -1135 8996 -1075
rect 8932 -1138 8996 -1135
rect 9160 -1075 9224 -1074
rect 9160 -1135 9168 -1075
rect 9168 -1135 9202 -1075
rect 9202 -1135 9224 -1075
rect 9160 -1138 9224 -1135
rect 10144 -1075 10208 -1074
rect 10144 -1135 10166 -1075
rect 10166 -1135 10200 -1075
rect 10200 -1135 10208 -1075
rect 10144 -1138 10208 -1135
rect 10372 -1075 10436 -1074
rect 10372 -1135 10380 -1075
rect 10380 -1135 10414 -1075
rect 10414 -1135 10436 -1075
rect 10372 -1138 10436 -1135
rect 11356 -1075 11420 -1074
rect 11356 -1135 11378 -1075
rect 11378 -1135 11412 -1075
rect 11412 -1135 11420 -1075
rect 11356 -1138 11420 -1135
rect 11584 -1075 11648 -1074
rect 11584 -1135 11592 -1075
rect 11592 -1135 11626 -1075
rect 11626 -1135 11648 -1075
rect 11584 -1138 11648 -1135
rect 12316 -1075 12380 -1074
rect 12316 -1135 12324 -1075
rect 12324 -1135 12358 -1075
rect 12358 -1135 12380 -1075
rect 12316 -1138 12380 -1135
rect 6397 -1363 6449 -1354
rect 6397 -1397 6403 -1363
rect 6403 -1397 6437 -1363
rect 6437 -1397 6449 -1363
rect 6397 -1406 6449 -1397
rect 7076 -1395 7128 -1343
rect 13140 -828 13192 -776
rect 13144 -1128 13196 -1119
rect 13287 -1128 13339 -1119
rect 13407 -1128 13459 -1119
rect 13144 -1162 13145 -1128
rect 13145 -1162 13196 -1128
rect 13287 -1162 13295 -1128
rect 13295 -1162 13329 -1128
rect 13329 -1162 13339 -1128
rect 13407 -1162 13421 -1128
rect 13421 -1162 13459 -1128
rect 13144 -1171 13196 -1162
rect 13287 -1171 13339 -1162
rect 13407 -1171 13459 -1162
rect 13152 -1363 13204 -1354
rect 13152 -1397 13158 -1363
rect 13158 -1397 13192 -1363
rect 13192 -1397 13204 -1363
rect 13152 -1406 13204 -1397
rect 6395 -1717 6447 -1665
rect 6539 -1672 6591 -1664
rect 6539 -1706 6540 -1672
rect 6540 -1706 6574 -1672
rect 6574 -1706 6591 -1672
rect 6539 -1716 6591 -1706
rect 6670 -1717 6722 -1665
rect 13150 -1717 13202 -1665
rect 13294 -1672 13346 -1664
rect 13294 -1706 13295 -1672
rect 13295 -1706 13329 -1672
rect 13329 -1706 13346 -1672
rect 13294 -1716 13346 -1706
rect 13425 -1717 13477 -1665
rect 6053 -2277 6102 -2270
rect 6102 -2277 6105 -2270
rect 6053 -2322 6105 -2277
rect 12808 -2277 12857 -2270
rect 12857 -2277 12860 -2270
rect 12808 -2322 12860 -2277
<< metal2 >>
rect 733 3272 807 3276
rect 733 3216 742 3272
rect 798 3216 807 3272
rect 733 3212 807 3216
rect 7422 3272 7496 3276
rect 7422 3216 7431 3272
rect 7487 3216 7496 3272
rect 7422 3212 7496 3216
rect 125 2667 181 2676
rect 125 2602 181 2611
rect 256 2666 312 2675
rect 256 2601 312 2610
rect 400 2667 456 2676
rect 400 2602 456 2611
rect 6814 2667 6870 2676
rect 6814 2602 6870 2611
rect 6945 2666 7001 2675
rect 6945 2601 7001 2610
rect 7089 2667 7145 2676
rect 7089 2602 7145 2611
rect 392 2302 400 2354
rect 452 2302 458 2354
rect 392 2301 458 2302
rect 6465 2345 6539 2349
rect 410 2225 456 2301
rect 6465 2289 6474 2345
rect 6530 2289 6539 2345
rect 7081 2302 7089 2354
rect 7141 2302 7147 2354
rect 7081 2301 7147 2302
rect 13154 2345 13228 2349
rect 6465 2285 6539 2289
rect 7099 2225 7145 2301
rect 13154 2289 13163 2345
rect 13219 2289 13228 2345
rect 13154 2285 13228 2289
rect 410 2179 649 2225
rect 7099 2179 7338 2225
rect 143 2121 199 2130
rect 143 2056 199 2065
rect 263 2121 319 2130
rect 263 2056 319 2065
rect 406 2121 462 2130
rect 406 2056 462 2065
rect 406 1776 471 1777
rect 406 1724 412 1776
rect 464 1773 471 1776
rect 603 1773 649 2179
rect 6832 2121 6888 2130
rect 1217 2086 1296 2087
rect 1949 2086 2028 2087
rect 2176 2086 2255 2087
rect 3161 2086 3240 2087
rect 3388 2086 3467 2087
rect 4373 2086 4452 2087
rect 4600 2086 4679 2087
rect 5585 2086 5664 2087
rect 5812 2086 5891 2087
rect 1214 2022 1224 2086
rect 1288 2022 1297 2086
rect 1946 2022 1956 2086
rect 2020 2022 2029 2086
rect 2175 2022 2184 2086
rect 2248 2022 2258 2086
rect 3158 2022 3168 2086
rect 3232 2022 3241 2086
rect 3387 2022 3396 2086
rect 3460 2022 3470 2086
rect 4370 2022 4380 2086
rect 4444 2022 4453 2086
rect 4599 2022 4608 2086
rect 4672 2022 4682 2086
rect 5582 2022 5592 2086
rect 5656 2022 5665 2086
rect 5811 2022 5820 2086
rect 5884 2022 5894 2086
rect 6553 2084 6627 2088
rect 6553 2028 6562 2084
rect 6618 2028 6627 2084
rect 6832 2056 6888 2065
rect 6952 2121 7008 2130
rect 6952 2056 7008 2065
rect 7095 2121 7151 2130
rect 7095 2056 7151 2065
rect 6553 2024 6627 2028
rect 1573 1820 1582 1884
rect 1646 1820 1655 1884
rect 1573 1819 1655 1820
rect 2305 1820 2314 1884
rect 2378 1820 2387 1884
rect 2305 1819 2387 1820
rect 2525 1820 2534 1884
rect 2598 1820 2607 1884
rect 2525 1819 2607 1820
rect 3517 1820 3526 1884
rect 3590 1820 3599 1884
rect 3517 1819 3599 1820
rect 3737 1820 3746 1884
rect 3810 1820 3819 1884
rect 3737 1819 3819 1820
rect 4855 1820 4864 1884
rect 4928 1820 4937 1884
rect 4855 1819 4937 1820
rect 5075 1820 5084 1884
rect 5148 1820 5157 1884
rect 5075 1819 5157 1820
rect 5807 1820 5816 1884
rect 5880 1820 5889 1884
rect 6553 1881 6627 1885
rect 6553 1825 6562 1881
rect 6618 1825 6627 1881
rect 6553 1821 6627 1825
rect 5807 1819 5889 1820
rect 7095 1776 7160 1777
rect 893 1773 900 1776
rect 464 1727 900 1773
rect 464 1724 471 1727
rect 893 1724 900 1727
rect 952 1724 958 1776
rect 7095 1724 7101 1776
rect 7153 1773 7160 1776
rect 7292 1773 7338 2179
rect 7906 2086 7985 2087
rect 8638 2086 8717 2087
rect 8865 2086 8944 2087
rect 9850 2086 9929 2087
rect 10077 2086 10156 2087
rect 11062 2086 11141 2087
rect 11289 2086 11368 2087
rect 12274 2086 12353 2087
rect 12501 2086 12580 2087
rect 7903 2022 7913 2086
rect 7977 2022 7986 2086
rect 8635 2022 8645 2086
rect 8709 2022 8718 2086
rect 8864 2022 8873 2086
rect 8937 2022 8947 2086
rect 9847 2022 9857 2086
rect 9921 2022 9930 2086
rect 10076 2022 10085 2086
rect 10149 2022 10159 2086
rect 11059 2022 11069 2086
rect 11133 2022 11142 2086
rect 11288 2022 11297 2086
rect 11361 2022 11371 2086
rect 12271 2022 12281 2086
rect 12345 2022 12354 2086
rect 12500 2022 12509 2086
rect 12573 2022 12583 2086
rect 13242 2084 13316 2088
rect 13242 2028 13251 2084
rect 13307 2028 13316 2084
rect 13242 2024 13316 2028
rect 8262 1820 8271 1884
rect 8335 1820 8344 1884
rect 8262 1819 8344 1820
rect 8994 1820 9003 1884
rect 9067 1820 9076 1884
rect 8994 1819 9076 1820
rect 9214 1820 9223 1884
rect 9287 1820 9296 1884
rect 9214 1819 9296 1820
rect 10206 1820 10215 1884
rect 10279 1820 10288 1884
rect 10206 1819 10288 1820
rect 10426 1820 10435 1884
rect 10499 1820 10508 1884
rect 10426 1819 10508 1820
rect 11544 1820 11553 1884
rect 11617 1820 11626 1884
rect 11544 1819 11626 1820
rect 11764 1820 11773 1884
rect 11837 1820 11846 1884
rect 11764 1819 11846 1820
rect 12496 1820 12505 1884
rect 12569 1820 12578 1884
rect 13242 1881 13316 1885
rect 13242 1825 13251 1881
rect 13307 1825 13316 1881
rect 13242 1821 13316 1825
rect 12496 1819 12578 1820
rect 7582 1773 7589 1776
rect 7153 1727 7589 1773
rect 7153 1724 7160 1727
rect 7582 1724 7589 1727
rect 7641 1724 7647 1776
rect 893 1723 958 1724
rect 7582 1723 7647 1724
rect 6462 1619 6536 1623
rect 6462 1563 6471 1619
rect 6527 1563 6536 1619
rect 6462 1559 6536 1563
rect 13151 1619 13225 1623
rect 13151 1563 13160 1619
rect 13216 1563 13225 1619
rect 13151 1559 13225 1563
rect 719 694 793 698
rect 719 638 728 694
rect 784 638 793 694
rect 719 634 793 638
rect 7408 694 7482 698
rect 7408 638 7417 694
rect 7473 638 7482 694
rect 7408 634 7482 638
rect 6056 310 6130 314
rect 6056 254 6065 310
rect 6121 254 6130 310
rect 6056 250 6130 254
rect 12811 310 12885 314
rect 12811 254 12820 310
rect 12876 254 12885 310
rect 12811 250 12885 254
rect 313 -615 387 -611
rect 313 -671 322 -615
rect 378 -671 387 -615
rect 313 -675 387 -671
rect 7068 -615 7142 -611
rect 7068 -671 7077 -615
rect 7133 -671 7142 -615
rect 7068 -675 7142 -671
rect 5891 -776 5956 -775
rect 12646 -776 12711 -775
rect 5891 -828 5897 -776
rect 5949 -779 5956 -776
rect 6378 -779 6385 -776
rect 5949 -825 6385 -779
rect 5949 -828 5956 -825
rect 960 -872 1042 -871
rect 222 -877 296 -873
rect 222 -933 231 -877
rect 287 -933 296 -877
rect 222 -937 296 -933
rect 960 -936 969 -872
rect 1033 -936 1042 -872
rect 1692 -872 1774 -871
rect 1692 -936 1701 -872
rect 1765 -936 1774 -872
rect 1912 -872 1994 -871
rect 1912 -936 1921 -872
rect 1985 -936 1994 -872
rect 3030 -872 3112 -871
rect 3030 -936 3039 -872
rect 3103 -936 3112 -872
rect 3250 -872 3332 -871
rect 3250 -936 3259 -872
rect 3323 -936 3332 -872
rect 4242 -872 4324 -871
rect 4242 -936 4251 -872
rect 4315 -936 4324 -872
rect 4462 -872 4544 -871
rect 4462 -936 4471 -872
rect 4535 -936 4544 -872
rect 5194 -872 5276 -871
rect 5194 -936 5203 -872
rect 5267 -936 5276 -872
rect 222 -1080 296 -1076
rect 222 -1136 231 -1080
rect 287 -1136 296 -1080
rect 222 -1140 296 -1136
rect 955 -1138 965 -1074
rect 1029 -1138 1038 -1074
rect 1184 -1138 1193 -1074
rect 1257 -1138 1267 -1074
rect 2167 -1138 2177 -1074
rect 2241 -1138 2250 -1074
rect 2396 -1138 2405 -1074
rect 2469 -1138 2479 -1074
rect 3379 -1138 3389 -1074
rect 3453 -1138 3462 -1074
rect 3608 -1138 3617 -1074
rect 3681 -1138 3691 -1074
rect 4591 -1138 4601 -1074
rect 4665 -1138 4674 -1074
rect 4820 -1138 4829 -1074
rect 4893 -1138 4903 -1074
rect 5552 -1138 5561 -1074
rect 5625 -1138 5635 -1074
rect 958 -1139 1037 -1138
rect 1185 -1139 1264 -1138
rect 2170 -1139 2249 -1138
rect 2397 -1139 2476 -1138
rect 3382 -1139 3461 -1138
rect 3609 -1139 3688 -1138
rect 4594 -1139 4673 -1138
rect 4821 -1139 4900 -1138
rect 5553 -1139 5632 -1138
rect 6200 -1231 6246 -825
rect 6378 -828 6385 -825
rect 6437 -828 6443 -776
rect 12646 -828 12652 -776
rect 12704 -779 12711 -776
rect 13133 -779 13140 -776
rect 12704 -825 13140 -779
rect 12704 -828 12711 -825
rect 6378 -829 6443 -828
rect 7715 -872 7797 -871
rect 6977 -877 7051 -873
rect 6977 -933 6986 -877
rect 7042 -933 7051 -877
rect 6977 -937 7051 -933
rect 7715 -936 7724 -872
rect 7788 -936 7797 -872
rect 8447 -872 8529 -871
rect 8447 -936 8456 -872
rect 8520 -936 8529 -872
rect 8667 -872 8749 -871
rect 8667 -936 8676 -872
rect 8740 -936 8749 -872
rect 9785 -872 9867 -871
rect 9785 -936 9794 -872
rect 9858 -936 9867 -872
rect 10005 -872 10087 -871
rect 10005 -936 10014 -872
rect 10078 -936 10087 -872
rect 10997 -872 11079 -871
rect 10997 -936 11006 -872
rect 11070 -936 11079 -872
rect 11217 -872 11299 -871
rect 11217 -936 11226 -872
rect 11290 -936 11299 -872
rect 11949 -872 12031 -871
rect 11949 -936 11958 -872
rect 12022 -936 12031 -872
rect 6977 -1080 7051 -1076
rect 6387 -1117 6443 -1108
rect 6387 -1182 6443 -1173
rect 6530 -1117 6586 -1108
rect 6530 -1182 6586 -1173
rect 6650 -1117 6706 -1108
rect 6977 -1136 6986 -1080
rect 7042 -1136 7051 -1080
rect 6977 -1140 7051 -1136
rect 7710 -1138 7720 -1074
rect 7784 -1138 7793 -1074
rect 7939 -1138 7948 -1074
rect 8012 -1138 8022 -1074
rect 8922 -1138 8932 -1074
rect 8996 -1138 9005 -1074
rect 9151 -1138 9160 -1074
rect 9224 -1138 9234 -1074
rect 10134 -1138 10144 -1074
rect 10208 -1138 10217 -1074
rect 10363 -1138 10372 -1074
rect 10436 -1138 10446 -1074
rect 11346 -1138 11356 -1074
rect 11420 -1138 11429 -1074
rect 11575 -1138 11584 -1074
rect 11648 -1138 11658 -1074
rect 12307 -1138 12316 -1074
rect 12380 -1138 12390 -1074
rect 7713 -1139 7792 -1138
rect 7940 -1139 8019 -1138
rect 8925 -1139 9004 -1138
rect 9152 -1139 9231 -1138
rect 10137 -1139 10216 -1138
rect 10364 -1139 10443 -1138
rect 11349 -1139 11428 -1138
rect 11576 -1139 11655 -1138
rect 12308 -1139 12387 -1138
rect 6650 -1182 6706 -1173
rect 12955 -1231 13001 -825
rect 13133 -828 13140 -825
rect 13192 -828 13198 -776
rect 13133 -829 13198 -828
rect 13142 -1117 13198 -1108
rect 13142 -1182 13198 -1173
rect 13285 -1117 13341 -1108
rect 13285 -1182 13341 -1173
rect 13405 -1117 13461 -1108
rect 13405 -1182 13461 -1173
rect 6200 -1277 6439 -1231
rect 12955 -1277 13194 -1231
rect 310 -1341 384 -1337
rect 310 -1397 319 -1341
rect 375 -1397 384 -1341
rect 6393 -1353 6439 -1277
rect 7065 -1341 7139 -1337
rect 310 -1401 384 -1397
rect 6391 -1354 6457 -1353
rect 6391 -1406 6397 -1354
rect 6449 -1406 6457 -1354
rect 7065 -1397 7074 -1341
rect 7130 -1397 7139 -1341
rect 13148 -1353 13194 -1277
rect 7065 -1401 7139 -1397
rect 13146 -1354 13212 -1353
rect 13146 -1406 13152 -1354
rect 13204 -1406 13212 -1354
rect 6393 -1663 6449 -1654
rect 6393 -1728 6449 -1719
rect 6537 -1662 6593 -1653
rect 6537 -1727 6593 -1718
rect 6668 -1663 6724 -1654
rect 6668 -1728 6724 -1719
rect 13148 -1663 13204 -1654
rect 13148 -1728 13204 -1719
rect 13292 -1662 13348 -1653
rect 13292 -1727 13348 -1718
rect 13423 -1663 13479 -1654
rect 13423 -1728 13479 -1719
rect 6042 -2268 6116 -2264
rect 6042 -2324 6051 -2268
rect 6107 -2324 6116 -2268
rect 6042 -2328 6116 -2324
rect 12797 -2268 12871 -2264
rect 12797 -2324 12806 -2268
rect 12862 -2324 12871 -2268
rect 12797 -2328 12871 -2324
<< via2 >>
rect 742 3270 798 3272
rect 742 3218 744 3270
rect 744 3218 796 3270
rect 796 3218 798 3270
rect 742 3216 798 3218
rect 7431 3270 7487 3272
rect 7431 3218 7433 3270
rect 7433 3218 7485 3270
rect 7485 3218 7487 3270
rect 7431 3216 7487 3218
rect 125 2665 181 2667
rect 125 2613 127 2665
rect 127 2613 179 2665
rect 179 2613 181 2665
rect 125 2611 181 2613
rect 256 2664 312 2666
rect 256 2612 258 2664
rect 258 2612 310 2664
rect 310 2612 312 2664
rect 256 2610 312 2612
rect 400 2665 456 2667
rect 400 2613 402 2665
rect 402 2613 454 2665
rect 454 2613 456 2665
rect 400 2611 456 2613
rect 6814 2665 6870 2667
rect 6814 2613 6816 2665
rect 6816 2613 6868 2665
rect 6868 2613 6870 2665
rect 6814 2611 6870 2613
rect 6945 2664 7001 2666
rect 6945 2612 6947 2664
rect 6947 2612 6999 2664
rect 6999 2612 7001 2664
rect 6945 2610 7001 2612
rect 7089 2665 7145 2667
rect 7089 2613 7091 2665
rect 7091 2613 7143 2665
rect 7143 2613 7145 2665
rect 7089 2611 7145 2613
rect 6474 2343 6530 2345
rect 6474 2291 6476 2343
rect 6476 2291 6528 2343
rect 6528 2291 6530 2343
rect 6474 2289 6530 2291
rect 13163 2343 13219 2345
rect 13163 2291 13165 2343
rect 13165 2291 13217 2343
rect 13217 2291 13219 2343
rect 13163 2289 13219 2291
rect 143 2119 199 2121
rect 143 2067 145 2119
rect 145 2067 197 2119
rect 197 2067 199 2119
rect 143 2065 199 2067
rect 263 2119 319 2121
rect 263 2067 265 2119
rect 265 2067 317 2119
rect 317 2067 319 2119
rect 263 2065 319 2067
rect 406 2119 462 2121
rect 406 2067 408 2119
rect 408 2067 460 2119
rect 460 2067 462 2119
rect 406 2065 462 2067
rect 6832 2119 6888 2121
rect 1224 2022 1288 2086
rect 1956 2022 2020 2086
rect 2184 2022 2248 2086
rect 3168 2022 3232 2086
rect 3396 2022 3460 2086
rect 4380 2022 4444 2086
rect 4608 2022 4672 2086
rect 5592 2022 5656 2086
rect 5820 2022 5884 2086
rect 6562 2082 6618 2084
rect 6562 2030 6564 2082
rect 6564 2030 6616 2082
rect 6616 2030 6618 2082
rect 6562 2028 6618 2030
rect 6832 2067 6834 2119
rect 6834 2067 6886 2119
rect 6886 2067 6888 2119
rect 6832 2065 6888 2067
rect 6952 2119 7008 2121
rect 6952 2067 6954 2119
rect 6954 2067 7006 2119
rect 7006 2067 7008 2119
rect 6952 2065 7008 2067
rect 7095 2119 7151 2121
rect 7095 2067 7097 2119
rect 7097 2067 7149 2119
rect 7149 2067 7151 2119
rect 7095 2065 7151 2067
rect 1582 1820 1646 1884
rect 2314 1820 2378 1884
rect 2534 1820 2598 1884
rect 3526 1820 3590 1884
rect 3746 1820 3810 1884
rect 4864 1820 4928 1884
rect 5084 1820 5148 1884
rect 5816 1820 5880 1884
rect 6562 1879 6618 1881
rect 6562 1827 6564 1879
rect 6564 1827 6616 1879
rect 6616 1827 6618 1879
rect 6562 1825 6618 1827
rect 7913 2022 7977 2086
rect 8645 2022 8709 2086
rect 8873 2022 8937 2086
rect 9857 2022 9921 2086
rect 10085 2022 10149 2086
rect 11069 2022 11133 2086
rect 11297 2022 11361 2086
rect 12281 2022 12345 2086
rect 12509 2022 12573 2086
rect 13251 2082 13307 2084
rect 13251 2030 13253 2082
rect 13253 2030 13305 2082
rect 13305 2030 13307 2082
rect 13251 2028 13307 2030
rect 8271 1820 8335 1884
rect 9003 1820 9067 1884
rect 9223 1820 9287 1884
rect 10215 1820 10279 1884
rect 10435 1820 10499 1884
rect 11553 1820 11617 1884
rect 11773 1820 11837 1884
rect 12505 1820 12569 1884
rect 13251 1879 13307 1881
rect 13251 1827 13253 1879
rect 13253 1827 13305 1879
rect 13305 1827 13307 1879
rect 13251 1825 13307 1827
rect 6471 1617 6527 1619
rect 6471 1565 6473 1617
rect 6473 1565 6525 1617
rect 6525 1565 6527 1617
rect 6471 1563 6527 1565
rect 13160 1617 13216 1619
rect 13160 1565 13162 1617
rect 13162 1565 13214 1617
rect 13214 1565 13216 1617
rect 13160 1563 13216 1565
rect 728 692 784 694
rect 728 640 730 692
rect 730 640 782 692
rect 782 640 784 692
rect 728 638 784 640
rect 7417 692 7473 694
rect 7417 640 7419 692
rect 7419 640 7471 692
rect 7471 640 7473 692
rect 7417 638 7473 640
rect 6065 308 6121 310
rect 6065 256 6067 308
rect 6067 256 6119 308
rect 6119 256 6121 308
rect 6065 254 6121 256
rect 12820 308 12876 310
rect 12820 256 12822 308
rect 12822 256 12874 308
rect 12874 256 12876 308
rect 12820 254 12876 256
rect 322 -617 378 -615
rect 322 -669 324 -617
rect 324 -669 376 -617
rect 376 -669 378 -617
rect 322 -671 378 -669
rect 7077 -617 7133 -615
rect 7077 -669 7079 -617
rect 7079 -669 7131 -617
rect 7131 -669 7133 -617
rect 7077 -671 7133 -669
rect 231 -879 287 -877
rect 231 -931 233 -879
rect 233 -931 285 -879
rect 285 -931 287 -879
rect 231 -933 287 -931
rect 969 -936 1033 -872
rect 1701 -936 1765 -872
rect 1921 -936 1985 -872
rect 3039 -936 3103 -872
rect 3259 -936 3323 -872
rect 4251 -936 4315 -872
rect 4471 -936 4535 -872
rect 5203 -936 5267 -872
rect 231 -1082 287 -1080
rect 231 -1134 233 -1082
rect 233 -1134 285 -1082
rect 285 -1134 287 -1082
rect 231 -1136 287 -1134
rect 965 -1138 1029 -1074
rect 1193 -1138 1257 -1074
rect 2177 -1138 2241 -1074
rect 2405 -1138 2469 -1074
rect 3389 -1138 3453 -1074
rect 3617 -1138 3681 -1074
rect 4601 -1138 4665 -1074
rect 4829 -1138 4893 -1074
rect 5561 -1138 5625 -1074
rect 6986 -879 7042 -877
rect 6986 -931 6988 -879
rect 6988 -931 7040 -879
rect 7040 -931 7042 -879
rect 6986 -933 7042 -931
rect 7724 -936 7788 -872
rect 8456 -936 8520 -872
rect 8676 -936 8740 -872
rect 9794 -936 9858 -872
rect 10014 -936 10078 -872
rect 11006 -936 11070 -872
rect 11226 -936 11290 -872
rect 11958 -936 12022 -872
rect 6387 -1119 6443 -1117
rect 6387 -1171 6389 -1119
rect 6389 -1171 6441 -1119
rect 6441 -1171 6443 -1119
rect 6387 -1173 6443 -1171
rect 6530 -1119 6586 -1117
rect 6530 -1171 6532 -1119
rect 6532 -1171 6584 -1119
rect 6584 -1171 6586 -1119
rect 6530 -1173 6586 -1171
rect 6650 -1119 6706 -1117
rect 6650 -1171 6652 -1119
rect 6652 -1171 6704 -1119
rect 6704 -1171 6706 -1119
rect 6986 -1082 7042 -1080
rect 6986 -1134 6988 -1082
rect 6988 -1134 7040 -1082
rect 7040 -1134 7042 -1082
rect 6986 -1136 7042 -1134
rect 7720 -1138 7784 -1074
rect 7948 -1138 8012 -1074
rect 8932 -1138 8996 -1074
rect 9160 -1138 9224 -1074
rect 10144 -1138 10208 -1074
rect 10372 -1138 10436 -1074
rect 11356 -1138 11420 -1074
rect 11584 -1138 11648 -1074
rect 12316 -1138 12380 -1074
rect 6650 -1173 6706 -1171
rect 13142 -1119 13198 -1117
rect 13142 -1171 13144 -1119
rect 13144 -1171 13196 -1119
rect 13196 -1171 13198 -1119
rect 13142 -1173 13198 -1171
rect 13285 -1119 13341 -1117
rect 13285 -1171 13287 -1119
rect 13287 -1171 13339 -1119
rect 13339 -1171 13341 -1119
rect 13285 -1173 13341 -1171
rect 13405 -1119 13461 -1117
rect 13405 -1171 13407 -1119
rect 13407 -1171 13459 -1119
rect 13459 -1171 13461 -1119
rect 13405 -1173 13461 -1171
rect 319 -1343 375 -1341
rect 319 -1395 321 -1343
rect 321 -1395 373 -1343
rect 373 -1395 375 -1343
rect 319 -1397 375 -1395
rect 7074 -1343 7130 -1341
rect 7074 -1395 7076 -1343
rect 7076 -1395 7128 -1343
rect 7128 -1395 7130 -1343
rect 7074 -1397 7130 -1395
rect 6393 -1665 6449 -1663
rect 6393 -1717 6395 -1665
rect 6395 -1717 6447 -1665
rect 6447 -1717 6449 -1665
rect 6393 -1719 6449 -1717
rect 6537 -1664 6593 -1662
rect 6537 -1716 6539 -1664
rect 6539 -1716 6591 -1664
rect 6591 -1716 6593 -1664
rect 6537 -1718 6593 -1716
rect 6668 -1665 6724 -1663
rect 6668 -1717 6670 -1665
rect 6670 -1717 6722 -1665
rect 6722 -1717 6724 -1665
rect 6668 -1719 6724 -1717
rect 13148 -1665 13204 -1663
rect 13148 -1717 13150 -1665
rect 13150 -1717 13202 -1665
rect 13202 -1717 13204 -1665
rect 13148 -1719 13204 -1717
rect 13292 -1664 13348 -1662
rect 13292 -1716 13294 -1664
rect 13294 -1716 13346 -1664
rect 13346 -1716 13348 -1664
rect 13292 -1718 13348 -1716
rect 13423 -1665 13479 -1663
rect 13423 -1717 13425 -1665
rect 13425 -1717 13477 -1665
rect 13477 -1717 13479 -1665
rect 13423 -1719 13479 -1717
rect 6051 -2270 6107 -2268
rect 6051 -2322 6053 -2270
rect 6053 -2322 6105 -2270
rect 6105 -2322 6107 -2270
rect 6051 -2324 6107 -2322
rect 12806 -2270 12862 -2268
rect 12806 -2322 12808 -2270
rect 12808 -2322 12860 -2270
rect 12860 -2322 12862 -2270
rect 12806 -2324 12862 -2322
<< metal3 >>
rect 707 3276 833 3286
rect 707 3212 738 3276
rect 802 3271 833 3276
rect 7396 3276 7522 3286
rect 802 3269 1403 3271
rect 802 3212 835 3269
rect 707 3205 835 3212
rect 899 3205 915 3269
rect 979 3205 995 3269
rect 1059 3205 1075 3269
rect 1139 3205 1155 3269
rect 1219 3205 1235 3269
rect 1299 3205 1403 3269
rect 707 3203 1403 3205
rect 1463 3269 6377 3271
rect 1463 3205 1567 3269
rect 1631 3205 1647 3269
rect 1711 3205 1727 3269
rect 1791 3205 1807 3269
rect 1871 3205 1887 3269
rect 1951 3205 1967 3269
rect 2031 3205 2173 3269
rect 2237 3205 2253 3269
rect 2317 3205 2333 3269
rect 2397 3205 2413 3269
rect 2477 3205 2493 3269
rect 2557 3205 2573 3269
rect 2637 3205 2779 3269
rect 2843 3205 2859 3269
rect 2923 3205 2939 3269
rect 3003 3205 3019 3269
rect 3083 3205 3099 3269
rect 3163 3205 3179 3269
rect 3243 3205 3385 3269
rect 3449 3205 3465 3269
rect 3529 3205 3545 3269
rect 3609 3205 3625 3269
rect 3689 3205 3705 3269
rect 3769 3205 3785 3269
rect 3849 3205 3991 3269
rect 4055 3205 4071 3269
rect 4135 3205 4151 3269
rect 4215 3205 4231 3269
rect 4295 3205 4311 3269
rect 4375 3205 4391 3269
rect 4455 3205 4597 3269
rect 4661 3205 4677 3269
rect 4741 3205 4757 3269
rect 4821 3205 4837 3269
rect 4901 3205 4917 3269
rect 4981 3205 4997 3269
rect 5061 3205 5203 3269
rect 5267 3205 5283 3269
rect 5347 3205 5363 3269
rect 5427 3205 5443 3269
rect 5507 3205 5523 3269
rect 5587 3205 5603 3269
rect 5667 3205 5809 3269
rect 5873 3205 5889 3269
rect 5953 3205 5969 3269
rect 6033 3205 6049 3269
rect 6113 3205 6129 3269
rect 6193 3205 6209 3269
rect 6273 3205 6377 3269
rect 1463 3203 6377 3205
rect 7396 3212 7427 3276
rect 7491 3271 7522 3276
rect 7491 3269 8092 3271
rect 7491 3212 7524 3269
rect 7396 3205 7524 3212
rect 7588 3205 7604 3269
rect 7668 3205 7684 3269
rect 7748 3205 7764 3269
rect 7828 3205 7844 3269
rect 7908 3205 7924 3269
rect 7988 3205 8092 3269
rect 7396 3203 8092 3205
rect 8152 3269 13066 3271
rect 8152 3205 8256 3269
rect 8320 3205 8336 3269
rect 8400 3205 8416 3269
rect 8480 3205 8496 3269
rect 8560 3205 8576 3269
rect 8640 3205 8656 3269
rect 8720 3205 8862 3269
rect 8926 3205 8942 3269
rect 9006 3205 9022 3269
rect 9086 3205 9102 3269
rect 9166 3205 9182 3269
rect 9246 3205 9262 3269
rect 9326 3205 9468 3269
rect 9532 3205 9548 3269
rect 9612 3205 9628 3269
rect 9692 3205 9708 3269
rect 9772 3205 9788 3269
rect 9852 3205 9868 3269
rect 9932 3205 10074 3269
rect 10138 3205 10154 3269
rect 10218 3205 10234 3269
rect 10298 3205 10314 3269
rect 10378 3205 10394 3269
rect 10458 3205 10474 3269
rect 10538 3205 10680 3269
rect 10744 3205 10760 3269
rect 10824 3205 10840 3269
rect 10904 3205 10920 3269
rect 10984 3205 11000 3269
rect 11064 3205 11080 3269
rect 11144 3205 11286 3269
rect 11350 3205 11366 3269
rect 11430 3205 11446 3269
rect 11510 3205 11526 3269
rect 11590 3205 11606 3269
rect 11670 3205 11686 3269
rect 11750 3205 11892 3269
rect 11956 3205 11972 3269
rect 12036 3205 12052 3269
rect 12116 3205 12132 3269
rect 12196 3205 12212 3269
rect 12276 3205 12292 3269
rect 12356 3205 12498 3269
rect 12562 3205 12578 3269
rect 12642 3205 12658 3269
rect 12722 3205 12738 3269
rect 12802 3205 12818 3269
rect 12882 3205 12898 3269
rect 12962 3205 13066 3269
rect 8152 3203 13066 3205
rect 731 3049 797 3139
rect 731 2985 732 3049
rect 796 2985 797 3049
rect 731 2969 797 2985
rect 731 2905 732 2969
rect 796 2905 797 2969
rect 731 2889 797 2905
rect 731 2825 732 2889
rect 796 2825 797 2889
rect 731 2809 797 2825
rect 731 2745 732 2809
rect 796 2745 797 2809
rect 731 2729 797 2745
rect 80 2685 224 2686
rect 355 2685 499 2686
rect 80 2671 499 2685
rect 80 2607 121 2671
rect 185 2670 396 2671
rect 185 2607 252 2670
rect 80 2606 252 2607
rect 316 2607 396 2670
rect 460 2607 499 2671
rect 316 2606 499 2607
rect 80 2590 499 2606
rect 731 2665 732 2729
rect 796 2665 797 2729
rect 731 2649 797 2665
rect 211 2589 355 2590
rect 731 2585 732 2649
rect 796 2585 797 2649
rect 731 2569 797 2585
rect 731 2505 732 2569
rect 796 2505 797 2569
rect 731 2489 797 2505
rect 731 2425 732 2489
rect 796 2425 797 2489
rect 731 2409 797 2425
rect 731 2345 732 2409
rect 796 2345 797 2409
rect 731 2329 797 2345
rect 731 2265 732 2329
rect 796 2265 797 2329
rect 246 2140 338 2141
rect 98 2125 505 2140
rect 98 2061 139 2125
rect 203 2061 259 2125
rect 323 2061 402 2125
rect 466 2061 505 2125
rect 98 2044 505 2061
rect 731 2111 797 2265
rect 857 2111 917 3143
rect 977 2173 1037 3203
rect 1097 2111 1157 3143
rect 1217 2173 1277 3203
rect 1337 3049 1403 3139
rect 1337 2985 1338 3049
rect 1402 2985 1403 3049
rect 1337 2969 1403 2985
rect 1337 2905 1338 2969
rect 1402 2905 1403 2969
rect 1337 2889 1403 2905
rect 1337 2825 1338 2889
rect 1402 2825 1403 2889
rect 1337 2809 1403 2825
rect 1337 2745 1338 2809
rect 1402 2745 1403 2809
rect 1337 2729 1403 2745
rect 1337 2665 1338 2729
rect 1402 2665 1403 2729
rect 1337 2649 1403 2665
rect 1337 2585 1338 2649
rect 1402 2585 1403 2649
rect 1337 2569 1403 2585
rect 1337 2505 1338 2569
rect 1402 2505 1403 2569
rect 1337 2489 1403 2505
rect 1337 2425 1338 2489
rect 1402 2425 1403 2489
rect 1337 2409 1403 2425
rect 1337 2345 1338 2409
rect 1402 2345 1403 2409
rect 1337 2329 1403 2345
rect 1337 2265 1338 2329
rect 1402 2265 1403 2329
rect 1337 2111 1403 2265
rect 731 2109 1403 2111
rect 731 2045 835 2109
rect 899 2045 915 2109
rect 979 2045 995 2109
rect 1059 2045 1075 2109
rect 1139 2045 1155 2109
rect 1219 2086 1235 2109
rect 1219 2045 1224 2086
rect 1299 2045 1403 2109
rect 731 2043 1224 2045
rect 1214 2022 1224 2043
rect 1288 2043 1403 2045
rect 1463 3049 1529 3139
rect 1463 2985 1464 3049
rect 1528 2985 1529 3049
rect 1463 2969 1529 2985
rect 1463 2905 1464 2969
rect 1528 2905 1529 2969
rect 1463 2889 1529 2905
rect 1463 2825 1464 2889
rect 1528 2825 1529 2889
rect 1463 2809 1529 2825
rect 1463 2745 1464 2809
rect 1528 2745 1529 2809
rect 1463 2729 1529 2745
rect 1463 2665 1464 2729
rect 1528 2665 1529 2729
rect 1463 2649 1529 2665
rect 1463 2585 1464 2649
rect 1528 2585 1529 2649
rect 1463 2569 1529 2585
rect 1463 2505 1464 2569
rect 1528 2505 1529 2569
rect 1463 2489 1529 2505
rect 1463 2425 1464 2489
rect 1528 2425 1529 2489
rect 1463 2409 1529 2425
rect 1463 2345 1464 2409
rect 1528 2345 1529 2409
rect 1463 2329 1529 2345
rect 1463 2265 1464 2329
rect 1528 2265 1529 2329
rect 1463 2111 1529 2265
rect 1589 2111 1649 3143
rect 1709 2173 1769 3203
rect 1829 2111 1889 3143
rect 1949 2173 2009 3203
rect 2069 3049 2135 3139
rect 2069 2985 2070 3049
rect 2134 2985 2135 3049
rect 2069 2969 2135 2985
rect 2069 2905 2070 2969
rect 2134 2905 2135 2969
rect 2069 2889 2135 2905
rect 2069 2825 2070 2889
rect 2134 2825 2135 2889
rect 2069 2809 2135 2825
rect 2069 2745 2070 2809
rect 2134 2745 2135 2809
rect 2069 2729 2135 2745
rect 2069 2665 2070 2729
rect 2134 2665 2135 2729
rect 2069 2649 2135 2665
rect 2069 2585 2070 2649
rect 2134 2585 2135 2649
rect 2069 2569 2135 2585
rect 2069 2505 2070 2569
rect 2134 2505 2135 2569
rect 2069 2489 2135 2505
rect 2069 2425 2070 2489
rect 2134 2425 2135 2489
rect 2069 2409 2135 2425
rect 2069 2345 2070 2409
rect 2134 2345 2135 2409
rect 2069 2329 2135 2345
rect 2069 2265 2070 2329
rect 2134 2265 2135 2329
rect 2069 2111 2135 2265
rect 2195 2173 2255 3203
rect 2315 2111 2375 3143
rect 2435 2173 2495 3203
rect 2555 2111 2615 3143
rect 2675 3049 2741 3139
rect 2675 2985 2676 3049
rect 2740 2985 2741 3049
rect 2675 2969 2741 2985
rect 2675 2905 2676 2969
rect 2740 2905 2741 2969
rect 2675 2889 2741 2905
rect 2675 2825 2676 2889
rect 2740 2825 2741 2889
rect 2675 2809 2741 2825
rect 2675 2745 2676 2809
rect 2740 2745 2741 2809
rect 2675 2729 2741 2745
rect 2675 2665 2676 2729
rect 2740 2665 2741 2729
rect 2675 2649 2741 2665
rect 2675 2585 2676 2649
rect 2740 2585 2741 2649
rect 2675 2569 2741 2585
rect 2675 2505 2676 2569
rect 2740 2505 2741 2569
rect 2675 2489 2741 2505
rect 2675 2425 2676 2489
rect 2740 2425 2741 2489
rect 2675 2409 2741 2425
rect 2675 2345 2676 2409
rect 2740 2345 2741 2409
rect 2675 2329 2741 2345
rect 2675 2265 2676 2329
rect 2740 2265 2741 2329
rect 2675 2111 2741 2265
rect 2801 2111 2861 3143
rect 2921 2173 2981 3203
rect 3041 2111 3101 3143
rect 3161 2173 3221 3203
rect 3281 3049 3347 3139
rect 3281 2985 3282 3049
rect 3346 2985 3347 3049
rect 3281 2969 3347 2985
rect 3281 2905 3282 2969
rect 3346 2905 3347 2969
rect 3281 2889 3347 2905
rect 3281 2825 3282 2889
rect 3346 2825 3347 2889
rect 3281 2809 3347 2825
rect 3281 2745 3282 2809
rect 3346 2745 3347 2809
rect 3281 2729 3347 2745
rect 3281 2665 3282 2729
rect 3346 2665 3347 2729
rect 3281 2649 3347 2665
rect 3281 2585 3282 2649
rect 3346 2585 3347 2649
rect 3281 2569 3347 2585
rect 3281 2505 3282 2569
rect 3346 2505 3347 2569
rect 3281 2489 3347 2505
rect 3281 2425 3282 2489
rect 3346 2425 3347 2489
rect 3281 2409 3347 2425
rect 3281 2345 3282 2409
rect 3346 2345 3347 2409
rect 3281 2329 3347 2345
rect 3281 2265 3282 2329
rect 3346 2265 3347 2329
rect 3281 2111 3347 2265
rect 3407 2173 3467 3203
rect 3527 2111 3587 3143
rect 3647 2173 3707 3203
rect 3767 2111 3827 3143
rect 3887 3049 3953 3139
rect 3887 2985 3888 3049
rect 3952 2985 3953 3049
rect 3887 2969 3953 2985
rect 3887 2905 3888 2969
rect 3952 2905 3953 2969
rect 3887 2889 3953 2905
rect 3887 2825 3888 2889
rect 3952 2825 3953 2889
rect 3887 2809 3953 2825
rect 3887 2745 3888 2809
rect 3952 2745 3953 2809
rect 3887 2729 3953 2745
rect 3887 2665 3888 2729
rect 3952 2665 3953 2729
rect 3887 2649 3953 2665
rect 3887 2585 3888 2649
rect 3952 2585 3953 2649
rect 3887 2569 3953 2585
rect 3887 2505 3888 2569
rect 3952 2505 3953 2569
rect 3887 2489 3953 2505
rect 3887 2425 3888 2489
rect 3952 2425 3953 2489
rect 3887 2409 3953 2425
rect 3887 2345 3888 2409
rect 3952 2345 3953 2409
rect 3887 2329 3953 2345
rect 3887 2265 3888 2329
rect 3952 2265 3953 2329
rect 3887 2111 3953 2265
rect 4013 2111 4073 3143
rect 4133 2173 4193 3203
rect 4253 2111 4313 3143
rect 4373 2173 4433 3203
rect 4493 3049 4559 3139
rect 4493 2985 4494 3049
rect 4558 2985 4559 3049
rect 4493 2969 4559 2985
rect 4493 2905 4494 2969
rect 4558 2905 4559 2969
rect 4493 2889 4559 2905
rect 4493 2825 4494 2889
rect 4558 2825 4559 2889
rect 4493 2809 4559 2825
rect 4493 2745 4494 2809
rect 4558 2745 4559 2809
rect 4493 2729 4559 2745
rect 4493 2665 4494 2729
rect 4558 2665 4559 2729
rect 4493 2649 4559 2665
rect 4493 2585 4494 2649
rect 4558 2585 4559 2649
rect 4493 2569 4559 2585
rect 4493 2505 4494 2569
rect 4558 2505 4559 2569
rect 4493 2489 4559 2505
rect 4493 2425 4494 2489
rect 4558 2425 4559 2489
rect 4493 2409 4559 2425
rect 4493 2345 4494 2409
rect 4558 2345 4559 2409
rect 4493 2329 4559 2345
rect 4493 2265 4494 2329
rect 4558 2265 4559 2329
rect 4493 2111 4559 2265
rect 4619 2173 4679 3203
rect 4739 2111 4799 3143
rect 4859 2173 4919 3203
rect 4979 2111 5039 3143
rect 5099 3049 5165 3139
rect 5099 2985 5100 3049
rect 5164 2985 5165 3049
rect 5099 2969 5165 2985
rect 5099 2905 5100 2969
rect 5164 2905 5165 2969
rect 5099 2889 5165 2905
rect 5099 2825 5100 2889
rect 5164 2825 5165 2889
rect 5099 2809 5165 2825
rect 5099 2745 5100 2809
rect 5164 2745 5165 2809
rect 5099 2729 5165 2745
rect 5099 2665 5100 2729
rect 5164 2665 5165 2729
rect 5099 2649 5165 2665
rect 5099 2585 5100 2649
rect 5164 2585 5165 2649
rect 5099 2569 5165 2585
rect 5099 2505 5100 2569
rect 5164 2505 5165 2569
rect 5099 2489 5165 2505
rect 5099 2425 5100 2489
rect 5164 2425 5165 2489
rect 5099 2409 5165 2425
rect 5099 2345 5100 2409
rect 5164 2345 5165 2409
rect 5099 2329 5165 2345
rect 5099 2265 5100 2329
rect 5164 2265 5165 2329
rect 5099 2111 5165 2265
rect 5225 2111 5285 3143
rect 5345 2173 5405 3203
rect 5465 2111 5525 3143
rect 5585 2173 5645 3203
rect 5705 3049 5771 3139
rect 5705 2985 5706 3049
rect 5770 2985 5771 3049
rect 5705 2969 5771 2985
rect 5705 2905 5706 2969
rect 5770 2905 5771 2969
rect 5705 2889 5771 2905
rect 5705 2825 5706 2889
rect 5770 2825 5771 2889
rect 5705 2809 5771 2825
rect 5705 2745 5706 2809
rect 5770 2745 5771 2809
rect 5705 2729 5771 2745
rect 5705 2665 5706 2729
rect 5770 2665 5771 2729
rect 5705 2649 5771 2665
rect 5705 2585 5706 2649
rect 5770 2585 5771 2649
rect 5705 2569 5771 2585
rect 5705 2505 5706 2569
rect 5770 2505 5771 2569
rect 5705 2489 5771 2505
rect 5705 2425 5706 2489
rect 5770 2425 5771 2489
rect 5705 2409 5771 2425
rect 5705 2345 5706 2409
rect 5770 2345 5771 2409
rect 5705 2329 5771 2345
rect 5705 2265 5706 2329
rect 5770 2265 5771 2329
rect 5705 2111 5771 2265
rect 5831 2173 5891 3203
rect 5951 2111 6011 3143
rect 6071 2173 6131 3203
rect 6191 2111 6251 3143
rect 6311 3049 6377 3139
rect 6311 2985 6312 3049
rect 6376 2985 6377 3049
rect 6311 2969 6377 2985
rect 6311 2905 6312 2969
rect 6376 2905 6377 2969
rect 6311 2889 6377 2905
rect 6311 2825 6312 2889
rect 6376 2825 6377 2889
rect 6311 2809 6377 2825
rect 6311 2745 6312 2809
rect 6376 2745 6377 2809
rect 6311 2729 6377 2745
rect 6311 2665 6312 2729
rect 6376 2665 6377 2729
rect 7420 3049 7486 3139
rect 7420 2985 7421 3049
rect 7485 2985 7486 3049
rect 7420 2969 7486 2985
rect 7420 2905 7421 2969
rect 7485 2905 7486 2969
rect 7420 2889 7486 2905
rect 7420 2825 7421 2889
rect 7485 2825 7486 2889
rect 7420 2809 7486 2825
rect 7420 2745 7421 2809
rect 7485 2745 7486 2809
rect 7420 2729 7486 2745
rect 6311 2649 6377 2665
rect 6311 2585 6312 2649
rect 6376 2585 6377 2649
rect 6769 2685 6913 2686
rect 7044 2685 7188 2686
rect 6769 2671 7188 2685
rect 6769 2607 6810 2671
rect 6874 2670 7085 2671
rect 6874 2607 6941 2670
rect 6769 2606 6941 2607
rect 7005 2607 7085 2670
rect 7149 2607 7188 2671
rect 7005 2606 7188 2607
rect 6769 2590 7188 2606
rect 7420 2665 7421 2729
rect 7485 2665 7486 2729
rect 7420 2649 7486 2665
rect 6900 2589 7044 2590
rect 6311 2569 6377 2585
rect 6311 2505 6312 2569
rect 6376 2505 6377 2569
rect 6311 2489 6377 2505
rect 6311 2425 6312 2489
rect 6376 2425 6377 2489
rect 6311 2409 6377 2425
rect 6311 2345 6312 2409
rect 6376 2345 6377 2409
rect 7420 2585 7421 2649
rect 7485 2585 7486 2649
rect 7420 2569 7486 2585
rect 7420 2505 7421 2569
rect 7485 2505 7486 2569
rect 7420 2489 7486 2505
rect 7420 2425 7421 2489
rect 7485 2425 7486 2489
rect 7420 2409 7486 2425
rect 6311 2329 6377 2345
rect 6311 2265 6312 2329
rect 6376 2265 6377 2329
rect 6439 2349 6565 2359
rect 6439 2285 6470 2349
rect 6534 2285 6565 2349
rect 6439 2275 6565 2285
rect 7420 2345 7421 2409
rect 7485 2345 7486 2409
rect 7420 2329 7486 2345
rect 6311 2111 6377 2265
rect 7420 2265 7421 2329
rect 7485 2265 7486 2329
rect 6935 2140 7027 2141
rect 1463 2109 6377 2111
rect 1463 2045 1567 2109
rect 1631 2045 1647 2109
rect 1711 2045 1727 2109
rect 1791 2045 1807 2109
rect 1871 2045 1887 2109
rect 1951 2086 1967 2109
rect 1951 2045 1956 2086
rect 2031 2045 2173 2109
rect 2237 2086 2253 2109
rect 2248 2045 2253 2086
rect 2317 2045 2333 2109
rect 2397 2045 2413 2109
rect 2477 2045 2493 2109
rect 2557 2045 2573 2109
rect 2637 2045 2779 2109
rect 2843 2045 2859 2109
rect 2923 2045 2939 2109
rect 3003 2045 3019 2109
rect 3083 2045 3099 2109
rect 3163 2086 3179 2109
rect 3163 2045 3168 2086
rect 3243 2045 3385 2109
rect 3449 2086 3465 2109
rect 3460 2045 3465 2086
rect 3529 2045 3545 2109
rect 3609 2045 3625 2109
rect 3689 2045 3705 2109
rect 3769 2045 3785 2109
rect 3849 2045 3991 2109
rect 4055 2045 4071 2109
rect 4135 2045 4151 2109
rect 4215 2045 4231 2109
rect 4295 2045 4311 2109
rect 4375 2086 4391 2109
rect 4375 2045 4380 2086
rect 4455 2045 4597 2109
rect 4661 2086 4677 2109
rect 4672 2045 4677 2086
rect 4741 2045 4757 2109
rect 4821 2045 4837 2109
rect 4901 2045 4917 2109
rect 4981 2045 4997 2109
rect 5061 2045 5203 2109
rect 5267 2045 5283 2109
rect 5347 2045 5363 2109
rect 5427 2045 5443 2109
rect 5507 2045 5523 2109
rect 5587 2086 5603 2109
rect 5587 2045 5592 2086
rect 5667 2045 5809 2109
rect 5873 2086 5889 2109
rect 5884 2045 5889 2086
rect 5953 2045 5969 2109
rect 6033 2045 6049 2109
rect 6113 2045 6129 2109
rect 6193 2045 6209 2109
rect 6273 2045 6377 2109
rect 6787 2125 7194 2140
rect 1463 2043 1956 2045
rect 1288 2022 1297 2043
rect 1214 2017 1297 2022
rect 1946 2022 1956 2043
rect 2020 2043 2184 2045
rect 2020 2022 2029 2043
rect 1946 2017 2029 2022
rect 2175 2022 2184 2043
rect 2248 2043 3168 2045
rect 2248 2022 2258 2043
rect 2175 2017 2258 2022
rect 3158 2022 3168 2043
rect 3232 2043 3396 2045
rect 3232 2022 3241 2043
rect 3158 2017 3241 2022
rect 3387 2022 3396 2043
rect 3460 2043 4380 2045
rect 3460 2022 3470 2043
rect 3387 2017 3470 2022
rect 4370 2022 4380 2043
rect 4444 2043 4608 2045
rect 4444 2022 4453 2043
rect 4370 2017 4453 2022
rect 4599 2022 4608 2043
rect 4672 2043 5592 2045
rect 4672 2022 4682 2043
rect 4599 2017 4682 2022
rect 5582 2022 5592 2043
rect 5656 2043 5820 2045
rect 5656 2022 5665 2043
rect 5582 2017 5665 2022
rect 5811 2022 5820 2043
rect 5884 2043 6377 2045
rect 6527 2088 6653 2098
rect 5884 2022 5894 2043
rect 5811 2017 5894 2022
rect 6527 2024 6558 2088
rect 6622 2024 6653 2088
rect 6787 2061 6828 2125
rect 6892 2061 6948 2125
rect 7012 2061 7091 2125
rect 7155 2061 7194 2125
rect 6787 2044 7194 2061
rect 7420 2111 7486 2265
rect 7546 2111 7606 3143
rect 7666 2173 7726 3203
rect 7786 2111 7846 3143
rect 7906 2173 7966 3203
rect 8026 3049 8092 3139
rect 8026 2985 8027 3049
rect 8091 2985 8092 3049
rect 8026 2969 8092 2985
rect 8026 2905 8027 2969
rect 8091 2905 8092 2969
rect 8026 2889 8092 2905
rect 8026 2825 8027 2889
rect 8091 2825 8092 2889
rect 8026 2809 8092 2825
rect 8026 2745 8027 2809
rect 8091 2745 8092 2809
rect 8026 2729 8092 2745
rect 8026 2665 8027 2729
rect 8091 2665 8092 2729
rect 8026 2649 8092 2665
rect 8026 2585 8027 2649
rect 8091 2585 8092 2649
rect 8026 2569 8092 2585
rect 8026 2505 8027 2569
rect 8091 2505 8092 2569
rect 8026 2489 8092 2505
rect 8026 2425 8027 2489
rect 8091 2425 8092 2489
rect 8026 2409 8092 2425
rect 8026 2345 8027 2409
rect 8091 2345 8092 2409
rect 8026 2329 8092 2345
rect 8026 2265 8027 2329
rect 8091 2265 8092 2329
rect 8026 2111 8092 2265
rect 7420 2109 8092 2111
rect 7420 2045 7524 2109
rect 7588 2045 7604 2109
rect 7668 2045 7684 2109
rect 7748 2045 7764 2109
rect 7828 2045 7844 2109
rect 7908 2086 7924 2109
rect 7908 2045 7913 2086
rect 7988 2045 8092 2109
rect 7420 2043 7913 2045
rect 6527 2014 6653 2024
rect 7903 2022 7913 2043
rect 7977 2043 8092 2045
rect 8152 3049 8218 3139
rect 8152 2985 8153 3049
rect 8217 2985 8218 3049
rect 8152 2969 8218 2985
rect 8152 2905 8153 2969
rect 8217 2905 8218 2969
rect 8152 2889 8218 2905
rect 8152 2825 8153 2889
rect 8217 2825 8218 2889
rect 8152 2809 8218 2825
rect 8152 2745 8153 2809
rect 8217 2745 8218 2809
rect 8152 2729 8218 2745
rect 8152 2665 8153 2729
rect 8217 2665 8218 2729
rect 8152 2649 8218 2665
rect 8152 2585 8153 2649
rect 8217 2585 8218 2649
rect 8152 2569 8218 2585
rect 8152 2505 8153 2569
rect 8217 2505 8218 2569
rect 8152 2489 8218 2505
rect 8152 2425 8153 2489
rect 8217 2425 8218 2489
rect 8152 2409 8218 2425
rect 8152 2345 8153 2409
rect 8217 2345 8218 2409
rect 8152 2329 8218 2345
rect 8152 2265 8153 2329
rect 8217 2265 8218 2329
rect 8152 2111 8218 2265
rect 8278 2111 8338 3143
rect 8398 2173 8458 3203
rect 8518 2111 8578 3143
rect 8638 2173 8698 3203
rect 8758 3049 8824 3139
rect 8758 2985 8759 3049
rect 8823 2985 8824 3049
rect 8758 2969 8824 2985
rect 8758 2905 8759 2969
rect 8823 2905 8824 2969
rect 8758 2889 8824 2905
rect 8758 2825 8759 2889
rect 8823 2825 8824 2889
rect 8758 2809 8824 2825
rect 8758 2745 8759 2809
rect 8823 2745 8824 2809
rect 8758 2729 8824 2745
rect 8758 2665 8759 2729
rect 8823 2665 8824 2729
rect 8758 2649 8824 2665
rect 8758 2585 8759 2649
rect 8823 2585 8824 2649
rect 8758 2569 8824 2585
rect 8758 2505 8759 2569
rect 8823 2505 8824 2569
rect 8758 2489 8824 2505
rect 8758 2425 8759 2489
rect 8823 2425 8824 2489
rect 8758 2409 8824 2425
rect 8758 2345 8759 2409
rect 8823 2345 8824 2409
rect 8758 2329 8824 2345
rect 8758 2265 8759 2329
rect 8823 2265 8824 2329
rect 8758 2111 8824 2265
rect 8884 2173 8944 3203
rect 9004 2111 9064 3143
rect 9124 2173 9184 3203
rect 9244 2111 9304 3143
rect 9364 3049 9430 3139
rect 9364 2985 9365 3049
rect 9429 2985 9430 3049
rect 9364 2969 9430 2985
rect 9364 2905 9365 2969
rect 9429 2905 9430 2969
rect 9364 2889 9430 2905
rect 9364 2825 9365 2889
rect 9429 2825 9430 2889
rect 9364 2809 9430 2825
rect 9364 2745 9365 2809
rect 9429 2745 9430 2809
rect 9364 2729 9430 2745
rect 9364 2665 9365 2729
rect 9429 2665 9430 2729
rect 9364 2649 9430 2665
rect 9364 2585 9365 2649
rect 9429 2585 9430 2649
rect 9364 2569 9430 2585
rect 9364 2505 9365 2569
rect 9429 2505 9430 2569
rect 9364 2489 9430 2505
rect 9364 2425 9365 2489
rect 9429 2425 9430 2489
rect 9364 2409 9430 2425
rect 9364 2345 9365 2409
rect 9429 2345 9430 2409
rect 9364 2329 9430 2345
rect 9364 2265 9365 2329
rect 9429 2265 9430 2329
rect 9364 2111 9430 2265
rect 9490 2111 9550 3143
rect 9610 2173 9670 3203
rect 9730 2111 9790 3143
rect 9850 2173 9910 3203
rect 9970 3049 10036 3139
rect 9970 2985 9971 3049
rect 10035 2985 10036 3049
rect 9970 2969 10036 2985
rect 9970 2905 9971 2969
rect 10035 2905 10036 2969
rect 9970 2889 10036 2905
rect 9970 2825 9971 2889
rect 10035 2825 10036 2889
rect 9970 2809 10036 2825
rect 9970 2745 9971 2809
rect 10035 2745 10036 2809
rect 9970 2729 10036 2745
rect 9970 2665 9971 2729
rect 10035 2665 10036 2729
rect 9970 2649 10036 2665
rect 9970 2585 9971 2649
rect 10035 2585 10036 2649
rect 9970 2569 10036 2585
rect 9970 2505 9971 2569
rect 10035 2505 10036 2569
rect 9970 2489 10036 2505
rect 9970 2425 9971 2489
rect 10035 2425 10036 2489
rect 9970 2409 10036 2425
rect 9970 2345 9971 2409
rect 10035 2345 10036 2409
rect 9970 2329 10036 2345
rect 9970 2265 9971 2329
rect 10035 2265 10036 2329
rect 9970 2111 10036 2265
rect 10096 2173 10156 3203
rect 10216 2111 10276 3143
rect 10336 2173 10396 3203
rect 10456 2111 10516 3143
rect 10576 3049 10642 3139
rect 10576 2985 10577 3049
rect 10641 2985 10642 3049
rect 10576 2969 10642 2985
rect 10576 2905 10577 2969
rect 10641 2905 10642 2969
rect 10576 2889 10642 2905
rect 10576 2825 10577 2889
rect 10641 2825 10642 2889
rect 10576 2809 10642 2825
rect 10576 2745 10577 2809
rect 10641 2745 10642 2809
rect 10576 2729 10642 2745
rect 10576 2665 10577 2729
rect 10641 2665 10642 2729
rect 10576 2649 10642 2665
rect 10576 2585 10577 2649
rect 10641 2585 10642 2649
rect 10576 2569 10642 2585
rect 10576 2505 10577 2569
rect 10641 2505 10642 2569
rect 10576 2489 10642 2505
rect 10576 2425 10577 2489
rect 10641 2425 10642 2489
rect 10576 2409 10642 2425
rect 10576 2345 10577 2409
rect 10641 2345 10642 2409
rect 10576 2329 10642 2345
rect 10576 2265 10577 2329
rect 10641 2265 10642 2329
rect 10576 2111 10642 2265
rect 10702 2111 10762 3143
rect 10822 2173 10882 3203
rect 10942 2111 11002 3143
rect 11062 2173 11122 3203
rect 11182 3049 11248 3139
rect 11182 2985 11183 3049
rect 11247 2985 11248 3049
rect 11182 2969 11248 2985
rect 11182 2905 11183 2969
rect 11247 2905 11248 2969
rect 11182 2889 11248 2905
rect 11182 2825 11183 2889
rect 11247 2825 11248 2889
rect 11182 2809 11248 2825
rect 11182 2745 11183 2809
rect 11247 2745 11248 2809
rect 11182 2729 11248 2745
rect 11182 2665 11183 2729
rect 11247 2665 11248 2729
rect 11182 2649 11248 2665
rect 11182 2585 11183 2649
rect 11247 2585 11248 2649
rect 11182 2569 11248 2585
rect 11182 2505 11183 2569
rect 11247 2505 11248 2569
rect 11182 2489 11248 2505
rect 11182 2425 11183 2489
rect 11247 2425 11248 2489
rect 11182 2409 11248 2425
rect 11182 2345 11183 2409
rect 11247 2345 11248 2409
rect 11182 2329 11248 2345
rect 11182 2265 11183 2329
rect 11247 2265 11248 2329
rect 11182 2111 11248 2265
rect 11308 2173 11368 3203
rect 11428 2111 11488 3143
rect 11548 2173 11608 3203
rect 11668 2111 11728 3143
rect 11788 3049 11854 3139
rect 11788 2985 11789 3049
rect 11853 2985 11854 3049
rect 11788 2969 11854 2985
rect 11788 2905 11789 2969
rect 11853 2905 11854 2969
rect 11788 2889 11854 2905
rect 11788 2825 11789 2889
rect 11853 2825 11854 2889
rect 11788 2809 11854 2825
rect 11788 2745 11789 2809
rect 11853 2745 11854 2809
rect 11788 2729 11854 2745
rect 11788 2665 11789 2729
rect 11853 2665 11854 2729
rect 11788 2649 11854 2665
rect 11788 2585 11789 2649
rect 11853 2585 11854 2649
rect 11788 2569 11854 2585
rect 11788 2505 11789 2569
rect 11853 2505 11854 2569
rect 11788 2489 11854 2505
rect 11788 2425 11789 2489
rect 11853 2425 11854 2489
rect 11788 2409 11854 2425
rect 11788 2345 11789 2409
rect 11853 2345 11854 2409
rect 11788 2329 11854 2345
rect 11788 2265 11789 2329
rect 11853 2265 11854 2329
rect 11788 2111 11854 2265
rect 11914 2111 11974 3143
rect 12034 2173 12094 3203
rect 12154 2111 12214 3143
rect 12274 2173 12334 3203
rect 12394 3049 12460 3139
rect 12394 2985 12395 3049
rect 12459 2985 12460 3049
rect 12394 2969 12460 2985
rect 12394 2905 12395 2969
rect 12459 2905 12460 2969
rect 12394 2889 12460 2905
rect 12394 2825 12395 2889
rect 12459 2825 12460 2889
rect 12394 2809 12460 2825
rect 12394 2745 12395 2809
rect 12459 2745 12460 2809
rect 12394 2729 12460 2745
rect 12394 2665 12395 2729
rect 12459 2665 12460 2729
rect 12394 2649 12460 2665
rect 12394 2585 12395 2649
rect 12459 2585 12460 2649
rect 12394 2569 12460 2585
rect 12394 2505 12395 2569
rect 12459 2505 12460 2569
rect 12394 2489 12460 2505
rect 12394 2425 12395 2489
rect 12459 2425 12460 2489
rect 12394 2409 12460 2425
rect 12394 2345 12395 2409
rect 12459 2345 12460 2409
rect 12394 2329 12460 2345
rect 12394 2265 12395 2329
rect 12459 2265 12460 2329
rect 12394 2111 12460 2265
rect 12520 2173 12580 3203
rect 12640 2111 12700 3143
rect 12760 2173 12820 3203
rect 12880 2111 12940 3143
rect 13000 3049 13066 3139
rect 13000 2985 13001 3049
rect 13065 2985 13066 3049
rect 13000 2969 13066 2985
rect 13000 2905 13001 2969
rect 13065 2905 13066 2969
rect 13000 2889 13066 2905
rect 13000 2825 13001 2889
rect 13065 2825 13066 2889
rect 13000 2809 13066 2825
rect 13000 2745 13001 2809
rect 13065 2745 13066 2809
rect 13000 2729 13066 2745
rect 13000 2665 13001 2729
rect 13065 2665 13066 2729
rect 13000 2649 13066 2665
rect 13000 2585 13001 2649
rect 13065 2585 13066 2649
rect 13000 2569 13066 2585
rect 13000 2505 13001 2569
rect 13065 2505 13066 2569
rect 13000 2489 13066 2505
rect 13000 2425 13001 2489
rect 13065 2425 13066 2489
rect 13000 2409 13066 2425
rect 13000 2345 13001 2409
rect 13065 2345 13066 2409
rect 13000 2329 13066 2345
rect 13000 2265 13001 2329
rect 13065 2265 13066 2329
rect 13128 2349 13254 2359
rect 13128 2285 13159 2349
rect 13223 2285 13254 2349
rect 13128 2275 13254 2285
rect 13000 2111 13066 2265
rect 8152 2109 13066 2111
rect 8152 2045 8256 2109
rect 8320 2045 8336 2109
rect 8400 2045 8416 2109
rect 8480 2045 8496 2109
rect 8560 2045 8576 2109
rect 8640 2086 8656 2109
rect 8640 2045 8645 2086
rect 8720 2045 8862 2109
rect 8926 2086 8942 2109
rect 8937 2045 8942 2086
rect 9006 2045 9022 2109
rect 9086 2045 9102 2109
rect 9166 2045 9182 2109
rect 9246 2045 9262 2109
rect 9326 2045 9468 2109
rect 9532 2045 9548 2109
rect 9612 2045 9628 2109
rect 9692 2045 9708 2109
rect 9772 2045 9788 2109
rect 9852 2086 9868 2109
rect 9852 2045 9857 2086
rect 9932 2045 10074 2109
rect 10138 2086 10154 2109
rect 10149 2045 10154 2086
rect 10218 2045 10234 2109
rect 10298 2045 10314 2109
rect 10378 2045 10394 2109
rect 10458 2045 10474 2109
rect 10538 2045 10680 2109
rect 10744 2045 10760 2109
rect 10824 2045 10840 2109
rect 10904 2045 10920 2109
rect 10984 2045 11000 2109
rect 11064 2086 11080 2109
rect 11064 2045 11069 2086
rect 11144 2045 11286 2109
rect 11350 2086 11366 2109
rect 11361 2045 11366 2086
rect 11430 2045 11446 2109
rect 11510 2045 11526 2109
rect 11590 2045 11606 2109
rect 11670 2045 11686 2109
rect 11750 2045 11892 2109
rect 11956 2045 11972 2109
rect 12036 2045 12052 2109
rect 12116 2045 12132 2109
rect 12196 2045 12212 2109
rect 12276 2086 12292 2109
rect 12276 2045 12281 2086
rect 12356 2045 12498 2109
rect 12562 2086 12578 2109
rect 12573 2045 12578 2086
rect 12642 2045 12658 2109
rect 12722 2045 12738 2109
rect 12802 2045 12818 2109
rect 12882 2045 12898 2109
rect 12962 2045 13066 2109
rect 8152 2043 8645 2045
rect 7977 2022 7986 2043
rect 7903 2017 7986 2022
rect 8635 2022 8645 2043
rect 8709 2043 8873 2045
rect 8709 2022 8718 2043
rect 8635 2017 8718 2022
rect 8864 2022 8873 2043
rect 8937 2043 9857 2045
rect 8937 2022 8947 2043
rect 8864 2017 8947 2022
rect 9847 2022 9857 2043
rect 9921 2043 10085 2045
rect 9921 2022 9930 2043
rect 9847 2017 9930 2022
rect 10076 2022 10085 2043
rect 10149 2043 11069 2045
rect 10149 2022 10159 2043
rect 10076 2017 10159 2022
rect 11059 2022 11069 2043
rect 11133 2043 11297 2045
rect 11133 2022 11142 2043
rect 11059 2017 11142 2022
rect 11288 2022 11297 2043
rect 11361 2043 12281 2045
rect 11361 2022 11371 2043
rect 11288 2017 11371 2022
rect 12271 2022 12281 2043
rect 12345 2043 12509 2045
rect 12345 2022 12354 2043
rect 12271 2017 12354 2022
rect 12500 2022 12509 2043
rect 12573 2043 13066 2045
rect 13216 2088 13342 2098
rect 12573 2022 12583 2043
rect 12500 2017 12583 2022
rect 13216 2024 13247 2088
rect 13311 2024 13342 2088
rect 13216 2014 13342 2024
rect 1573 1884 1655 1890
rect 1573 1862 1582 1884
rect 1085 1860 1582 1862
rect 1646 1862 1655 1884
rect 2305 1884 2387 1890
rect 2305 1862 2314 1884
rect 1646 1860 1757 1862
rect 1085 1796 1189 1860
rect 1253 1796 1269 1860
rect 1333 1796 1349 1860
rect 1413 1796 1429 1860
rect 1493 1796 1509 1860
rect 1573 1820 1582 1860
rect 1573 1796 1589 1820
rect 1653 1796 1757 1860
rect 1085 1794 1757 1796
rect 1085 1640 1151 1794
rect 1085 1576 1086 1640
rect 1150 1576 1151 1640
rect 1085 1560 1151 1576
rect 1085 1496 1086 1560
rect 1150 1496 1151 1560
rect 1085 1480 1151 1496
rect 1085 1416 1086 1480
rect 1150 1416 1151 1480
rect 1085 1400 1151 1416
rect 1085 1336 1086 1400
rect 1150 1336 1151 1400
rect 1085 1320 1151 1336
rect 1085 1256 1086 1320
rect 1150 1256 1151 1320
rect 1085 1240 1151 1256
rect 1085 1176 1086 1240
rect 1150 1176 1151 1240
rect 1085 1160 1151 1176
rect 1085 1096 1086 1160
rect 1150 1096 1151 1160
rect 1085 1080 1151 1096
rect 1085 1016 1086 1080
rect 1150 1016 1151 1080
rect 1085 1000 1151 1016
rect 1085 936 1086 1000
rect 1150 936 1151 1000
rect 1085 920 1151 936
rect 1085 856 1086 920
rect 1150 856 1151 920
rect 1085 766 1151 856
rect 1211 762 1271 1794
rect 694 698 819 708
rect 1331 702 1391 1732
rect 1451 762 1511 1794
rect 1571 702 1631 1732
rect 1691 1640 1757 1794
rect 1691 1576 1692 1640
rect 1756 1576 1757 1640
rect 1691 1560 1757 1576
rect 1691 1496 1692 1560
rect 1756 1496 1757 1560
rect 1691 1480 1757 1496
rect 1691 1416 1692 1480
rect 1756 1416 1757 1480
rect 1691 1400 1757 1416
rect 1691 1336 1692 1400
rect 1756 1336 1757 1400
rect 1691 1320 1757 1336
rect 1691 1256 1692 1320
rect 1756 1256 1757 1320
rect 1691 1240 1757 1256
rect 1691 1176 1692 1240
rect 1756 1176 1757 1240
rect 1691 1160 1757 1176
rect 1691 1096 1692 1160
rect 1756 1096 1757 1160
rect 1691 1080 1757 1096
rect 1691 1016 1692 1080
rect 1756 1016 1757 1080
rect 1691 1000 1757 1016
rect 1691 936 1692 1000
rect 1756 936 1757 1000
rect 1691 920 1757 936
rect 1691 856 1692 920
rect 1756 856 1757 920
rect 1691 766 1757 856
rect 1817 1860 2314 1862
rect 2378 1862 2387 1884
rect 2525 1884 2607 1890
rect 2525 1862 2534 1884
rect 2378 1860 2534 1862
rect 2598 1862 2607 1884
rect 3517 1884 3599 1890
rect 3517 1862 3526 1884
rect 2598 1860 3526 1862
rect 3590 1862 3599 1884
rect 3737 1884 3819 1890
rect 3737 1862 3746 1884
rect 3590 1860 3746 1862
rect 3810 1862 3819 1884
rect 4855 1884 4937 1890
rect 4855 1862 4864 1884
rect 3810 1860 4307 1862
rect 1817 1796 1921 1860
rect 1985 1796 2001 1860
rect 2065 1796 2081 1860
rect 2145 1796 2161 1860
rect 2225 1796 2241 1860
rect 2305 1820 2314 1860
rect 2305 1796 2321 1820
rect 2385 1796 2527 1860
rect 2598 1820 2607 1860
rect 2591 1796 2607 1820
rect 2671 1796 2687 1860
rect 2751 1796 2767 1860
rect 2831 1796 2847 1860
rect 2911 1796 2927 1860
rect 2991 1796 3133 1860
rect 3197 1796 3213 1860
rect 3277 1796 3293 1860
rect 3357 1796 3373 1860
rect 3437 1796 3453 1860
rect 3517 1820 3526 1860
rect 3517 1796 3533 1820
rect 3597 1796 3739 1860
rect 3810 1820 3819 1860
rect 3803 1796 3819 1820
rect 3883 1796 3899 1860
rect 3963 1796 3979 1860
rect 4043 1796 4059 1860
rect 4123 1796 4139 1860
rect 4203 1796 4307 1860
rect 1817 1794 4307 1796
rect 1817 1640 1883 1794
rect 1817 1576 1818 1640
rect 1882 1576 1883 1640
rect 1817 1560 1883 1576
rect 1817 1496 1818 1560
rect 1882 1496 1883 1560
rect 1817 1480 1883 1496
rect 1817 1416 1818 1480
rect 1882 1416 1883 1480
rect 1817 1400 1883 1416
rect 1817 1336 1818 1400
rect 1882 1336 1883 1400
rect 1817 1320 1883 1336
rect 1817 1256 1818 1320
rect 1882 1256 1883 1320
rect 1817 1240 1883 1256
rect 1817 1176 1818 1240
rect 1882 1176 1883 1240
rect 1817 1160 1883 1176
rect 1817 1096 1818 1160
rect 1882 1096 1883 1160
rect 1817 1080 1883 1096
rect 1817 1016 1818 1080
rect 1882 1016 1883 1080
rect 1817 1000 1883 1016
rect 1817 936 1818 1000
rect 1882 936 1883 1000
rect 1817 920 1883 936
rect 1817 856 1818 920
rect 1882 856 1883 920
rect 1817 766 1883 856
rect 1943 762 2003 1794
rect 2063 702 2123 1732
rect 2183 762 2243 1794
rect 2303 702 2363 1732
rect 2423 1640 2489 1794
rect 2423 1576 2424 1640
rect 2488 1576 2489 1640
rect 2423 1560 2489 1576
rect 2423 1496 2424 1560
rect 2488 1496 2489 1560
rect 2423 1480 2489 1496
rect 2423 1416 2424 1480
rect 2488 1416 2489 1480
rect 2423 1400 2489 1416
rect 2423 1336 2424 1400
rect 2488 1336 2489 1400
rect 2423 1320 2489 1336
rect 2423 1256 2424 1320
rect 2488 1256 2489 1320
rect 2423 1240 2489 1256
rect 2423 1176 2424 1240
rect 2488 1176 2489 1240
rect 2423 1160 2489 1176
rect 2423 1096 2424 1160
rect 2488 1096 2489 1160
rect 2423 1080 2489 1096
rect 2423 1016 2424 1080
rect 2488 1016 2489 1080
rect 2423 1000 2489 1016
rect 2423 936 2424 1000
rect 2488 936 2489 1000
rect 2423 920 2489 936
rect 2423 856 2424 920
rect 2488 856 2489 920
rect 2423 766 2489 856
rect 2549 702 2609 1732
rect 2669 762 2729 1794
rect 2789 702 2849 1732
rect 2909 762 2969 1794
rect 3029 1640 3095 1794
rect 3029 1576 3030 1640
rect 3094 1576 3095 1640
rect 3029 1560 3095 1576
rect 3029 1496 3030 1560
rect 3094 1496 3095 1560
rect 3029 1480 3095 1496
rect 3029 1416 3030 1480
rect 3094 1416 3095 1480
rect 3029 1400 3095 1416
rect 3029 1336 3030 1400
rect 3094 1336 3095 1400
rect 3029 1320 3095 1336
rect 3029 1256 3030 1320
rect 3094 1256 3095 1320
rect 3029 1240 3095 1256
rect 3029 1176 3030 1240
rect 3094 1176 3095 1240
rect 3029 1160 3095 1176
rect 3029 1096 3030 1160
rect 3094 1096 3095 1160
rect 3029 1080 3095 1096
rect 3029 1016 3030 1080
rect 3094 1016 3095 1080
rect 3029 1000 3095 1016
rect 3029 936 3030 1000
rect 3094 936 3095 1000
rect 3029 920 3095 936
rect 3029 856 3030 920
rect 3094 856 3095 920
rect 3029 766 3095 856
rect 3155 762 3215 1794
rect 3275 702 3335 1732
rect 3395 762 3455 1794
rect 3515 702 3575 1732
rect 3635 1640 3701 1794
rect 3635 1576 3636 1640
rect 3700 1576 3701 1640
rect 3635 1560 3701 1576
rect 3635 1496 3636 1560
rect 3700 1496 3701 1560
rect 3635 1480 3701 1496
rect 3635 1416 3636 1480
rect 3700 1416 3701 1480
rect 3635 1400 3701 1416
rect 3635 1336 3636 1400
rect 3700 1336 3701 1400
rect 3635 1320 3701 1336
rect 3635 1256 3636 1320
rect 3700 1256 3701 1320
rect 3635 1240 3701 1256
rect 3635 1176 3636 1240
rect 3700 1176 3701 1240
rect 3635 1160 3701 1176
rect 3635 1096 3636 1160
rect 3700 1096 3701 1160
rect 3635 1080 3701 1096
rect 3635 1016 3636 1080
rect 3700 1016 3701 1080
rect 3635 1000 3701 1016
rect 3635 936 3636 1000
rect 3700 936 3701 1000
rect 3635 920 3701 936
rect 3635 856 3636 920
rect 3700 856 3701 920
rect 3635 766 3701 856
rect 3761 702 3821 1732
rect 3881 762 3941 1794
rect 4001 702 4061 1732
rect 4121 762 4181 1794
rect 4241 1640 4307 1794
rect 4241 1576 4242 1640
rect 4306 1576 4307 1640
rect 4241 1560 4307 1576
rect 4241 1496 4242 1560
rect 4306 1496 4307 1560
rect 4241 1480 4307 1496
rect 4241 1416 4242 1480
rect 4306 1416 4307 1480
rect 4241 1400 4307 1416
rect 4241 1336 4242 1400
rect 4306 1336 4307 1400
rect 4241 1320 4307 1336
rect 4241 1256 4242 1320
rect 4306 1256 4307 1320
rect 4241 1240 4307 1256
rect 4241 1176 4242 1240
rect 4306 1176 4307 1240
rect 4241 1160 4307 1176
rect 4241 1096 4242 1160
rect 4306 1096 4307 1160
rect 4241 1080 4307 1096
rect 4241 1016 4242 1080
rect 4306 1016 4307 1080
rect 4241 1000 4307 1016
rect 4241 936 4242 1000
rect 4306 936 4307 1000
rect 4241 920 4307 936
rect 4241 856 4242 920
rect 4306 856 4307 920
rect 4241 766 4307 856
rect 4367 1860 4864 1862
rect 4928 1862 4937 1884
rect 5075 1884 5157 1890
rect 5075 1862 5084 1884
rect 4928 1860 5084 1862
rect 5148 1862 5157 1884
rect 5807 1884 5889 1890
rect 5807 1862 5816 1884
rect 5148 1860 5645 1862
rect 4367 1796 4471 1860
rect 4535 1796 4551 1860
rect 4615 1796 4631 1860
rect 4695 1796 4711 1860
rect 4775 1796 4791 1860
rect 4855 1820 4864 1860
rect 4855 1796 4871 1820
rect 4935 1796 5077 1860
rect 5148 1820 5157 1860
rect 5141 1796 5157 1820
rect 5221 1796 5237 1860
rect 5301 1796 5317 1860
rect 5381 1796 5397 1860
rect 5461 1796 5477 1860
rect 5541 1796 5645 1860
rect 4367 1794 5645 1796
rect 4367 1640 4433 1794
rect 4367 1576 4368 1640
rect 4432 1576 4433 1640
rect 4367 1560 4433 1576
rect 4367 1496 4368 1560
rect 4432 1496 4433 1560
rect 4367 1480 4433 1496
rect 4367 1416 4368 1480
rect 4432 1416 4433 1480
rect 4367 1400 4433 1416
rect 4367 1336 4368 1400
rect 4432 1336 4433 1400
rect 4367 1320 4433 1336
rect 4367 1256 4368 1320
rect 4432 1256 4433 1320
rect 4367 1240 4433 1256
rect 4367 1176 4368 1240
rect 4432 1176 4433 1240
rect 4367 1160 4433 1176
rect 4367 1096 4368 1160
rect 4432 1096 4433 1160
rect 4367 1080 4433 1096
rect 4367 1016 4368 1080
rect 4432 1016 4433 1080
rect 4367 1000 4433 1016
rect 4367 936 4368 1000
rect 4432 936 4433 1000
rect 4367 920 4433 936
rect 4367 856 4368 920
rect 4432 856 4433 920
rect 4367 766 4433 856
rect 4493 762 4553 1794
rect 4613 702 4673 1732
rect 4733 762 4793 1794
rect 4853 702 4913 1732
rect 4973 1640 5039 1794
rect 4973 1576 4974 1640
rect 5038 1576 5039 1640
rect 4973 1560 5039 1576
rect 4973 1496 4974 1560
rect 5038 1496 5039 1560
rect 4973 1480 5039 1496
rect 4973 1416 4974 1480
rect 5038 1416 5039 1480
rect 4973 1400 5039 1416
rect 4973 1336 4974 1400
rect 5038 1336 5039 1400
rect 4973 1320 5039 1336
rect 4973 1256 4974 1320
rect 5038 1256 5039 1320
rect 4973 1240 5039 1256
rect 4973 1176 4974 1240
rect 5038 1176 5039 1240
rect 4973 1160 5039 1176
rect 4973 1096 4974 1160
rect 5038 1096 5039 1160
rect 4973 1080 5039 1096
rect 4973 1016 4974 1080
rect 5038 1016 5039 1080
rect 4973 1000 5039 1016
rect 4973 936 4974 1000
rect 5038 936 5039 1000
rect 4973 920 5039 936
rect 4973 856 4974 920
rect 5038 856 5039 920
rect 4973 766 5039 856
rect 5099 702 5159 1732
rect 5219 762 5279 1794
rect 5339 702 5399 1732
rect 5459 762 5519 1794
rect 5579 1640 5645 1794
rect 5579 1576 5580 1640
rect 5644 1576 5645 1640
rect 5579 1560 5645 1576
rect 5579 1496 5580 1560
rect 5644 1496 5645 1560
rect 5579 1480 5645 1496
rect 5579 1416 5580 1480
rect 5644 1416 5645 1480
rect 5579 1400 5645 1416
rect 5579 1336 5580 1400
rect 5644 1336 5645 1400
rect 5579 1320 5645 1336
rect 5579 1256 5580 1320
rect 5644 1256 5645 1320
rect 5579 1240 5645 1256
rect 5579 1176 5580 1240
rect 5644 1176 5645 1240
rect 5579 1160 5645 1176
rect 5579 1096 5580 1160
rect 5644 1096 5645 1160
rect 5579 1080 5645 1096
rect 5579 1016 5580 1080
rect 5644 1016 5645 1080
rect 5579 1000 5645 1016
rect 5579 936 5580 1000
rect 5644 936 5645 1000
rect 5579 920 5645 936
rect 5579 856 5580 920
rect 5644 856 5645 920
rect 5579 766 5645 856
rect 5705 1860 5816 1862
rect 5880 1862 5889 1884
rect 6527 1885 6653 1895
rect 5880 1860 6377 1862
rect 5705 1796 5809 1860
rect 5880 1820 5889 1860
rect 5873 1796 5889 1820
rect 5953 1796 5969 1860
rect 6033 1796 6049 1860
rect 6113 1796 6129 1860
rect 6193 1796 6209 1860
rect 6273 1796 6377 1860
rect 6527 1821 6558 1885
rect 6622 1821 6653 1885
rect 8262 1884 8344 1890
rect 8262 1862 8271 1884
rect 6527 1811 6653 1821
rect 7774 1860 8271 1862
rect 8335 1862 8344 1884
rect 8994 1884 9076 1890
rect 8994 1862 9003 1884
rect 8335 1860 8446 1862
rect 6553 1810 6627 1811
rect 5705 1794 6377 1796
rect 5705 1640 5771 1794
rect 5705 1576 5706 1640
rect 5770 1576 5771 1640
rect 5705 1560 5771 1576
rect 5705 1496 5706 1560
rect 5770 1496 5771 1560
rect 5705 1480 5771 1496
rect 5705 1416 5706 1480
rect 5770 1416 5771 1480
rect 5705 1400 5771 1416
rect 5705 1336 5706 1400
rect 5770 1336 5771 1400
rect 5705 1320 5771 1336
rect 5705 1256 5706 1320
rect 5770 1256 5771 1320
rect 5705 1240 5771 1256
rect 5705 1176 5706 1240
rect 5770 1176 5771 1240
rect 5705 1160 5771 1176
rect 5705 1096 5706 1160
rect 5770 1096 5771 1160
rect 5705 1080 5771 1096
rect 5705 1016 5706 1080
rect 5770 1016 5771 1080
rect 5705 1000 5771 1016
rect 5705 936 5706 1000
rect 5770 936 5771 1000
rect 5705 920 5771 936
rect 5705 856 5706 920
rect 5770 856 5771 920
rect 5705 766 5771 856
rect 5831 702 5891 1732
rect 5951 762 6011 1794
rect 6071 702 6131 1732
rect 6191 762 6251 1794
rect 6311 1640 6377 1794
rect 6311 1576 6312 1640
rect 6376 1576 6377 1640
rect 7774 1796 7878 1860
rect 7942 1796 7958 1860
rect 8022 1796 8038 1860
rect 8102 1796 8118 1860
rect 8182 1796 8198 1860
rect 8262 1820 8271 1860
rect 8262 1796 8278 1820
rect 8342 1796 8446 1860
rect 7774 1794 8446 1796
rect 7774 1640 7840 1794
rect 6311 1560 6377 1576
rect 6311 1496 6312 1560
rect 6376 1496 6377 1560
rect 6437 1623 6562 1633
rect 6437 1559 6467 1623
rect 6531 1559 6562 1623
rect 6437 1549 6562 1559
rect 7774 1576 7775 1640
rect 7839 1576 7840 1640
rect 7774 1560 7840 1576
rect 6311 1480 6377 1496
rect 6311 1416 6312 1480
rect 6376 1416 6377 1480
rect 6311 1400 6377 1416
rect 6311 1336 6312 1400
rect 6376 1336 6377 1400
rect 6311 1320 6377 1336
rect 6311 1256 6312 1320
rect 6376 1256 6377 1320
rect 6311 1240 6377 1256
rect 6311 1176 6312 1240
rect 6376 1176 6377 1240
rect 6311 1160 6377 1176
rect 6311 1096 6312 1160
rect 6376 1096 6377 1160
rect 6311 1080 6377 1096
rect 6311 1016 6312 1080
rect 6376 1016 6377 1080
rect 6311 1000 6377 1016
rect 6311 936 6312 1000
rect 6376 936 6377 1000
rect 6311 920 6377 936
rect 6311 856 6312 920
rect 6376 856 6377 920
rect 6311 766 6377 856
rect 7774 1496 7775 1560
rect 7839 1496 7840 1560
rect 7774 1480 7840 1496
rect 7774 1416 7775 1480
rect 7839 1416 7840 1480
rect 7774 1400 7840 1416
rect 7774 1336 7775 1400
rect 7839 1336 7840 1400
rect 7774 1320 7840 1336
rect 7774 1256 7775 1320
rect 7839 1256 7840 1320
rect 7774 1240 7840 1256
rect 7774 1176 7775 1240
rect 7839 1176 7840 1240
rect 7774 1160 7840 1176
rect 7774 1096 7775 1160
rect 7839 1096 7840 1160
rect 7774 1080 7840 1096
rect 7774 1016 7775 1080
rect 7839 1016 7840 1080
rect 7774 1000 7840 1016
rect 7774 936 7775 1000
rect 7839 936 7840 1000
rect 7774 920 7840 936
rect 7774 856 7775 920
rect 7839 856 7840 920
rect 7774 766 7840 856
rect 7900 762 7960 1794
rect 694 634 724 698
rect 788 634 819 698
rect 1085 700 1757 702
rect 1085 636 1189 700
rect 1253 636 1269 700
rect 1333 636 1349 700
rect 1413 636 1429 700
rect 1493 636 1509 700
rect 1573 636 1589 700
rect 1653 636 1757 700
rect 1085 634 1757 636
rect 1817 700 4307 702
rect 1817 636 1921 700
rect 1985 636 2001 700
rect 2065 636 2081 700
rect 2145 636 2161 700
rect 2225 636 2241 700
rect 2305 636 2321 700
rect 2385 636 2527 700
rect 2591 636 2607 700
rect 2671 636 2687 700
rect 2751 636 2767 700
rect 2831 636 2847 700
rect 2911 636 2927 700
rect 2991 636 3133 700
rect 3197 636 3213 700
rect 3277 636 3293 700
rect 3357 636 3373 700
rect 3437 636 3453 700
rect 3517 636 3533 700
rect 3597 636 3739 700
rect 3803 636 3819 700
rect 3883 636 3899 700
rect 3963 636 3979 700
rect 4043 636 4059 700
rect 4123 636 4139 700
rect 4203 636 4307 700
rect 1817 634 4307 636
rect 4367 700 5645 702
rect 4367 636 4471 700
rect 4535 636 4551 700
rect 4615 636 4631 700
rect 4695 636 4711 700
rect 4775 636 4791 700
rect 4855 636 4871 700
rect 4935 636 5077 700
rect 5141 636 5157 700
rect 5221 636 5237 700
rect 5301 636 5317 700
rect 5381 636 5397 700
rect 5461 636 5477 700
rect 5541 636 5645 700
rect 4367 634 5645 636
rect 5705 700 6377 702
rect 5705 636 5809 700
rect 5873 636 5889 700
rect 5953 636 5969 700
rect 6033 636 6049 700
rect 6113 636 6129 700
rect 6193 636 6209 700
rect 6273 636 6377 700
rect 5705 634 6377 636
rect 7383 698 7508 708
rect 8020 702 8080 1732
rect 8140 762 8200 1794
rect 8260 702 8320 1732
rect 8380 1640 8446 1794
rect 8380 1576 8381 1640
rect 8445 1576 8446 1640
rect 8380 1560 8446 1576
rect 8380 1496 8381 1560
rect 8445 1496 8446 1560
rect 8380 1480 8446 1496
rect 8380 1416 8381 1480
rect 8445 1416 8446 1480
rect 8380 1400 8446 1416
rect 8380 1336 8381 1400
rect 8445 1336 8446 1400
rect 8380 1320 8446 1336
rect 8380 1256 8381 1320
rect 8445 1256 8446 1320
rect 8380 1240 8446 1256
rect 8380 1176 8381 1240
rect 8445 1176 8446 1240
rect 8380 1160 8446 1176
rect 8380 1096 8381 1160
rect 8445 1096 8446 1160
rect 8380 1080 8446 1096
rect 8380 1016 8381 1080
rect 8445 1016 8446 1080
rect 8380 1000 8446 1016
rect 8380 936 8381 1000
rect 8445 936 8446 1000
rect 8380 920 8446 936
rect 8380 856 8381 920
rect 8445 856 8446 920
rect 8380 766 8446 856
rect 8506 1860 9003 1862
rect 9067 1862 9076 1884
rect 9214 1884 9296 1890
rect 9214 1862 9223 1884
rect 9067 1860 9223 1862
rect 9287 1862 9296 1884
rect 10206 1884 10288 1890
rect 10206 1862 10215 1884
rect 9287 1860 10215 1862
rect 10279 1862 10288 1884
rect 10426 1884 10508 1890
rect 10426 1862 10435 1884
rect 10279 1860 10435 1862
rect 10499 1862 10508 1884
rect 11544 1884 11626 1890
rect 11544 1862 11553 1884
rect 10499 1860 10996 1862
rect 8506 1796 8610 1860
rect 8674 1796 8690 1860
rect 8754 1796 8770 1860
rect 8834 1796 8850 1860
rect 8914 1796 8930 1860
rect 8994 1820 9003 1860
rect 8994 1796 9010 1820
rect 9074 1796 9216 1860
rect 9287 1820 9296 1860
rect 9280 1796 9296 1820
rect 9360 1796 9376 1860
rect 9440 1796 9456 1860
rect 9520 1796 9536 1860
rect 9600 1796 9616 1860
rect 9680 1796 9822 1860
rect 9886 1796 9902 1860
rect 9966 1796 9982 1860
rect 10046 1796 10062 1860
rect 10126 1796 10142 1860
rect 10206 1820 10215 1860
rect 10206 1796 10222 1820
rect 10286 1796 10428 1860
rect 10499 1820 10508 1860
rect 10492 1796 10508 1820
rect 10572 1796 10588 1860
rect 10652 1796 10668 1860
rect 10732 1796 10748 1860
rect 10812 1796 10828 1860
rect 10892 1796 10996 1860
rect 8506 1794 10996 1796
rect 8506 1640 8572 1794
rect 8506 1576 8507 1640
rect 8571 1576 8572 1640
rect 8506 1560 8572 1576
rect 8506 1496 8507 1560
rect 8571 1496 8572 1560
rect 8506 1480 8572 1496
rect 8506 1416 8507 1480
rect 8571 1416 8572 1480
rect 8506 1400 8572 1416
rect 8506 1336 8507 1400
rect 8571 1336 8572 1400
rect 8506 1320 8572 1336
rect 8506 1256 8507 1320
rect 8571 1256 8572 1320
rect 8506 1240 8572 1256
rect 8506 1176 8507 1240
rect 8571 1176 8572 1240
rect 8506 1160 8572 1176
rect 8506 1096 8507 1160
rect 8571 1096 8572 1160
rect 8506 1080 8572 1096
rect 8506 1016 8507 1080
rect 8571 1016 8572 1080
rect 8506 1000 8572 1016
rect 8506 936 8507 1000
rect 8571 936 8572 1000
rect 8506 920 8572 936
rect 8506 856 8507 920
rect 8571 856 8572 920
rect 8506 766 8572 856
rect 8632 762 8692 1794
rect 8752 702 8812 1732
rect 8872 762 8932 1794
rect 8992 702 9052 1732
rect 9112 1640 9178 1794
rect 9112 1576 9113 1640
rect 9177 1576 9178 1640
rect 9112 1560 9178 1576
rect 9112 1496 9113 1560
rect 9177 1496 9178 1560
rect 9112 1480 9178 1496
rect 9112 1416 9113 1480
rect 9177 1416 9178 1480
rect 9112 1400 9178 1416
rect 9112 1336 9113 1400
rect 9177 1336 9178 1400
rect 9112 1320 9178 1336
rect 9112 1256 9113 1320
rect 9177 1256 9178 1320
rect 9112 1240 9178 1256
rect 9112 1176 9113 1240
rect 9177 1176 9178 1240
rect 9112 1160 9178 1176
rect 9112 1096 9113 1160
rect 9177 1096 9178 1160
rect 9112 1080 9178 1096
rect 9112 1016 9113 1080
rect 9177 1016 9178 1080
rect 9112 1000 9178 1016
rect 9112 936 9113 1000
rect 9177 936 9178 1000
rect 9112 920 9178 936
rect 9112 856 9113 920
rect 9177 856 9178 920
rect 9112 766 9178 856
rect 9238 702 9298 1732
rect 9358 762 9418 1794
rect 9478 702 9538 1732
rect 9598 762 9658 1794
rect 9718 1640 9784 1794
rect 9718 1576 9719 1640
rect 9783 1576 9784 1640
rect 9718 1560 9784 1576
rect 9718 1496 9719 1560
rect 9783 1496 9784 1560
rect 9718 1480 9784 1496
rect 9718 1416 9719 1480
rect 9783 1416 9784 1480
rect 9718 1400 9784 1416
rect 9718 1336 9719 1400
rect 9783 1336 9784 1400
rect 9718 1320 9784 1336
rect 9718 1256 9719 1320
rect 9783 1256 9784 1320
rect 9718 1240 9784 1256
rect 9718 1176 9719 1240
rect 9783 1176 9784 1240
rect 9718 1160 9784 1176
rect 9718 1096 9719 1160
rect 9783 1096 9784 1160
rect 9718 1080 9784 1096
rect 9718 1016 9719 1080
rect 9783 1016 9784 1080
rect 9718 1000 9784 1016
rect 9718 936 9719 1000
rect 9783 936 9784 1000
rect 9718 920 9784 936
rect 9718 856 9719 920
rect 9783 856 9784 920
rect 9718 766 9784 856
rect 9844 762 9904 1794
rect 9964 702 10024 1732
rect 10084 762 10144 1794
rect 10204 702 10264 1732
rect 10324 1640 10390 1794
rect 10324 1576 10325 1640
rect 10389 1576 10390 1640
rect 10324 1560 10390 1576
rect 10324 1496 10325 1560
rect 10389 1496 10390 1560
rect 10324 1480 10390 1496
rect 10324 1416 10325 1480
rect 10389 1416 10390 1480
rect 10324 1400 10390 1416
rect 10324 1336 10325 1400
rect 10389 1336 10390 1400
rect 10324 1320 10390 1336
rect 10324 1256 10325 1320
rect 10389 1256 10390 1320
rect 10324 1240 10390 1256
rect 10324 1176 10325 1240
rect 10389 1176 10390 1240
rect 10324 1160 10390 1176
rect 10324 1096 10325 1160
rect 10389 1096 10390 1160
rect 10324 1080 10390 1096
rect 10324 1016 10325 1080
rect 10389 1016 10390 1080
rect 10324 1000 10390 1016
rect 10324 936 10325 1000
rect 10389 936 10390 1000
rect 10324 920 10390 936
rect 10324 856 10325 920
rect 10389 856 10390 920
rect 10324 766 10390 856
rect 10450 702 10510 1732
rect 10570 762 10630 1794
rect 10690 702 10750 1732
rect 10810 762 10870 1794
rect 10930 1640 10996 1794
rect 10930 1576 10931 1640
rect 10995 1576 10996 1640
rect 10930 1560 10996 1576
rect 10930 1496 10931 1560
rect 10995 1496 10996 1560
rect 10930 1480 10996 1496
rect 10930 1416 10931 1480
rect 10995 1416 10996 1480
rect 10930 1400 10996 1416
rect 10930 1336 10931 1400
rect 10995 1336 10996 1400
rect 10930 1320 10996 1336
rect 10930 1256 10931 1320
rect 10995 1256 10996 1320
rect 10930 1240 10996 1256
rect 10930 1176 10931 1240
rect 10995 1176 10996 1240
rect 10930 1160 10996 1176
rect 10930 1096 10931 1160
rect 10995 1096 10996 1160
rect 10930 1080 10996 1096
rect 10930 1016 10931 1080
rect 10995 1016 10996 1080
rect 10930 1000 10996 1016
rect 10930 936 10931 1000
rect 10995 936 10996 1000
rect 10930 920 10996 936
rect 10930 856 10931 920
rect 10995 856 10996 920
rect 10930 766 10996 856
rect 11056 1860 11553 1862
rect 11617 1862 11626 1884
rect 11764 1884 11846 1890
rect 11764 1862 11773 1884
rect 11617 1860 11773 1862
rect 11837 1862 11846 1884
rect 12496 1884 12578 1890
rect 12496 1862 12505 1884
rect 11837 1860 12334 1862
rect 11056 1796 11160 1860
rect 11224 1796 11240 1860
rect 11304 1796 11320 1860
rect 11384 1796 11400 1860
rect 11464 1796 11480 1860
rect 11544 1820 11553 1860
rect 11544 1796 11560 1820
rect 11624 1796 11766 1860
rect 11837 1820 11846 1860
rect 11830 1796 11846 1820
rect 11910 1796 11926 1860
rect 11990 1796 12006 1860
rect 12070 1796 12086 1860
rect 12150 1796 12166 1860
rect 12230 1796 12334 1860
rect 11056 1794 12334 1796
rect 11056 1640 11122 1794
rect 11056 1576 11057 1640
rect 11121 1576 11122 1640
rect 11056 1560 11122 1576
rect 11056 1496 11057 1560
rect 11121 1496 11122 1560
rect 11056 1480 11122 1496
rect 11056 1416 11057 1480
rect 11121 1416 11122 1480
rect 11056 1400 11122 1416
rect 11056 1336 11057 1400
rect 11121 1336 11122 1400
rect 11056 1320 11122 1336
rect 11056 1256 11057 1320
rect 11121 1256 11122 1320
rect 11056 1240 11122 1256
rect 11056 1176 11057 1240
rect 11121 1176 11122 1240
rect 11056 1160 11122 1176
rect 11056 1096 11057 1160
rect 11121 1096 11122 1160
rect 11056 1080 11122 1096
rect 11056 1016 11057 1080
rect 11121 1016 11122 1080
rect 11056 1000 11122 1016
rect 11056 936 11057 1000
rect 11121 936 11122 1000
rect 11056 920 11122 936
rect 11056 856 11057 920
rect 11121 856 11122 920
rect 11056 766 11122 856
rect 11182 762 11242 1794
rect 11302 702 11362 1732
rect 11422 762 11482 1794
rect 11542 702 11602 1732
rect 11662 1640 11728 1794
rect 11662 1576 11663 1640
rect 11727 1576 11728 1640
rect 11662 1560 11728 1576
rect 11662 1496 11663 1560
rect 11727 1496 11728 1560
rect 11662 1480 11728 1496
rect 11662 1416 11663 1480
rect 11727 1416 11728 1480
rect 11662 1400 11728 1416
rect 11662 1336 11663 1400
rect 11727 1336 11728 1400
rect 11662 1320 11728 1336
rect 11662 1256 11663 1320
rect 11727 1256 11728 1320
rect 11662 1240 11728 1256
rect 11662 1176 11663 1240
rect 11727 1176 11728 1240
rect 11662 1160 11728 1176
rect 11662 1096 11663 1160
rect 11727 1096 11728 1160
rect 11662 1080 11728 1096
rect 11662 1016 11663 1080
rect 11727 1016 11728 1080
rect 11662 1000 11728 1016
rect 11662 936 11663 1000
rect 11727 936 11728 1000
rect 11662 920 11728 936
rect 11662 856 11663 920
rect 11727 856 11728 920
rect 11662 766 11728 856
rect 11788 702 11848 1732
rect 11908 762 11968 1794
rect 12028 702 12088 1732
rect 12148 762 12208 1794
rect 12268 1640 12334 1794
rect 12268 1576 12269 1640
rect 12333 1576 12334 1640
rect 12268 1560 12334 1576
rect 12268 1496 12269 1560
rect 12333 1496 12334 1560
rect 12268 1480 12334 1496
rect 12268 1416 12269 1480
rect 12333 1416 12334 1480
rect 12268 1400 12334 1416
rect 12268 1336 12269 1400
rect 12333 1336 12334 1400
rect 12268 1320 12334 1336
rect 12268 1256 12269 1320
rect 12333 1256 12334 1320
rect 12268 1240 12334 1256
rect 12268 1176 12269 1240
rect 12333 1176 12334 1240
rect 12268 1160 12334 1176
rect 12268 1096 12269 1160
rect 12333 1096 12334 1160
rect 12268 1080 12334 1096
rect 12268 1016 12269 1080
rect 12333 1016 12334 1080
rect 12268 1000 12334 1016
rect 12268 936 12269 1000
rect 12333 936 12334 1000
rect 12268 920 12334 936
rect 12268 856 12269 920
rect 12333 856 12334 920
rect 12268 766 12334 856
rect 12394 1860 12505 1862
rect 12569 1862 12578 1884
rect 13216 1885 13342 1895
rect 12569 1860 13066 1862
rect 12394 1796 12498 1860
rect 12569 1820 12578 1860
rect 12562 1796 12578 1820
rect 12642 1796 12658 1860
rect 12722 1796 12738 1860
rect 12802 1796 12818 1860
rect 12882 1796 12898 1860
rect 12962 1796 13066 1860
rect 13216 1821 13247 1885
rect 13311 1821 13342 1885
rect 13216 1811 13342 1821
rect 13242 1810 13316 1811
rect 12394 1794 13066 1796
rect 12394 1640 12460 1794
rect 12394 1576 12395 1640
rect 12459 1576 12460 1640
rect 12394 1560 12460 1576
rect 12394 1496 12395 1560
rect 12459 1496 12460 1560
rect 12394 1480 12460 1496
rect 12394 1416 12395 1480
rect 12459 1416 12460 1480
rect 12394 1400 12460 1416
rect 12394 1336 12395 1400
rect 12459 1336 12460 1400
rect 12394 1320 12460 1336
rect 12394 1256 12395 1320
rect 12459 1256 12460 1320
rect 12394 1240 12460 1256
rect 12394 1176 12395 1240
rect 12459 1176 12460 1240
rect 12394 1160 12460 1176
rect 12394 1096 12395 1160
rect 12459 1096 12460 1160
rect 12394 1080 12460 1096
rect 12394 1016 12395 1080
rect 12459 1016 12460 1080
rect 12394 1000 12460 1016
rect 12394 936 12395 1000
rect 12459 936 12460 1000
rect 12394 920 12460 936
rect 12394 856 12395 920
rect 12459 856 12460 920
rect 12394 766 12460 856
rect 12520 702 12580 1732
rect 12640 762 12700 1794
rect 12760 702 12820 1732
rect 12880 762 12940 1794
rect 13000 1640 13066 1794
rect 13000 1576 13001 1640
rect 13065 1576 13066 1640
rect 13000 1560 13066 1576
rect 13000 1496 13001 1560
rect 13065 1496 13066 1560
rect 13126 1623 13251 1633
rect 13126 1559 13156 1623
rect 13220 1559 13251 1623
rect 13126 1549 13251 1559
rect 13000 1480 13066 1496
rect 13000 1416 13001 1480
rect 13065 1416 13066 1480
rect 13000 1400 13066 1416
rect 13000 1336 13001 1400
rect 13065 1336 13066 1400
rect 13000 1320 13066 1336
rect 13000 1256 13001 1320
rect 13065 1256 13066 1320
rect 13000 1240 13066 1256
rect 13000 1176 13001 1240
rect 13065 1176 13066 1240
rect 13000 1160 13066 1176
rect 13000 1096 13001 1160
rect 13065 1096 13066 1160
rect 13000 1080 13066 1096
rect 13000 1016 13001 1080
rect 13065 1016 13066 1080
rect 13000 1000 13066 1016
rect 13000 936 13001 1000
rect 13065 936 13066 1000
rect 13000 920 13066 936
rect 13000 856 13001 920
rect 13065 856 13066 920
rect 13000 766 13066 856
rect 7383 634 7413 698
rect 7477 634 7508 698
rect 7774 700 8446 702
rect 7774 636 7878 700
rect 7942 636 7958 700
rect 8022 636 8038 700
rect 8102 636 8118 700
rect 8182 636 8198 700
rect 8262 636 8278 700
rect 8342 636 8446 700
rect 7774 634 8446 636
rect 8506 700 10996 702
rect 8506 636 8610 700
rect 8674 636 8690 700
rect 8754 636 8770 700
rect 8834 636 8850 700
rect 8914 636 8930 700
rect 8994 636 9010 700
rect 9074 636 9216 700
rect 9280 636 9296 700
rect 9360 636 9376 700
rect 9440 636 9456 700
rect 9520 636 9536 700
rect 9600 636 9616 700
rect 9680 636 9822 700
rect 9886 636 9902 700
rect 9966 636 9982 700
rect 10046 636 10062 700
rect 10126 636 10142 700
rect 10206 636 10222 700
rect 10286 636 10428 700
rect 10492 636 10508 700
rect 10572 636 10588 700
rect 10652 636 10668 700
rect 10732 636 10748 700
rect 10812 636 10828 700
rect 10892 636 10996 700
rect 8506 634 10996 636
rect 11056 700 12334 702
rect 11056 636 11160 700
rect 11224 636 11240 700
rect 11304 636 11320 700
rect 11384 636 11400 700
rect 11464 636 11480 700
rect 11544 636 11560 700
rect 11624 636 11766 700
rect 11830 636 11846 700
rect 11910 636 11926 700
rect 11990 636 12006 700
rect 12070 636 12086 700
rect 12150 636 12166 700
rect 12230 636 12334 700
rect 11056 634 12334 636
rect 12394 700 13066 702
rect 12394 636 12498 700
rect 12562 636 12578 700
rect 12642 636 12658 700
rect 12722 636 12738 700
rect 12802 636 12818 700
rect 12882 636 12898 700
rect 12962 636 13066 700
rect 12394 634 13066 636
rect 694 624 819 634
rect 7383 624 7508 634
rect 6030 314 6155 324
rect 12785 314 12910 324
rect 472 312 1144 314
rect 472 248 576 312
rect 640 248 656 312
rect 720 248 736 312
rect 800 248 816 312
rect 880 248 896 312
rect 960 248 976 312
rect 1040 248 1144 312
rect 472 246 1144 248
rect 1204 312 2482 314
rect 1204 248 1308 312
rect 1372 248 1388 312
rect 1452 248 1468 312
rect 1532 248 1548 312
rect 1612 248 1628 312
rect 1692 248 1708 312
rect 1772 248 1914 312
rect 1978 248 1994 312
rect 2058 248 2074 312
rect 2138 248 2154 312
rect 2218 248 2234 312
rect 2298 248 2314 312
rect 2378 248 2482 312
rect 1204 246 2482 248
rect 2542 312 5032 314
rect 2542 248 2646 312
rect 2710 248 2726 312
rect 2790 248 2806 312
rect 2870 248 2886 312
rect 2950 248 2966 312
rect 3030 248 3046 312
rect 3110 248 3252 312
rect 3316 248 3332 312
rect 3396 248 3412 312
rect 3476 248 3492 312
rect 3556 248 3572 312
rect 3636 248 3652 312
rect 3716 248 3858 312
rect 3922 248 3938 312
rect 4002 248 4018 312
rect 4082 248 4098 312
rect 4162 248 4178 312
rect 4242 248 4258 312
rect 4322 248 4464 312
rect 4528 248 4544 312
rect 4608 248 4624 312
rect 4688 248 4704 312
rect 4768 248 4784 312
rect 4848 248 4864 312
rect 4928 248 5032 312
rect 2542 246 5032 248
rect 5092 312 5764 314
rect 5092 248 5196 312
rect 5260 248 5276 312
rect 5340 248 5356 312
rect 5420 248 5436 312
rect 5500 248 5516 312
rect 5580 248 5596 312
rect 5660 248 5764 312
rect 5092 246 5764 248
rect 6030 250 6061 314
rect 6125 250 6155 314
rect 472 92 538 182
rect 472 28 473 92
rect 537 28 538 92
rect 472 12 538 28
rect 472 -52 473 12
rect 537 -52 538 12
rect 472 -68 538 -52
rect 472 -132 473 -68
rect 537 -132 538 -68
rect 472 -148 538 -132
rect 472 -212 473 -148
rect 537 -212 538 -148
rect 472 -228 538 -212
rect 472 -292 473 -228
rect 537 -292 538 -228
rect 472 -308 538 -292
rect 472 -372 473 -308
rect 537 -372 538 -308
rect 472 -388 538 -372
rect 472 -452 473 -388
rect 537 -452 538 -388
rect 472 -468 538 -452
rect 472 -532 473 -468
rect 537 -532 538 -468
rect 472 -548 538 -532
rect 287 -611 412 -601
rect 287 -675 318 -611
rect 382 -675 412 -611
rect 287 -685 412 -675
rect 472 -612 473 -548
rect 537 -612 538 -548
rect 472 -628 538 -612
rect 472 -692 473 -628
rect 537 -692 538 -628
rect 472 -846 538 -692
rect 598 -846 658 186
rect 718 -784 778 246
rect 838 -846 898 186
rect 958 -784 1018 246
rect 1078 92 1144 182
rect 1078 28 1079 92
rect 1143 28 1144 92
rect 1078 12 1144 28
rect 1078 -52 1079 12
rect 1143 -52 1144 12
rect 1078 -68 1144 -52
rect 1078 -132 1079 -68
rect 1143 -132 1144 -68
rect 1078 -148 1144 -132
rect 1078 -212 1079 -148
rect 1143 -212 1144 -148
rect 1078 -228 1144 -212
rect 1078 -292 1079 -228
rect 1143 -292 1144 -228
rect 1078 -308 1144 -292
rect 1078 -372 1079 -308
rect 1143 -372 1144 -308
rect 1078 -388 1144 -372
rect 1078 -452 1079 -388
rect 1143 -452 1144 -388
rect 1078 -468 1144 -452
rect 1078 -532 1079 -468
rect 1143 -532 1144 -468
rect 1078 -548 1144 -532
rect 1078 -612 1079 -548
rect 1143 -612 1144 -548
rect 1078 -628 1144 -612
rect 1078 -692 1079 -628
rect 1143 -692 1144 -628
rect 1078 -846 1144 -692
rect 472 -848 1144 -846
rect 222 -863 296 -862
rect 196 -873 322 -863
rect 196 -937 227 -873
rect 291 -937 322 -873
rect 472 -912 576 -848
rect 640 -912 656 -848
rect 720 -912 736 -848
rect 800 -912 816 -848
rect 880 -912 896 -848
rect 960 -872 976 -848
rect 960 -912 969 -872
rect 1040 -912 1144 -848
rect 472 -914 969 -912
rect 196 -947 322 -937
rect 960 -936 969 -914
rect 1033 -914 1144 -912
rect 1204 92 1270 182
rect 1204 28 1205 92
rect 1269 28 1270 92
rect 1204 12 1270 28
rect 1204 -52 1205 12
rect 1269 -52 1270 12
rect 1204 -68 1270 -52
rect 1204 -132 1205 -68
rect 1269 -132 1270 -68
rect 1204 -148 1270 -132
rect 1204 -212 1205 -148
rect 1269 -212 1270 -148
rect 1204 -228 1270 -212
rect 1204 -292 1205 -228
rect 1269 -292 1270 -228
rect 1204 -308 1270 -292
rect 1204 -372 1205 -308
rect 1269 -372 1270 -308
rect 1204 -388 1270 -372
rect 1204 -452 1205 -388
rect 1269 -452 1270 -388
rect 1204 -468 1270 -452
rect 1204 -532 1205 -468
rect 1269 -532 1270 -468
rect 1204 -548 1270 -532
rect 1204 -612 1205 -548
rect 1269 -612 1270 -548
rect 1204 -628 1270 -612
rect 1204 -692 1205 -628
rect 1269 -692 1270 -628
rect 1204 -846 1270 -692
rect 1330 -846 1390 186
rect 1450 -784 1510 246
rect 1570 -846 1630 186
rect 1690 -784 1750 246
rect 1810 92 1876 182
rect 1810 28 1811 92
rect 1875 28 1876 92
rect 1810 12 1876 28
rect 1810 -52 1811 12
rect 1875 -52 1876 12
rect 1810 -68 1876 -52
rect 1810 -132 1811 -68
rect 1875 -132 1876 -68
rect 1810 -148 1876 -132
rect 1810 -212 1811 -148
rect 1875 -212 1876 -148
rect 1810 -228 1876 -212
rect 1810 -292 1811 -228
rect 1875 -292 1876 -228
rect 1810 -308 1876 -292
rect 1810 -372 1811 -308
rect 1875 -372 1876 -308
rect 1810 -388 1876 -372
rect 1810 -452 1811 -388
rect 1875 -452 1876 -388
rect 1810 -468 1876 -452
rect 1810 -532 1811 -468
rect 1875 -532 1876 -468
rect 1810 -548 1876 -532
rect 1810 -612 1811 -548
rect 1875 -612 1876 -548
rect 1810 -628 1876 -612
rect 1810 -692 1811 -628
rect 1875 -692 1876 -628
rect 1810 -846 1876 -692
rect 1936 -784 1996 246
rect 2056 -846 2116 186
rect 2176 -784 2236 246
rect 2296 -846 2356 186
rect 2416 92 2482 182
rect 2416 28 2417 92
rect 2481 28 2482 92
rect 2416 12 2482 28
rect 2416 -52 2417 12
rect 2481 -52 2482 12
rect 2416 -68 2482 -52
rect 2416 -132 2417 -68
rect 2481 -132 2482 -68
rect 2416 -148 2482 -132
rect 2416 -212 2417 -148
rect 2481 -212 2482 -148
rect 2416 -228 2482 -212
rect 2416 -292 2417 -228
rect 2481 -292 2482 -228
rect 2416 -308 2482 -292
rect 2416 -372 2417 -308
rect 2481 -372 2482 -308
rect 2416 -388 2482 -372
rect 2416 -452 2417 -388
rect 2481 -452 2482 -388
rect 2416 -468 2482 -452
rect 2416 -532 2417 -468
rect 2481 -532 2482 -468
rect 2416 -548 2482 -532
rect 2416 -612 2417 -548
rect 2481 -612 2482 -548
rect 2416 -628 2482 -612
rect 2416 -692 2417 -628
rect 2481 -692 2482 -628
rect 2416 -846 2482 -692
rect 1204 -848 2482 -846
rect 1204 -912 1308 -848
rect 1372 -912 1388 -848
rect 1452 -912 1468 -848
rect 1532 -912 1548 -848
rect 1612 -912 1628 -848
rect 1692 -872 1708 -848
rect 1692 -912 1701 -872
rect 1772 -912 1914 -848
rect 1978 -872 1994 -848
rect 1985 -912 1994 -872
rect 2058 -912 2074 -848
rect 2138 -912 2154 -848
rect 2218 -912 2234 -848
rect 2298 -912 2314 -848
rect 2378 -912 2482 -848
rect 1204 -914 1701 -912
rect 1033 -936 1042 -914
rect 960 -942 1042 -936
rect 1692 -936 1701 -914
rect 1765 -914 1921 -912
rect 1765 -936 1774 -914
rect 1692 -942 1774 -936
rect 1912 -936 1921 -914
rect 1985 -914 2482 -912
rect 2542 92 2608 182
rect 2542 28 2543 92
rect 2607 28 2608 92
rect 2542 12 2608 28
rect 2542 -52 2543 12
rect 2607 -52 2608 12
rect 2542 -68 2608 -52
rect 2542 -132 2543 -68
rect 2607 -132 2608 -68
rect 2542 -148 2608 -132
rect 2542 -212 2543 -148
rect 2607 -212 2608 -148
rect 2542 -228 2608 -212
rect 2542 -292 2543 -228
rect 2607 -292 2608 -228
rect 2542 -308 2608 -292
rect 2542 -372 2543 -308
rect 2607 -372 2608 -308
rect 2542 -388 2608 -372
rect 2542 -452 2543 -388
rect 2607 -452 2608 -388
rect 2542 -468 2608 -452
rect 2542 -532 2543 -468
rect 2607 -532 2608 -468
rect 2542 -548 2608 -532
rect 2542 -612 2543 -548
rect 2607 -612 2608 -548
rect 2542 -628 2608 -612
rect 2542 -692 2543 -628
rect 2607 -692 2608 -628
rect 2542 -846 2608 -692
rect 2668 -846 2728 186
rect 2788 -784 2848 246
rect 2908 -846 2968 186
rect 3028 -784 3088 246
rect 3148 92 3214 182
rect 3148 28 3149 92
rect 3213 28 3214 92
rect 3148 12 3214 28
rect 3148 -52 3149 12
rect 3213 -52 3214 12
rect 3148 -68 3214 -52
rect 3148 -132 3149 -68
rect 3213 -132 3214 -68
rect 3148 -148 3214 -132
rect 3148 -212 3149 -148
rect 3213 -212 3214 -148
rect 3148 -228 3214 -212
rect 3148 -292 3149 -228
rect 3213 -292 3214 -228
rect 3148 -308 3214 -292
rect 3148 -372 3149 -308
rect 3213 -372 3214 -308
rect 3148 -388 3214 -372
rect 3148 -452 3149 -388
rect 3213 -452 3214 -388
rect 3148 -468 3214 -452
rect 3148 -532 3149 -468
rect 3213 -532 3214 -468
rect 3148 -548 3214 -532
rect 3148 -612 3149 -548
rect 3213 -612 3214 -548
rect 3148 -628 3214 -612
rect 3148 -692 3149 -628
rect 3213 -692 3214 -628
rect 3148 -846 3214 -692
rect 3274 -784 3334 246
rect 3394 -846 3454 186
rect 3514 -784 3574 246
rect 3634 -846 3694 186
rect 3754 92 3820 182
rect 3754 28 3755 92
rect 3819 28 3820 92
rect 3754 12 3820 28
rect 3754 -52 3755 12
rect 3819 -52 3820 12
rect 3754 -68 3820 -52
rect 3754 -132 3755 -68
rect 3819 -132 3820 -68
rect 3754 -148 3820 -132
rect 3754 -212 3755 -148
rect 3819 -212 3820 -148
rect 3754 -228 3820 -212
rect 3754 -292 3755 -228
rect 3819 -292 3820 -228
rect 3754 -308 3820 -292
rect 3754 -372 3755 -308
rect 3819 -372 3820 -308
rect 3754 -388 3820 -372
rect 3754 -452 3755 -388
rect 3819 -452 3820 -388
rect 3754 -468 3820 -452
rect 3754 -532 3755 -468
rect 3819 -532 3820 -468
rect 3754 -548 3820 -532
rect 3754 -612 3755 -548
rect 3819 -612 3820 -548
rect 3754 -628 3820 -612
rect 3754 -692 3755 -628
rect 3819 -692 3820 -628
rect 3754 -846 3820 -692
rect 3880 -846 3940 186
rect 4000 -784 4060 246
rect 4120 -846 4180 186
rect 4240 -784 4300 246
rect 4360 92 4426 182
rect 4360 28 4361 92
rect 4425 28 4426 92
rect 4360 12 4426 28
rect 4360 -52 4361 12
rect 4425 -52 4426 12
rect 4360 -68 4426 -52
rect 4360 -132 4361 -68
rect 4425 -132 4426 -68
rect 4360 -148 4426 -132
rect 4360 -212 4361 -148
rect 4425 -212 4426 -148
rect 4360 -228 4426 -212
rect 4360 -292 4361 -228
rect 4425 -292 4426 -228
rect 4360 -308 4426 -292
rect 4360 -372 4361 -308
rect 4425 -372 4426 -308
rect 4360 -388 4426 -372
rect 4360 -452 4361 -388
rect 4425 -452 4426 -388
rect 4360 -468 4426 -452
rect 4360 -532 4361 -468
rect 4425 -532 4426 -468
rect 4360 -548 4426 -532
rect 4360 -612 4361 -548
rect 4425 -612 4426 -548
rect 4360 -628 4426 -612
rect 4360 -692 4361 -628
rect 4425 -692 4426 -628
rect 4360 -846 4426 -692
rect 4486 -784 4546 246
rect 4606 -846 4666 186
rect 4726 -784 4786 246
rect 4846 -846 4906 186
rect 4966 92 5032 182
rect 4966 28 4967 92
rect 5031 28 5032 92
rect 4966 12 5032 28
rect 4966 -52 4967 12
rect 5031 -52 5032 12
rect 4966 -68 5032 -52
rect 4966 -132 4967 -68
rect 5031 -132 5032 -68
rect 4966 -148 5032 -132
rect 4966 -212 4967 -148
rect 5031 -212 5032 -148
rect 4966 -228 5032 -212
rect 4966 -292 4967 -228
rect 5031 -292 5032 -228
rect 4966 -308 5032 -292
rect 4966 -372 4967 -308
rect 5031 -372 5032 -308
rect 4966 -388 5032 -372
rect 4966 -452 4967 -388
rect 5031 -452 5032 -388
rect 4966 -468 5032 -452
rect 4966 -532 4967 -468
rect 5031 -532 5032 -468
rect 4966 -548 5032 -532
rect 4966 -612 4967 -548
rect 5031 -612 5032 -548
rect 4966 -628 5032 -612
rect 4966 -692 4967 -628
rect 5031 -692 5032 -628
rect 4966 -846 5032 -692
rect 2542 -848 5032 -846
rect 2542 -912 2646 -848
rect 2710 -912 2726 -848
rect 2790 -912 2806 -848
rect 2870 -912 2886 -848
rect 2950 -912 2966 -848
rect 3030 -872 3046 -848
rect 3030 -912 3039 -872
rect 3110 -912 3252 -848
rect 3316 -872 3332 -848
rect 3323 -912 3332 -872
rect 3396 -912 3412 -848
rect 3476 -912 3492 -848
rect 3556 -912 3572 -848
rect 3636 -912 3652 -848
rect 3716 -912 3858 -848
rect 3922 -912 3938 -848
rect 4002 -912 4018 -848
rect 4082 -912 4098 -848
rect 4162 -912 4178 -848
rect 4242 -872 4258 -848
rect 4242 -912 4251 -872
rect 4322 -912 4464 -848
rect 4528 -872 4544 -848
rect 4535 -912 4544 -872
rect 4608 -912 4624 -848
rect 4688 -912 4704 -848
rect 4768 -912 4784 -848
rect 4848 -912 4864 -848
rect 4928 -912 5032 -848
rect 2542 -914 3039 -912
rect 1985 -936 1994 -914
rect 1912 -942 1994 -936
rect 3030 -936 3039 -914
rect 3103 -914 3259 -912
rect 3103 -936 3112 -914
rect 3030 -942 3112 -936
rect 3250 -936 3259 -914
rect 3323 -914 4251 -912
rect 3323 -936 3332 -914
rect 3250 -942 3332 -936
rect 4242 -936 4251 -914
rect 4315 -914 4471 -912
rect 4315 -936 4324 -914
rect 4242 -942 4324 -936
rect 4462 -936 4471 -914
rect 4535 -914 5032 -912
rect 5092 92 5158 182
rect 5092 28 5093 92
rect 5157 28 5158 92
rect 5092 12 5158 28
rect 5092 -52 5093 12
rect 5157 -52 5158 12
rect 5092 -68 5158 -52
rect 5092 -132 5093 -68
rect 5157 -132 5158 -68
rect 5092 -148 5158 -132
rect 5092 -212 5093 -148
rect 5157 -212 5158 -148
rect 5092 -228 5158 -212
rect 5092 -292 5093 -228
rect 5157 -292 5158 -228
rect 5092 -308 5158 -292
rect 5092 -372 5093 -308
rect 5157 -372 5158 -308
rect 5092 -388 5158 -372
rect 5092 -452 5093 -388
rect 5157 -452 5158 -388
rect 5092 -468 5158 -452
rect 5092 -532 5093 -468
rect 5157 -532 5158 -468
rect 5092 -548 5158 -532
rect 5092 -612 5093 -548
rect 5157 -612 5158 -548
rect 5092 -628 5158 -612
rect 5092 -692 5093 -628
rect 5157 -692 5158 -628
rect 5092 -846 5158 -692
rect 5218 -784 5278 246
rect 5338 -846 5398 186
rect 5458 -784 5518 246
rect 6030 240 6155 250
rect 7227 312 7899 314
rect 7227 248 7331 312
rect 7395 248 7411 312
rect 7475 248 7491 312
rect 7555 248 7571 312
rect 7635 248 7651 312
rect 7715 248 7731 312
rect 7795 248 7899 312
rect 7227 246 7899 248
rect 7959 312 9237 314
rect 7959 248 8063 312
rect 8127 248 8143 312
rect 8207 248 8223 312
rect 8287 248 8303 312
rect 8367 248 8383 312
rect 8447 248 8463 312
rect 8527 248 8669 312
rect 8733 248 8749 312
rect 8813 248 8829 312
rect 8893 248 8909 312
rect 8973 248 8989 312
rect 9053 248 9069 312
rect 9133 248 9237 312
rect 7959 246 9237 248
rect 9297 312 11787 314
rect 9297 248 9401 312
rect 9465 248 9481 312
rect 9545 248 9561 312
rect 9625 248 9641 312
rect 9705 248 9721 312
rect 9785 248 9801 312
rect 9865 248 10007 312
rect 10071 248 10087 312
rect 10151 248 10167 312
rect 10231 248 10247 312
rect 10311 248 10327 312
rect 10391 248 10407 312
rect 10471 248 10613 312
rect 10677 248 10693 312
rect 10757 248 10773 312
rect 10837 248 10853 312
rect 10917 248 10933 312
rect 10997 248 11013 312
rect 11077 248 11219 312
rect 11283 248 11299 312
rect 11363 248 11379 312
rect 11443 248 11459 312
rect 11523 248 11539 312
rect 11603 248 11619 312
rect 11683 248 11787 312
rect 9297 246 11787 248
rect 11847 312 12519 314
rect 11847 248 11951 312
rect 12015 248 12031 312
rect 12095 248 12111 312
rect 12175 248 12191 312
rect 12255 248 12271 312
rect 12335 248 12351 312
rect 12415 248 12519 312
rect 11847 246 12519 248
rect 12785 250 12816 314
rect 12880 250 12910 314
rect 5578 -846 5638 186
rect 5698 92 5764 182
rect 5698 28 5699 92
rect 5763 28 5764 92
rect 5698 12 5764 28
rect 5698 -52 5699 12
rect 5763 -52 5764 12
rect 5698 -68 5764 -52
rect 5698 -132 5699 -68
rect 5763 -132 5764 -68
rect 5698 -148 5764 -132
rect 5698 -212 5699 -148
rect 5763 -212 5764 -148
rect 5698 -228 5764 -212
rect 5698 -292 5699 -228
rect 5763 -292 5764 -228
rect 5698 -308 5764 -292
rect 5698 -372 5699 -308
rect 5763 -372 5764 -308
rect 5698 -388 5764 -372
rect 5698 -452 5699 -388
rect 5763 -452 5764 -388
rect 5698 -468 5764 -452
rect 5698 -532 5699 -468
rect 5763 -532 5764 -468
rect 5698 -548 5764 -532
rect 5698 -612 5699 -548
rect 5763 -612 5764 -548
rect 7227 92 7293 182
rect 7227 28 7228 92
rect 7292 28 7293 92
rect 7227 12 7293 28
rect 7227 -52 7228 12
rect 7292 -52 7293 12
rect 7227 -68 7293 -52
rect 7227 -132 7228 -68
rect 7292 -132 7293 -68
rect 7227 -148 7293 -132
rect 7227 -212 7228 -148
rect 7292 -212 7293 -148
rect 7227 -228 7293 -212
rect 7227 -292 7228 -228
rect 7292 -292 7293 -228
rect 7227 -308 7293 -292
rect 7227 -372 7228 -308
rect 7292 -372 7293 -308
rect 7227 -388 7293 -372
rect 7227 -452 7228 -388
rect 7292 -452 7293 -388
rect 7227 -468 7293 -452
rect 7227 -532 7228 -468
rect 7292 -532 7293 -468
rect 7227 -548 7293 -532
rect 5698 -628 5764 -612
rect 5698 -692 5699 -628
rect 5763 -692 5764 -628
rect 7042 -611 7167 -601
rect 7042 -675 7073 -611
rect 7137 -675 7167 -611
rect 7042 -685 7167 -675
rect 7227 -612 7228 -548
rect 7292 -612 7293 -548
rect 7227 -628 7293 -612
rect 5698 -846 5764 -692
rect 5092 -848 5764 -846
rect 5092 -912 5196 -848
rect 5260 -872 5276 -848
rect 5267 -912 5276 -872
rect 5340 -912 5356 -848
rect 5420 -912 5436 -848
rect 5500 -912 5516 -848
rect 5580 -912 5596 -848
rect 5660 -912 5764 -848
rect 7227 -692 7228 -628
rect 7292 -692 7293 -628
rect 7227 -846 7293 -692
rect 7353 -846 7413 186
rect 7473 -784 7533 246
rect 7593 -846 7653 186
rect 7713 -784 7773 246
rect 7833 92 7899 182
rect 7833 28 7834 92
rect 7898 28 7899 92
rect 7833 12 7899 28
rect 7833 -52 7834 12
rect 7898 -52 7899 12
rect 7833 -68 7899 -52
rect 7833 -132 7834 -68
rect 7898 -132 7899 -68
rect 7833 -148 7899 -132
rect 7833 -212 7834 -148
rect 7898 -212 7899 -148
rect 7833 -228 7899 -212
rect 7833 -292 7834 -228
rect 7898 -292 7899 -228
rect 7833 -308 7899 -292
rect 7833 -372 7834 -308
rect 7898 -372 7899 -308
rect 7833 -388 7899 -372
rect 7833 -452 7834 -388
rect 7898 -452 7899 -388
rect 7833 -468 7899 -452
rect 7833 -532 7834 -468
rect 7898 -532 7899 -468
rect 7833 -548 7899 -532
rect 7833 -612 7834 -548
rect 7898 -612 7899 -548
rect 7833 -628 7899 -612
rect 7833 -692 7834 -628
rect 7898 -692 7899 -628
rect 7833 -846 7899 -692
rect 7227 -848 7899 -846
rect 6977 -863 7051 -862
rect 5092 -914 5203 -912
rect 4535 -936 4544 -914
rect 4462 -942 4544 -936
rect 5194 -936 5203 -914
rect 5267 -914 5764 -912
rect 6951 -873 7077 -863
rect 5267 -936 5276 -914
rect 5194 -942 5276 -936
rect 6951 -937 6982 -873
rect 7046 -937 7077 -873
rect 7227 -912 7331 -848
rect 7395 -912 7411 -848
rect 7475 -912 7491 -848
rect 7555 -912 7571 -848
rect 7635 -912 7651 -848
rect 7715 -872 7731 -848
rect 7715 -912 7724 -872
rect 7795 -912 7899 -848
rect 7227 -914 7724 -912
rect 6951 -947 7077 -937
rect 7715 -936 7724 -914
rect 7788 -914 7899 -912
rect 7959 92 8025 182
rect 7959 28 7960 92
rect 8024 28 8025 92
rect 7959 12 8025 28
rect 7959 -52 7960 12
rect 8024 -52 8025 12
rect 7959 -68 8025 -52
rect 7959 -132 7960 -68
rect 8024 -132 8025 -68
rect 7959 -148 8025 -132
rect 7959 -212 7960 -148
rect 8024 -212 8025 -148
rect 7959 -228 8025 -212
rect 7959 -292 7960 -228
rect 8024 -292 8025 -228
rect 7959 -308 8025 -292
rect 7959 -372 7960 -308
rect 8024 -372 8025 -308
rect 7959 -388 8025 -372
rect 7959 -452 7960 -388
rect 8024 -452 8025 -388
rect 7959 -468 8025 -452
rect 7959 -532 7960 -468
rect 8024 -532 8025 -468
rect 7959 -548 8025 -532
rect 7959 -612 7960 -548
rect 8024 -612 8025 -548
rect 7959 -628 8025 -612
rect 7959 -692 7960 -628
rect 8024 -692 8025 -628
rect 7959 -846 8025 -692
rect 8085 -846 8145 186
rect 8205 -784 8265 246
rect 8325 -846 8385 186
rect 8445 -784 8505 246
rect 8565 92 8631 182
rect 8565 28 8566 92
rect 8630 28 8631 92
rect 8565 12 8631 28
rect 8565 -52 8566 12
rect 8630 -52 8631 12
rect 8565 -68 8631 -52
rect 8565 -132 8566 -68
rect 8630 -132 8631 -68
rect 8565 -148 8631 -132
rect 8565 -212 8566 -148
rect 8630 -212 8631 -148
rect 8565 -228 8631 -212
rect 8565 -292 8566 -228
rect 8630 -292 8631 -228
rect 8565 -308 8631 -292
rect 8565 -372 8566 -308
rect 8630 -372 8631 -308
rect 8565 -388 8631 -372
rect 8565 -452 8566 -388
rect 8630 -452 8631 -388
rect 8565 -468 8631 -452
rect 8565 -532 8566 -468
rect 8630 -532 8631 -468
rect 8565 -548 8631 -532
rect 8565 -612 8566 -548
rect 8630 -612 8631 -548
rect 8565 -628 8631 -612
rect 8565 -692 8566 -628
rect 8630 -692 8631 -628
rect 8565 -846 8631 -692
rect 8691 -784 8751 246
rect 8811 -846 8871 186
rect 8931 -784 8991 246
rect 9051 -846 9111 186
rect 9171 92 9237 182
rect 9171 28 9172 92
rect 9236 28 9237 92
rect 9171 12 9237 28
rect 9171 -52 9172 12
rect 9236 -52 9237 12
rect 9171 -68 9237 -52
rect 9171 -132 9172 -68
rect 9236 -132 9237 -68
rect 9171 -148 9237 -132
rect 9171 -212 9172 -148
rect 9236 -212 9237 -148
rect 9171 -228 9237 -212
rect 9171 -292 9172 -228
rect 9236 -292 9237 -228
rect 9171 -308 9237 -292
rect 9171 -372 9172 -308
rect 9236 -372 9237 -308
rect 9171 -388 9237 -372
rect 9171 -452 9172 -388
rect 9236 -452 9237 -388
rect 9171 -468 9237 -452
rect 9171 -532 9172 -468
rect 9236 -532 9237 -468
rect 9171 -548 9237 -532
rect 9171 -612 9172 -548
rect 9236 -612 9237 -548
rect 9171 -628 9237 -612
rect 9171 -692 9172 -628
rect 9236 -692 9237 -628
rect 9171 -846 9237 -692
rect 7959 -848 9237 -846
rect 7959 -912 8063 -848
rect 8127 -912 8143 -848
rect 8207 -912 8223 -848
rect 8287 -912 8303 -848
rect 8367 -912 8383 -848
rect 8447 -872 8463 -848
rect 8447 -912 8456 -872
rect 8527 -912 8669 -848
rect 8733 -872 8749 -848
rect 8740 -912 8749 -872
rect 8813 -912 8829 -848
rect 8893 -912 8909 -848
rect 8973 -912 8989 -848
rect 9053 -912 9069 -848
rect 9133 -912 9237 -848
rect 7959 -914 8456 -912
rect 7788 -936 7797 -914
rect 7715 -942 7797 -936
rect 8447 -936 8456 -914
rect 8520 -914 8676 -912
rect 8520 -936 8529 -914
rect 8447 -942 8529 -936
rect 8667 -936 8676 -914
rect 8740 -914 9237 -912
rect 9297 92 9363 182
rect 9297 28 9298 92
rect 9362 28 9363 92
rect 9297 12 9363 28
rect 9297 -52 9298 12
rect 9362 -52 9363 12
rect 9297 -68 9363 -52
rect 9297 -132 9298 -68
rect 9362 -132 9363 -68
rect 9297 -148 9363 -132
rect 9297 -212 9298 -148
rect 9362 -212 9363 -148
rect 9297 -228 9363 -212
rect 9297 -292 9298 -228
rect 9362 -292 9363 -228
rect 9297 -308 9363 -292
rect 9297 -372 9298 -308
rect 9362 -372 9363 -308
rect 9297 -388 9363 -372
rect 9297 -452 9298 -388
rect 9362 -452 9363 -388
rect 9297 -468 9363 -452
rect 9297 -532 9298 -468
rect 9362 -532 9363 -468
rect 9297 -548 9363 -532
rect 9297 -612 9298 -548
rect 9362 -612 9363 -548
rect 9297 -628 9363 -612
rect 9297 -692 9298 -628
rect 9362 -692 9363 -628
rect 9297 -846 9363 -692
rect 9423 -846 9483 186
rect 9543 -784 9603 246
rect 9663 -846 9723 186
rect 9783 -784 9843 246
rect 9903 92 9969 182
rect 9903 28 9904 92
rect 9968 28 9969 92
rect 9903 12 9969 28
rect 9903 -52 9904 12
rect 9968 -52 9969 12
rect 9903 -68 9969 -52
rect 9903 -132 9904 -68
rect 9968 -132 9969 -68
rect 9903 -148 9969 -132
rect 9903 -212 9904 -148
rect 9968 -212 9969 -148
rect 9903 -228 9969 -212
rect 9903 -292 9904 -228
rect 9968 -292 9969 -228
rect 9903 -308 9969 -292
rect 9903 -372 9904 -308
rect 9968 -372 9969 -308
rect 9903 -388 9969 -372
rect 9903 -452 9904 -388
rect 9968 -452 9969 -388
rect 9903 -468 9969 -452
rect 9903 -532 9904 -468
rect 9968 -532 9969 -468
rect 9903 -548 9969 -532
rect 9903 -612 9904 -548
rect 9968 -612 9969 -548
rect 9903 -628 9969 -612
rect 9903 -692 9904 -628
rect 9968 -692 9969 -628
rect 9903 -846 9969 -692
rect 10029 -784 10089 246
rect 10149 -846 10209 186
rect 10269 -784 10329 246
rect 10389 -846 10449 186
rect 10509 92 10575 182
rect 10509 28 10510 92
rect 10574 28 10575 92
rect 10509 12 10575 28
rect 10509 -52 10510 12
rect 10574 -52 10575 12
rect 10509 -68 10575 -52
rect 10509 -132 10510 -68
rect 10574 -132 10575 -68
rect 10509 -148 10575 -132
rect 10509 -212 10510 -148
rect 10574 -212 10575 -148
rect 10509 -228 10575 -212
rect 10509 -292 10510 -228
rect 10574 -292 10575 -228
rect 10509 -308 10575 -292
rect 10509 -372 10510 -308
rect 10574 -372 10575 -308
rect 10509 -388 10575 -372
rect 10509 -452 10510 -388
rect 10574 -452 10575 -388
rect 10509 -468 10575 -452
rect 10509 -532 10510 -468
rect 10574 -532 10575 -468
rect 10509 -548 10575 -532
rect 10509 -612 10510 -548
rect 10574 -612 10575 -548
rect 10509 -628 10575 -612
rect 10509 -692 10510 -628
rect 10574 -692 10575 -628
rect 10509 -846 10575 -692
rect 10635 -846 10695 186
rect 10755 -784 10815 246
rect 10875 -846 10935 186
rect 10995 -784 11055 246
rect 11115 92 11181 182
rect 11115 28 11116 92
rect 11180 28 11181 92
rect 11115 12 11181 28
rect 11115 -52 11116 12
rect 11180 -52 11181 12
rect 11115 -68 11181 -52
rect 11115 -132 11116 -68
rect 11180 -132 11181 -68
rect 11115 -148 11181 -132
rect 11115 -212 11116 -148
rect 11180 -212 11181 -148
rect 11115 -228 11181 -212
rect 11115 -292 11116 -228
rect 11180 -292 11181 -228
rect 11115 -308 11181 -292
rect 11115 -372 11116 -308
rect 11180 -372 11181 -308
rect 11115 -388 11181 -372
rect 11115 -452 11116 -388
rect 11180 -452 11181 -388
rect 11115 -468 11181 -452
rect 11115 -532 11116 -468
rect 11180 -532 11181 -468
rect 11115 -548 11181 -532
rect 11115 -612 11116 -548
rect 11180 -612 11181 -548
rect 11115 -628 11181 -612
rect 11115 -692 11116 -628
rect 11180 -692 11181 -628
rect 11115 -846 11181 -692
rect 11241 -784 11301 246
rect 11361 -846 11421 186
rect 11481 -784 11541 246
rect 11601 -846 11661 186
rect 11721 92 11787 182
rect 11721 28 11722 92
rect 11786 28 11787 92
rect 11721 12 11787 28
rect 11721 -52 11722 12
rect 11786 -52 11787 12
rect 11721 -68 11787 -52
rect 11721 -132 11722 -68
rect 11786 -132 11787 -68
rect 11721 -148 11787 -132
rect 11721 -212 11722 -148
rect 11786 -212 11787 -148
rect 11721 -228 11787 -212
rect 11721 -292 11722 -228
rect 11786 -292 11787 -228
rect 11721 -308 11787 -292
rect 11721 -372 11722 -308
rect 11786 -372 11787 -308
rect 11721 -388 11787 -372
rect 11721 -452 11722 -388
rect 11786 -452 11787 -388
rect 11721 -468 11787 -452
rect 11721 -532 11722 -468
rect 11786 -532 11787 -468
rect 11721 -548 11787 -532
rect 11721 -612 11722 -548
rect 11786 -612 11787 -548
rect 11721 -628 11787 -612
rect 11721 -692 11722 -628
rect 11786 -692 11787 -628
rect 11721 -846 11787 -692
rect 9297 -848 11787 -846
rect 9297 -912 9401 -848
rect 9465 -912 9481 -848
rect 9545 -912 9561 -848
rect 9625 -912 9641 -848
rect 9705 -912 9721 -848
rect 9785 -872 9801 -848
rect 9785 -912 9794 -872
rect 9865 -912 10007 -848
rect 10071 -872 10087 -848
rect 10078 -912 10087 -872
rect 10151 -912 10167 -848
rect 10231 -912 10247 -848
rect 10311 -912 10327 -848
rect 10391 -912 10407 -848
rect 10471 -912 10613 -848
rect 10677 -912 10693 -848
rect 10757 -912 10773 -848
rect 10837 -912 10853 -848
rect 10917 -912 10933 -848
rect 10997 -872 11013 -848
rect 10997 -912 11006 -872
rect 11077 -912 11219 -848
rect 11283 -872 11299 -848
rect 11290 -912 11299 -872
rect 11363 -912 11379 -848
rect 11443 -912 11459 -848
rect 11523 -912 11539 -848
rect 11603 -912 11619 -848
rect 11683 -912 11787 -848
rect 9297 -914 9794 -912
rect 8740 -936 8749 -914
rect 8667 -942 8749 -936
rect 9785 -936 9794 -914
rect 9858 -914 10014 -912
rect 9858 -936 9867 -914
rect 9785 -942 9867 -936
rect 10005 -936 10014 -914
rect 10078 -914 11006 -912
rect 10078 -936 10087 -914
rect 10005 -942 10087 -936
rect 10997 -936 11006 -914
rect 11070 -914 11226 -912
rect 11070 -936 11079 -914
rect 10997 -942 11079 -936
rect 11217 -936 11226 -914
rect 11290 -914 11787 -912
rect 11847 92 11913 182
rect 11847 28 11848 92
rect 11912 28 11913 92
rect 11847 12 11913 28
rect 11847 -52 11848 12
rect 11912 -52 11913 12
rect 11847 -68 11913 -52
rect 11847 -132 11848 -68
rect 11912 -132 11913 -68
rect 11847 -148 11913 -132
rect 11847 -212 11848 -148
rect 11912 -212 11913 -148
rect 11847 -228 11913 -212
rect 11847 -292 11848 -228
rect 11912 -292 11913 -228
rect 11847 -308 11913 -292
rect 11847 -372 11848 -308
rect 11912 -372 11913 -308
rect 11847 -388 11913 -372
rect 11847 -452 11848 -388
rect 11912 -452 11913 -388
rect 11847 -468 11913 -452
rect 11847 -532 11848 -468
rect 11912 -532 11913 -468
rect 11847 -548 11913 -532
rect 11847 -612 11848 -548
rect 11912 -612 11913 -548
rect 11847 -628 11913 -612
rect 11847 -692 11848 -628
rect 11912 -692 11913 -628
rect 11847 -846 11913 -692
rect 11973 -784 12033 246
rect 12093 -846 12153 186
rect 12213 -784 12273 246
rect 12785 240 12910 250
rect 12333 -846 12393 186
rect 12453 92 12519 182
rect 12453 28 12454 92
rect 12518 28 12519 92
rect 12453 12 12519 28
rect 12453 -52 12454 12
rect 12518 -52 12519 12
rect 12453 -68 12519 -52
rect 12453 -132 12454 -68
rect 12518 -132 12519 -68
rect 12453 -148 12519 -132
rect 12453 -212 12454 -148
rect 12518 -212 12519 -148
rect 12453 -228 12519 -212
rect 12453 -292 12454 -228
rect 12518 -292 12519 -228
rect 12453 -308 12519 -292
rect 12453 -372 12454 -308
rect 12518 -372 12519 -308
rect 12453 -388 12519 -372
rect 12453 -452 12454 -388
rect 12518 -452 12519 -388
rect 12453 -468 12519 -452
rect 12453 -532 12454 -468
rect 12518 -532 12519 -468
rect 12453 -548 12519 -532
rect 12453 -612 12454 -548
rect 12518 -612 12519 -548
rect 12453 -628 12519 -612
rect 12453 -692 12454 -628
rect 12518 -692 12519 -628
rect 12453 -846 12519 -692
rect 11847 -848 12519 -846
rect 11847 -912 11951 -848
rect 12015 -872 12031 -848
rect 12022 -912 12031 -872
rect 12095 -912 12111 -848
rect 12175 -912 12191 -848
rect 12255 -912 12271 -848
rect 12335 -912 12351 -848
rect 12415 -912 12519 -848
rect 11847 -914 11958 -912
rect 11290 -936 11299 -914
rect 11217 -942 11299 -936
rect 11949 -936 11958 -914
rect 12022 -914 12519 -912
rect 12022 -936 12031 -914
rect 11949 -942 12031 -936
rect 196 -1076 322 -1066
rect 196 -1140 227 -1076
rect 291 -1140 322 -1076
rect 955 -1074 1038 -1069
rect 955 -1095 965 -1074
rect 196 -1150 322 -1140
rect 472 -1097 965 -1095
rect 1029 -1095 1038 -1074
rect 1184 -1074 1267 -1069
rect 1184 -1095 1193 -1074
rect 1029 -1097 1193 -1095
rect 1257 -1095 1267 -1074
rect 2167 -1074 2250 -1069
rect 2167 -1095 2177 -1074
rect 1257 -1097 2177 -1095
rect 2241 -1095 2250 -1074
rect 2396 -1074 2479 -1069
rect 2396 -1095 2405 -1074
rect 2241 -1097 2405 -1095
rect 2469 -1095 2479 -1074
rect 3379 -1074 3462 -1069
rect 3379 -1095 3389 -1074
rect 2469 -1097 3389 -1095
rect 3453 -1095 3462 -1074
rect 3608 -1074 3691 -1069
rect 3608 -1095 3617 -1074
rect 3453 -1097 3617 -1095
rect 3681 -1095 3691 -1074
rect 4591 -1074 4674 -1069
rect 4591 -1095 4601 -1074
rect 3681 -1097 4601 -1095
rect 4665 -1095 4674 -1074
rect 4820 -1074 4903 -1069
rect 4820 -1095 4829 -1074
rect 4665 -1097 4829 -1095
rect 4893 -1095 4903 -1074
rect 5552 -1074 5635 -1069
rect 5552 -1095 5561 -1074
rect 4893 -1097 5386 -1095
rect 472 -1161 576 -1097
rect 640 -1161 656 -1097
rect 720 -1161 736 -1097
rect 800 -1161 816 -1097
rect 880 -1161 896 -1097
rect 960 -1138 965 -1097
rect 960 -1161 976 -1138
rect 1040 -1161 1182 -1097
rect 1257 -1138 1262 -1097
rect 1246 -1161 1262 -1138
rect 1326 -1161 1342 -1097
rect 1406 -1161 1422 -1097
rect 1486 -1161 1502 -1097
rect 1566 -1161 1582 -1097
rect 1646 -1161 1788 -1097
rect 1852 -1161 1868 -1097
rect 1932 -1161 1948 -1097
rect 2012 -1161 2028 -1097
rect 2092 -1161 2108 -1097
rect 2172 -1138 2177 -1097
rect 2172 -1161 2188 -1138
rect 2252 -1161 2394 -1097
rect 2469 -1138 2474 -1097
rect 2458 -1161 2474 -1138
rect 2538 -1161 2554 -1097
rect 2618 -1161 2634 -1097
rect 2698 -1161 2714 -1097
rect 2778 -1161 2794 -1097
rect 2858 -1161 3000 -1097
rect 3064 -1161 3080 -1097
rect 3144 -1161 3160 -1097
rect 3224 -1161 3240 -1097
rect 3304 -1161 3320 -1097
rect 3384 -1138 3389 -1097
rect 3384 -1161 3400 -1138
rect 3464 -1161 3606 -1097
rect 3681 -1138 3686 -1097
rect 3670 -1161 3686 -1138
rect 3750 -1161 3766 -1097
rect 3830 -1161 3846 -1097
rect 3910 -1161 3926 -1097
rect 3990 -1161 4006 -1097
rect 4070 -1161 4212 -1097
rect 4276 -1161 4292 -1097
rect 4356 -1161 4372 -1097
rect 4436 -1161 4452 -1097
rect 4516 -1161 4532 -1097
rect 4596 -1138 4601 -1097
rect 4596 -1161 4612 -1138
rect 4676 -1161 4818 -1097
rect 4893 -1138 4898 -1097
rect 4882 -1161 4898 -1138
rect 4962 -1161 4978 -1097
rect 5042 -1161 5058 -1097
rect 5122 -1161 5138 -1097
rect 5202 -1161 5218 -1097
rect 5282 -1161 5386 -1097
rect 472 -1163 5386 -1161
rect 472 -1317 538 -1163
rect 284 -1337 410 -1327
rect 284 -1401 315 -1337
rect 379 -1401 410 -1337
rect 284 -1411 410 -1401
rect 472 -1381 473 -1317
rect 537 -1381 538 -1317
rect 472 -1397 538 -1381
rect 472 -1461 473 -1397
rect 537 -1461 538 -1397
rect 472 -1477 538 -1461
rect 472 -1541 473 -1477
rect 537 -1541 538 -1477
rect 472 -1557 538 -1541
rect 472 -1621 473 -1557
rect 537 -1621 538 -1557
rect 472 -1637 538 -1621
rect 472 -1701 473 -1637
rect 537 -1701 538 -1637
rect 472 -1717 538 -1701
rect 472 -1781 473 -1717
rect 537 -1781 538 -1717
rect 472 -1797 538 -1781
rect 472 -1861 473 -1797
rect 537 -1861 538 -1797
rect 472 -1877 538 -1861
rect 472 -1941 473 -1877
rect 537 -1941 538 -1877
rect 472 -1957 538 -1941
rect 472 -2021 473 -1957
rect 537 -2021 538 -1957
rect 472 -2037 538 -2021
rect 472 -2101 473 -2037
rect 537 -2101 538 -2037
rect 472 -2191 538 -2101
rect 598 -2195 658 -1163
rect 718 -2255 778 -1225
rect 838 -2195 898 -1163
rect 958 -2255 1018 -1225
rect 1078 -1317 1144 -1163
rect 1078 -1381 1079 -1317
rect 1143 -1381 1144 -1317
rect 1078 -1397 1144 -1381
rect 1078 -1461 1079 -1397
rect 1143 -1461 1144 -1397
rect 1078 -1477 1144 -1461
rect 1078 -1541 1079 -1477
rect 1143 -1541 1144 -1477
rect 1078 -1557 1144 -1541
rect 1078 -1621 1079 -1557
rect 1143 -1621 1144 -1557
rect 1078 -1637 1144 -1621
rect 1078 -1701 1079 -1637
rect 1143 -1701 1144 -1637
rect 1078 -1717 1144 -1701
rect 1078 -1781 1079 -1717
rect 1143 -1781 1144 -1717
rect 1078 -1797 1144 -1781
rect 1078 -1861 1079 -1797
rect 1143 -1861 1144 -1797
rect 1078 -1877 1144 -1861
rect 1078 -1941 1079 -1877
rect 1143 -1941 1144 -1877
rect 1078 -1957 1144 -1941
rect 1078 -2021 1079 -1957
rect 1143 -2021 1144 -1957
rect 1078 -2037 1144 -2021
rect 1078 -2101 1079 -2037
rect 1143 -2101 1144 -2037
rect 1078 -2191 1144 -2101
rect 1204 -2255 1264 -1225
rect 1324 -2195 1384 -1163
rect 1444 -2255 1504 -1225
rect 1564 -2195 1624 -1163
rect 1684 -1317 1750 -1163
rect 1684 -1381 1685 -1317
rect 1749 -1381 1750 -1317
rect 1684 -1397 1750 -1381
rect 1684 -1461 1685 -1397
rect 1749 -1461 1750 -1397
rect 1684 -1477 1750 -1461
rect 1684 -1541 1685 -1477
rect 1749 -1541 1750 -1477
rect 1684 -1557 1750 -1541
rect 1684 -1621 1685 -1557
rect 1749 -1621 1750 -1557
rect 1684 -1637 1750 -1621
rect 1684 -1701 1685 -1637
rect 1749 -1701 1750 -1637
rect 1684 -1717 1750 -1701
rect 1684 -1781 1685 -1717
rect 1749 -1781 1750 -1717
rect 1684 -1797 1750 -1781
rect 1684 -1861 1685 -1797
rect 1749 -1861 1750 -1797
rect 1684 -1877 1750 -1861
rect 1684 -1941 1685 -1877
rect 1749 -1941 1750 -1877
rect 1684 -1957 1750 -1941
rect 1684 -2021 1685 -1957
rect 1749 -2021 1750 -1957
rect 1684 -2037 1750 -2021
rect 1684 -2101 1685 -2037
rect 1749 -2101 1750 -2037
rect 1684 -2191 1750 -2101
rect 1810 -2195 1870 -1163
rect 1930 -2255 1990 -1225
rect 2050 -2195 2110 -1163
rect 2170 -2255 2230 -1225
rect 2290 -1317 2356 -1163
rect 2290 -1381 2291 -1317
rect 2355 -1381 2356 -1317
rect 2290 -1397 2356 -1381
rect 2290 -1461 2291 -1397
rect 2355 -1461 2356 -1397
rect 2290 -1477 2356 -1461
rect 2290 -1541 2291 -1477
rect 2355 -1541 2356 -1477
rect 2290 -1557 2356 -1541
rect 2290 -1621 2291 -1557
rect 2355 -1621 2356 -1557
rect 2290 -1637 2356 -1621
rect 2290 -1701 2291 -1637
rect 2355 -1701 2356 -1637
rect 2290 -1717 2356 -1701
rect 2290 -1781 2291 -1717
rect 2355 -1781 2356 -1717
rect 2290 -1797 2356 -1781
rect 2290 -1861 2291 -1797
rect 2355 -1861 2356 -1797
rect 2290 -1877 2356 -1861
rect 2290 -1941 2291 -1877
rect 2355 -1941 2356 -1877
rect 2290 -1957 2356 -1941
rect 2290 -2021 2291 -1957
rect 2355 -2021 2356 -1957
rect 2290 -2037 2356 -2021
rect 2290 -2101 2291 -2037
rect 2355 -2101 2356 -2037
rect 2290 -2191 2356 -2101
rect 2416 -2255 2476 -1225
rect 2536 -2195 2596 -1163
rect 2656 -2255 2716 -1225
rect 2776 -2195 2836 -1163
rect 2896 -1317 2962 -1163
rect 2896 -1381 2897 -1317
rect 2961 -1381 2962 -1317
rect 2896 -1397 2962 -1381
rect 2896 -1461 2897 -1397
rect 2961 -1461 2962 -1397
rect 2896 -1477 2962 -1461
rect 2896 -1541 2897 -1477
rect 2961 -1541 2962 -1477
rect 2896 -1557 2962 -1541
rect 2896 -1621 2897 -1557
rect 2961 -1621 2962 -1557
rect 2896 -1637 2962 -1621
rect 2896 -1701 2897 -1637
rect 2961 -1701 2962 -1637
rect 2896 -1717 2962 -1701
rect 2896 -1781 2897 -1717
rect 2961 -1781 2962 -1717
rect 2896 -1797 2962 -1781
rect 2896 -1861 2897 -1797
rect 2961 -1861 2962 -1797
rect 2896 -1877 2962 -1861
rect 2896 -1941 2897 -1877
rect 2961 -1941 2962 -1877
rect 2896 -1957 2962 -1941
rect 2896 -2021 2897 -1957
rect 2961 -2021 2962 -1957
rect 2896 -2037 2962 -2021
rect 2896 -2101 2897 -2037
rect 2961 -2101 2962 -2037
rect 2896 -2191 2962 -2101
rect 3022 -2195 3082 -1163
rect 3142 -2255 3202 -1225
rect 3262 -2195 3322 -1163
rect 3382 -2255 3442 -1225
rect 3502 -1317 3568 -1163
rect 3502 -1381 3503 -1317
rect 3567 -1381 3568 -1317
rect 3502 -1397 3568 -1381
rect 3502 -1461 3503 -1397
rect 3567 -1461 3568 -1397
rect 3502 -1477 3568 -1461
rect 3502 -1541 3503 -1477
rect 3567 -1541 3568 -1477
rect 3502 -1557 3568 -1541
rect 3502 -1621 3503 -1557
rect 3567 -1621 3568 -1557
rect 3502 -1637 3568 -1621
rect 3502 -1701 3503 -1637
rect 3567 -1701 3568 -1637
rect 3502 -1717 3568 -1701
rect 3502 -1781 3503 -1717
rect 3567 -1781 3568 -1717
rect 3502 -1797 3568 -1781
rect 3502 -1861 3503 -1797
rect 3567 -1861 3568 -1797
rect 3502 -1877 3568 -1861
rect 3502 -1941 3503 -1877
rect 3567 -1941 3568 -1877
rect 3502 -1957 3568 -1941
rect 3502 -2021 3503 -1957
rect 3567 -2021 3568 -1957
rect 3502 -2037 3568 -2021
rect 3502 -2101 3503 -2037
rect 3567 -2101 3568 -2037
rect 3502 -2191 3568 -2101
rect 3628 -2255 3688 -1225
rect 3748 -2195 3808 -1163
rect 3868 -2255 3928 -1225
rect 3988 -2195 4048 -1163
rect 4108 -1317 4174 -1163
rect 4108 -1381 4109 -1317
rect 4173 -1381 4174 -1317
rect 4108 -1397 4174 -1381
rect 4108 -1461 4109 -1397
rect 4173 -1461 4174 -1397
rect 4108 -1477 4174 -1461
rect 4108 -1541 4109 -1477
rect 4173 -1541 4174 -1477
rect 4108 -1557 4174 -1541
rect 4108 -1621 4109 -1557
rect 4173 -1621 4174 -1557
rect 4108 -1637 4174 -1621
rect 4108 -1701 4109 -1637
rect 4173 -1701 4174 -1637
rect 4108 -1717 4174 -1701
rect 4108 -1781 4109 -1717
rect 4173 -1781 4174 -1717
rect 4108 -1797 4174 -1781
rect 4108 -1861 4109 -1797
rect 4173 -1861 4174 -1797
rect 4108 -1877 4174 -1861
rect 4108 -1941 4109 -1877
rect 4173 -1941 4174 -1877
rect 4108 -1957 4174 -1941
rect 4108 -2021 4109 -1957
rect 4173 -2021 4174 -1957
rect 4108 -2037 4174 -2021
rect 4108 -2101 4109 -2037
rect 4173 -2101 4174 -2037
rect 4108 -2191 4174 -2101
rect 4234 -2195 4294 -1163
rect 4354 -2255 4414 -1225
rect 4474 -2195 4534 -1163
rect 4594 -2255 4654 -1225
rect 4714 -1317 4780 -1163
rect 4714 -1381 4715 -1317
rect 4779 -1381 4780 -1317
rect 4714 -1397 4780 -1381
rect 4714 -1461 4715 -1397
rect 4779 -1461 4780 -1397
rect 4714 -1477 4780 -1461
rect 4714 -1541 4715 -1477
rect 4779 -1541 4780 -1477
rect 4714 -1557 4780 -1541
rect 4714 -1621 4715 -1557
rect 4779 -1621 4780 -1557
rect 4714 -1637 4780 -1621
rect 4714 -1701 4715 -1637
rect 4779 -1701 4780 -1637
rect 4714 -1717 4780 -1701
rect 4714 -1781 4715 -1717
rect 4779 -1781 4780 -1717
rect 4714 -1797 4780 -1781
rect 4714 -1861 4715 -1797
rect 4779 -1861 4780 -1797
rect 4714 -1877 4780 -1861
rect 4714 -1941 4715 -1877
rect 4779 -1941 4780 -1877
rect 4714 -1957 4780 -1941
rect 4714 -2021 4715 -1957
rect 4779 -2021 4780 -1957
rect 4714 -2037 4780 -2021
rect 4714 -2101 4715 -2037
rect 4779 -2101 4780 -2037
rect 4714 -2191 4780 -2101
rect 4840 -2255 4900 -1225
rect 4960 -2195 5020 -1163
rect 5080 -2255 5140 -1225
rect 5200 -2195 5260 -1163
rect 5320 -1317 5386 -1163
rect 5320 -1381 5321 -1317
rect 5385 -1381 5386 -1317
rect 5320 -1397 5386 -1381
rect 5320 -1461 5321 -1397
rect 5385 -1461 5386 -1397
rect 5320 -1477 5386 -1461
rect 5320 -1541 5321 -1477
rect 5385 -1541 5386 -1477
rect 5320 -1557 5386 -1541
rect 5320 -1621 5321 -1557
rect 5385 -1621 5386 -1557
rect 5320 -1637 5386 -1621
rect 5320 -1701 5321 -1637
rect 5385 -1701 5386 -1637
rect 5320 -1717 5386 -1701
rect 5320 -1781 5321 -1717
rect 5385 -1781 5386 -1717
rect 5320 -1797 5386 -1781
rect 5320 -1861 5321 -1797
rect 5385 -1861 5386 -1797
rect 5320 -1877 5386 -1861
rect 5320 -1941 5321 -1877
rect 5385 -1941 5386 -1877
rect 5320 -1957 5386 -1941
rect 5320 -2021 5321 -1957
rect 5385 -2021 5386 -1957
rect 5320 -2037 5386 -2021
rect 5320 -2101 5321 -2037
rect 5385 -2101 5386 -2037
rect 5320 -2191 5386 -2101
rect 5446 -1097 5561 -1095
rect 5625 -1095 5635 -1074
rect 6951 -1076 7077 -1066
rect 5625 -1097 6118 -1095
rect 5446 -1161 5550 -1097
rect 5625 -1138 5630 -1097
rect 5614 -1161 5630 -1138
rect 5694 -1161 5710 -1097
rect 5774 -1161 5790 -1097
rect 5854 -1161 5870 -1097
rect 5934 -1161 5950 -1097
rect 6014 -1161 6118 -1097
rect 5446 -1163 6118 -1161
rect 5446 -1317 5512 -1163
rect 5446 -1381 5447 -1317
rect 5511 -1381 5512 -1317
rect 5446 -1397 5512 -1381
rect 5446 -1461 5447 -1397
rect 5511 -1461 5512 -1397
rect 5446 -1477 5512 -1461
rect 5446 -1541 5447 -1477
rect 5511 -1541 5512 -1477
rect 5446 -1557 5512 -1541
rect 5446 -1621 5447 -1557
rect 5511 -1621 5512 -1557
rect 5446 -1637 5512 -1621
rect 5446 -1701 5447 -1637
rect 5511 -1701 5512 -1637
rect 5446 -1717 5512 -1701
rect 5446 -1781 5447 -1717
rect 5511 -1781 5512 -1717
rect 5446 -1797 5512 -1781
rect 5446 -1861 5447 -1797
rect 5511 -1861 5512 -1797
rect 5446 -1877 5512 -1861
rect 5446 -1941 5447 -1877
rect 5511 -1941 5512 -1877
rect 5446 -1957 5512 -1941
rect 5446 -2021 5447 -1957
rect 5511 -2021 5512 -1957
rect 5446 -2037 5512 -2021
rect 5446 -2101 5447 -2037
rect 5511 -2101 5512 -2037
rect 5446 -2191 5512 -2101
rect 5572 -2255 5632 -1225
rect 5692 -2195 5752 -1163
rect 5812 -2255 5872 -1225
rect 5932 -2195 5992 -1163
rect 6052 -1317 6118 -1163
rect 6344 -1113 6751 -1096
rect 6344 -1177 6383 -1113
rect 6447 -1177 6526 -1113
rect 6590 -1177 6646 -1113
rect 6710 -1177 6751 -1113
rect 6951 -1140 6982 -1076
rect 7046 -1140 7077 -1076
rect 7710 -1074 7793 -1069
rect 7710 -1095 7720 -1074
rect 6951 -1150 7077 -1140
rect 7227 -1097 7720 -1095
rect 7784 -1095 7793 -1074
rect 7939 -1074 8022 -1069
rect 7939 -1095 7948 -1074
rect 7784 -1097 7948 -1095
rect 8012 -1095 8022 -1074
rect 8922 -1074 9005 -1069
rect 8922 -1095 8932 -1074
rect 8012 -1097 8932 -1095
rect 8996 -1095 9005 -1074
rect 9151 -1074 9234 -1069
rect 9151 -1095 9160 -1074
rect 8996 -1097 9160 -1095
rect 9224 -1095 9234 -1074
rect 10134 -1074 10217 -1069
rect 10134 -1095 10144 -1074
rect 9224 -1097 10144 -1095
rect 10208 -1095 10217 -1074
rect 10363 -1074 10446 -1069
rect 10363 -1095 10372 -1074
rect 10208 -1097 10372 -1095
rect 10436 -1095 10446 -1074
rect 11346 -1074 11429 -1069
rect 11346 -1095 11356 -1074
rect 10436 -1097 11356 -1095
rect 11420 -1095 11429 -1074
rect 11575 -1074 11658 -1069
rect 11575 -1095 11584 -1074
rect 11420 -1097 11584 -1095
rect 11648 -1095 11658 -1074
rect 12307 -1074 12390 -1069
rect 12307 -1095 12316 -1074
rect 11648 -1097 12141 -1095
rect 6344 -1192 6751 -1177
rect 7227 -1161 7331 -1097
rect 7395 -1161 7411 -1097
rect 7475 -1161 7491 -1097
rect 7555 -1161 7571 -1097
rect 7635 -1161 7651 -1097
rect 7715 -1138 7720 -1097
rect 7715 -1161 7731 -1138
rect 7795 -1161 7937 -1097
rect 8012 -1138 8017 -1097
rect 8001 -1161 8017 -1138
rect 8081 -1161 8097 -1097
rect 8161 -1161 8177 -1097
rect 8241 -1161 8257 -1097
rect 8321 -1161 8337 -1097
rect 8401 -1161 8543 -1097
rect 8607 -1161 8623 -1097
rect 8687 -1161 8703 -1097
rect 8767 -1161 8783 -1097
rect 8847 -1161 8863 -1097
rect 8927 -1138 8932 -1097
rect 8927 -1161 8943 -1138
rect 9007 -1161 9149 -1097
rect 9224 -1138 9229 -1097
rect 9213 -1161 9229 -1138
rect 9293 -1161 9309 -1097
rect 9373 -1161 9389 -1097
rect 9453 -1161 9469 -1097
rect 9533 -1161 9549 -1097
rect 9613 -1161 9755 -1097
rect 9819 -1161 9835 -1097
rect 9899 -1161 9915 -1097
rect 9979 -1161 9995 -1097
rect 10059 -1161 10075 -1097
rect 10139 -1138 10144 -1097
rect 10139 -1161 10155 -1138
rect 10219 -1161 10361 -1097
rect 10436 -1138 10441 -1097
rect 10425 -1161 10441 -1138
rect 10505 -1161 10521 -1097
rect 10585 -1161 10601 -1097
rect 10665 -1161 10681 -1097
rect 10745 -1161 10761 -1097
rect 10825 -1161 10967 -1097
rect 11031 -1161 11047 -1097
rect 11111 -1161 11127 -1097
rect 11191 -1161 11207 -1097
rect 11271 -1161 11287 -1097
rect 11351 -1138 11356 -1097
rect 11351 -1161 11367 -1138
rect 11431 -1161 11573 -1097
rect 11648 -1138 11653 -1097
rect 11637 -1161 11653 -1138
rect 11717 -1161 11733 -1097
rect 11797 -1161 11813 -1097
rect 11877 -1161 11893 -1097
rect 11957 -1161 11973 -1097
rect 12037 -1161 12141 -1097
rect 7227 -1163 12141 -1161
rect 6511 -1193 6603 -1192
rect 6052 -1381 6053 -1317
rect 6117 -1381 6118 -1317
rect 7227 -1317 7293 -1163
rect 6052 -1397 6118 -1381
rect 6052 -1461 6053 -1397
rect 6117 -1461 6118 -1397
rect 7039 -1337 7165 -1327
rect 7039 -1401 7070 -1337
rect 7134 -1401 7165 -1337
rect 7039 -1411 7165 -1401
rect 7227 -1381 7228 -1317
rect 7292 -1381 7293 -1317
rect 7227 -1397 7293 -1381
rect 6052 -1477 6118 -1461
rect 6052 -1541 6053 -1477
rect 6117 -1541 6118 -1477
rect 6052 -1557 6118 -1541
rect 6052 -1621 6053 -1557
rect 6117 -1621 6118 -1557
rect 6052 -1637 6118 -1621
rect 6052 -1701 6053 -1637
rect 6117 -1701 6118 -1637
rect 7227 -1461 7228 -1397
rect 7292 -1461 7293 -1397
rect 7227 -1477 7293 -1461
rect 7227 -1541 7228 -1477
rect 7292 -1541 7293 -1477
rect 7227 -1557 7293 -1541
rect 7227 -1621 7228 -1557
rect 7292 -1621 7293 -1557
rect 7227 -1637 7293 -1621
rect 6494 -1642 6638 -1641
rect 6052 -1717 6118 -1701
rect 6052 -1781 6053 -1717
rect 6117 -1781 6118 -1717
rect 6350 -1658 6769 -1642
rect 6350 -1659 6533 -1658
rect 6350 -1723 6389 -1659
rect 6453 -1722 6533 -1659
rect 6597 -1659 6769 -1658
rect 6597 -1722 6664 -1659
rect 6453 -1723 6664 -1722
rect 6728 -1723 6769 -1659
rect 6350 -1737 6769 -1723
rect 6350 -1738 6494 -1737
rect 6625 -1738 6769 -1737
rect 7227 -1701 7228 -1637
rect 7292 -1701 7293 -1637
rect 7227 -1717 7293 -1701
rect 6052 -1797 6118 -1781
rect 6052 -1861 6053 -1797
rect 6117 -1861 6118 -1797
rect 6052 -1877 6118 -1861
rect 6052 -1941 6053 -1877
rect 6117 -1941 6118 -1877
rect 6052 -1957 6118 -1941
rect 6052 -2021 6053 -1957
rect 6117 -2021 6118 -1957
rect 6052 -2037 6118 -2021
rect 6052 -2101 6053 -2037
rect 6117 -2101 6118 -2037
rect 6052 -2191 6118 -2101
rect 7227 -1781 7228 -1717
rect 7292 -1781 7293 -1717
rect 7227 -1797 7293 -1781
rect 7227 -1861 7228 -1797
rect 7292 -1861 7293 -1797
rect 7227 -1877 7293 -1861
rect 7227 -1941 7228 -1877
rect 7292 -1941 7293 -1877
rect 7227 -1957 7293 -1941
rect 7227 -2021 7228 -1957
rect 7292 -2021 7293 -1957
rect 7227 -2037 7293 -2021
rect 7227 -2101 7228 -2037
rect 7292 -2101 7293 -2037
rect 7227 -2191 7293 -2101
rect 7353 -2195 7413 -1163
rect 7473 -2255 7533 -1225
rect 7593 -2195 7653 -1163
rect 7713 -2255 7773 -1225
rect 7833 -1317 7899 -1163
rect 7833 -1381 7834 -1317
rect 7898 -1381 7899 -1317
rect 7833 -1397 7899 -1381
rect 7833 -1461 7834 -1397
rect 7898 -1461 7899 -1397
rect 7833 -1477 7899 -1461
rect 7833 -1541 7834 -1477
rect 7898 -1541 7899 -1477
rect 7833 -1557 7899 -1541
rect 7833 -1621 7834 -1557
rect 7898 -1621 7899 -1557
rect 7833 -1637 7899 -1621
rect 7833 -1701 7834 -1637
rect 7898 -1701 7899 -1637
rect 7833 -1717 7899 -1701
rect 7833 -1781 7834 -1717
rect 7898 -1781 7899 -1717
rect 7833 -1797 7899 -1781
rect 7833 -1861 7834 -1797
rect 7898 -1861 7899 -1797
rect 7833 -1877 7899 -1861
rect 7833 -1941 7834 -1877
rect 7898 -1941 7899 -1877
rect 7833 -1957 7899 -1941
rect 7833 -2021 7834 -1957
rect 7898 -2021 7899 -1957
rect 7833 -2037 7899 -2021
rect 7833 -2101 7834 -2037
rect 7898 -2101 7899 -2037
rect 7833 -2191 7899 -2101
rect 7959 -2255 8019 -1225
rect 8079 -2195 8139 -1163
rect 8199 -2255 8259 -1225
rect 8319 -2195 8379 -1163
rect 8439 -1317 8505 -1163
rect 8439 -1381 8440 -1317
rect 8504 -1381 8505 -1317
rect 8439 -1397 8505 -1381
rect 8439 -1461 8440 -1397
rect 8504 -1461 8505 -1397
rect 8439 -1477 8505 -1461
rect 8439 -1541 8440 -1477
rect 8504 -1541 8505 -1477
rect 8439 -1557 8505 -1541
rect 8439 -1621 8440 -1557
rect 8504 -1621 8505 -1557
rect 8439 -1637 8505 -1621
rect 8439 -1701 8440 -1637
rect 8504 -1701 8505 -1637
rect 8439 -1717 8505 -1701
rect 8439 -1781 8440 -1717
rect 8504 -1781 8505 -1717
rect 8439 -1797 8505 -1781
rect 8439 -1861 8440 -1797
rect 8504 -1861 8505 -1797
rect 8439 -1877 8505 -1861
rect 8439 -1941 8440 -1877
rect 8504 -1941 8505 -1877
rect 8439 -1957 8505 -1941
rect 8439 -2021 8440 -1957
rect 8504 -2021 8505 -1957
rect 8439 -2037 8505 -2021
rect 8439 -2101 8440 -2037
rect 8504 -2101 8505 -2037
rect 8439 -2191 8505 -2101
rect 8565 -2195 8625 -1163
rect 8685 -2255 8745 -1225
rect 8805 -2195 8865 -1163
rect 8925 -2255 8985 -1225
rect 9045 -1317 9111 -1163
rect 9045 -1381 9046 -1317
rect 9110 -1381 9111 -1317
rect 9045 -1397 9111 -1381
rect 9045 -1461 9046 -1397
rect 9110 -1461 9111 -1397
rect 9045 -1477 9111 -1461
rect 9045 -1541 9046 -1477
rect 9110 -1541 9111 -1477
rect 9045 -1557 9111 -1541
rect 9045 -1621 9046 -1557
rect 9110 -1621 9111 -1557
rect 9045 -1637 9111 -1621
rect 9045 -1701 9046 -1637
rect 9110 -1701 9111 -1637
rect 9045 -1717 9111 -1701
rect 9045 -1781 9046 -1717
rect 9110 -1781 9111 -1717
rect 9045 -1797 9111 -1781
rect 9045 -1861 9046 -1797
rect 9110 -1861 9111 -1797
rect 9045 -1877 9111 -1861
rect 9045 -1941 9046 -1877
rect 9110 -1941 9111 -1877
rect 9045 -1957 9111 -1941
rect 9045 -2021 9046 -1957
rect 9110 -2021 9111 -1957
rect 9045 -2037 9111 -2021
rect 9045 -2101 9046 -2037
rect 9110 -2101 9111 -2037
rect 9045 -2191 9111 -2101
rect 9171 -2255 9231 -1225
rect 9291 -2195 9351 -1163
rect 9411 -2255 9471 -1225
rect 9531 -2195 9591 -1163
rect 9651 -1317 9717 -1163
rect 9651 -1381 9652 -1317
rect 9716 -1381 9717 -1317
rect 9651 -1397 9717 -1381
rect 9651 -1461 9652 -1397
rect 9716 -1461 9717 -1397
rect 9651 -1477 9717 -1461
rect 9651 -1541 9652 -1477
rect 9716 -1541 9717 -1477
rect 9651 -1557 9717 -1541
rect 9651 -1621 9652 -1557
rect 9716 -1621 9717 -1557
rect 9651 -1637 9717 -1621
rect 9651 -1701 9652 -1637
rect 9716 -1701 9717 -1637
rect 9651 -1717 9717 -1701
rect 9651 -1781 9652 -1717
rect 9716 -1781 9717 -1717
rect 9651 -1797 9717 -1781
rect 9651 -1861 9652 -1797
rect 9716 -1861 9717 -1797
rect 9651 -1877 9717 -1861
rect 9651 -1941 9652 -1877
rect 9716 -1941 9717 -1877
rect 9651 -1957 9717 -1941
rect 9651 -2021 9652 -1957
rect 9716 -2021 9717 -1957
rect 9651 -2037 9717 -2021
rect 9651 -2101 9652 -2037
rect 9716 -2101 9717 -2037
rect 9651 -2191 9717 -2101
rect 9777 -2195 9837 -1163
rect 9897 -2255 9957 -1225
rect 10017 -2195 10077 -1163
rect 10137 -2255 10197 -1225
rect 10257 -1317 10323 -1163
rect 10257 -1381 10258 -1317
rect 10322 -1381 10323 -1317
rect 10257 -1397 10323 -1381
rect 10257 -1461 10258 -1397
rect 10322 -1461 10323 -1397
rect 10257 -1477 10323 -1461
rect 10257 -1541 10258 -1477
rect 10322 -1541 10323 -1477
rect 10257 -1557 10323 -1541
rect 10257 -1621 10258 -1557
rect 10322 -1621 10323 -1557
rect 10257 -1637 10323 -1621
rect 10257 -1701 10258 -1637
rect 10322 -1701 10323 -1637
rect 10257 -1717 10323 -1701
rect 10257 -1781 10258 -1717
rect 10322 -1781 10323 -1717
rect 10257 -1797 10323 -1781
rect 10257 -1861 10258 -1797
rect 10322 -1861 10323 -1797
rect 10257 -1877 10323 -1861
rect 10257 -1941 10258 -1877
rect 10322 -1941 10323 -1877
rect 10257 -1957 10323 -1941
rect 10257 -2021 10258 -1957
rect 10322 -2021 10323 -1957
rect 10257 -2037 10323 -2021
rect 10257 -2101 10258 -2037
rect 10322 -2101 10323 -2037
rect 10257 -2191 10323 -2101
rect 10383 -2255 10443 -1225
rect 10503 -2195 10563 -1163
rect 10623 -2255 10683 -1225
rect 10743 -2195 10803 -1163
rect 10863 -1317 10929 -1163
rect 10863 -1381 10864 -1317
rect 10928 -1381 10929 -1317
rect 10863 -1397 10929 -1381
rect 10863 -1461 10864 -1397
rect 10928 -1461 10929 -1397
rect 10863 -1477 10929 -1461
rect 10863 -1541 10864 -1477
rect 10928 -1541 10929 -1477
rect 10863 -1557 10929 -1541
rect 10863 -1621 10864 -1557
rect 10928 -1621 10929 -1557
rect 10863 -1637 10929 -1621
rect 10863 -1701 10864 -1637
rect 10928 -1701 10929 -1637
rect 10863 -1717 10929 -1701
rect 10863 -1781 10864 -1717
rect 10928 -1781 10929 -1717
rect 10863 -1797 10929 -1781
rect 10863 -1861 10864 -1797
rect 10928 -1861 10929 -1797
rect 10863 -1877 10929 -1861
rect 10863 -1941 10864 -1877
rect 10928 -1941 10929 -1877
rect 10863 -1957 10929 -1941
rect 10863 -2021 10864 -1957
rect 10928 -2021 10929 -1957
rect 10863 -2037 10929 -2021
rect 10863 -2101 10864 -2037
rect 10928 -2101 10929 -2037
rect 10863 -2191 10929 -2101
rect 10989 -2195 11049 -1163
rect 11109 -2255 11169 -1225
rect 11229 -2195 11289 -1163
rect 11349 -2255 11409 -1225
rect 11469 -1317 11535 -1163
rect 11469 -1381 11470 -1317
rect 11534 -1381 11535 -1317
rect 11469 -1397 11535 -1381
rect 11469 -1461 11470 -1397
rect 11534 -1461 11535 -1397
rect 11469 -1477 11535 -1461
rect 11469 -1541 11470 -1477
rect 11534 -1541 11535 -1477
rect 11469 -1557 11535 -1541
rect 11469 -1621 11470 -1557
rect 11534 -1621 11535 -1557
rect 11469 -1637 11535 -1621
rect 11469 -1701 11470 -1637
rect 11534 -1701 11535 -1637
rect 11469 -1717 11535 -1701
rect 11469 -1781 11470 -1717
rect 11534 -1781 11535 -1717
rect 11469 -1797 11535 -1781
rect 11469 -1861 11470 -1797
rect 11534 -1861 11535 -1797
rect 11469 -1877 11535 -1861
rect 11469 -1941 11470 -1877
rect 11534 -1941 11535 -1877
rect 11469 -1957 11535 -1941
rect 11469 -2021 11470 -1957
rect 11534 -2021 11535 -1957
rect 11469 -2037 11535 -2021
rect 11469 -2101 11470 -2037
rect 11534 -2101 11535 -2037
rect 11469 -2191 11535 -2101
rect 11595 -2255 11655 -1225
rect 11715 -2195 11775 -1163
rect 11835 -2255 11895 -1225
rect 11955 -2195 12015 -1163
rect 12075 -1317 12141 -1163
rect 12075 -1381 12076 -1317
rect 12140 -1381 12141 -1317
rect 12075 -1397 12141 -1381
rect 12075 -1461 12076 -1397
rect 12140 -1461 12141 -1397
rect 12075 -1477 12141 -1461
rect 12075 -1541 12076 -1477
rect 12140 -1541 12141 -1477
rect 12075 -1557 12141 -1541
rect 12075 -1621 12076 -1557
rect 12140 -1621 12141 -1557
rect 12075 -1637 12141 -1621
rect 12075 -1701 12076 -1637
rect 12140 -1701 12141 -1637
rect 12075 -1717 12141 -1701
rect 12075 -1781 12076 -1717
rect 12140 -1781 12141 -1717
rect 12075 -1797 12141 -1781
rect 12075 -1861 12076 -1797
rect 12140 -1861 12141 -1797
rect 12075 -1877 12141 -1861
rect 12075 -1941 12076 -1877
rect 12140 -1941 12141 -1877
rect 12075 -1957 12141 -1941
rect 12075 -2021 12076 -1957
rect 12140 -2021 12141 -1957
rect 12075 -2037 12141 -2021
rect 12075 -2101 12076 -2037
rect 12140 -2101 12141 -2037
rect 12075 -2191 12141 -2101
rect 12201 -1097 12316 -1095
rect 12380 -1095 12390 -1074
rect 12380 -1097 12873 -1095
rect 12201 -1161 12305 -1097
rect 12380 -1138 12385 -1097
rect 12369 -1161 12385 -1138
rect 12449 -1161 12465 -1097
rect 12529 -1161 12545 -1097
rect 12609 -1161 12625 -1097
rect 12689 -1161 12705 -1097
rect 12769 -1161 12873 -1097
rect 12201 -1163 12873 -1161
rect 12201 -1317 12267 -1163
rect 12201 -1381 12202 -1317
rect 12266 -1381 12267 -1317
rect 12201 -1397 12267 -1381
rect 12201 -1461 12202 -1397
rect 12266 -1461 12267 -1397
rect 12201 -1477 12267 -1461
rect 12201 -1541 12202 -1477
rect 12266 -1541 12267 -1477
rect 12201 -1557 12267 -1541
rect 12201 -1621 12202 -1557
rect 12266 -1621 12267 -1557
rect 12201 -1637 12267 -1621
rect 12201 -1701 12202 -1637
rect 12266 -1701 12267 -1637
rect 12201 -1717 12267 -1701
rect 12201 -1781 12202 -1717
rect 12266 -1781 12267 -1717
rect 12201 -1797 12267 -1781
rect 12201 -1861 12202 -1797
rect 12266 -1861 12267 -1797
rect 12201 -1877 12267 -1861
rect 12201 -1941 12202 -1877
rect 12266 -1941 12267 -1877
rect 12201 -1957 12267 -1941
rect 12201 -2021 12202 -1957
rect 12266 -2021 12267 -1957
rect 12201 -2037 12267 -2021
rect 12201 -2101 12202 -2037
rect 12266 -2101 12267 -2037
rect 12201 -2191 12267 -2101
rect 12327 -2255 12387 -1225
rect 12447 -2195 12507 -1163
rect 12567 -2255 12627 -1225
rect 12687 -2195 12747 -1163
rect 12807 -1317 12873 -1163
rect 13099 -1113 13506 -1096
rect 13099 -1177 13138 -1113
rect 13202 -1177 13281 -1113
rect 13345 -1177 13401 -1113
rect 13465 -1177 13506 -1113
rect 13099 -1192 13506 -1177
rect 13266 -1193 13358 -1192
rect 12807 -1381 12808 -1317
rect 12872 -1381 12873 -1317
rect 12807 -1397 12873 -1381
rect 12807 -1461 12808 -1397
rect 12872 -1461 12873 -1397
rect 12807 -1477 12873 -1461
rect 12807 -1541 12808 -1477
rect 12872 -1541 12873 -1477
rect 12807 -1557 12873 -1541
rect 12807 -1621 12808 -1557
rect 12872 -1621 12873 -1557
rect 12807 -1637 12873 -1621
rect 12807 -1701 12808 -1637
rect 12872 -1701 12873 -1637
rect 13249 -1642 13393 -1641
rect 12807 -1717 12873 -1701
rect 12807 -1781 12808 -1717
rect 12872 -1781 12873 -1717
rect 13105 -1658 13524 -1642
rect 13105 -1659 13288 -1658
rect 13105 -1723 13144 -1659
rect 13208 -1722 13288 -1659
rect 13352 -1659 13524 -1658
rect 13352 -1722 13419 -1659
rect 13208 -1723 13419 -1722
rect 13483 -1723 13524 -1659
rect 13105 -1737 13524 -1723
rect 13105 -1738 13249 -1737
rect 13380 -1738 13524 -1737
rect 12807 -1797 12873 -1781
rect 12807 -1861 12808 -1797
rect 12872 -1861 12873 -1797
rect 12807 -1877 12873 -1861
rect 12807 -1941 12808 -1877
rect 12872 -1941 12873 -1877
rect 12807 -1957 12873 -1941
rect 12807 -2021 12808 -1957
rect 12872 -2021 12873 -1957
rect 12807 -2037 12873 -2021
rect 12807 -2101 12808 -2037
rect 12872 -2101 12873 -2037
rect 12807 -2191 12873 -2101
rect 472 -2257 5386 -2255
rect 472 -2321 576 -2257
rect 640 -2321 656 -2257
rect 720 -2321 736 -2257
rect 800 -2321 816 -2257
rect 880 -2321 896 -2257
rect 960 -2321 976 -2257
rect 1040 -2321 1182 -2257
rect 1246 -2321 1262 -2257
rect 1326 -2321 1342 -2257
rect 1406 -2321 1422 -2257
rect 1486 -2321 1502 -2257
rect 1566 -2321 1582 -2257
rect 1646 -2321 1788 -2257
rect 1852 -2321 1868 -2257
rect 1932 -2321 1948 -2257
rect 2012 -2321 2028 -2257
rect 2092 -2321 2108 -2257
rect 2172 -2321 2188 -2257
rect 2252 -2321 2394 -2257
rect 2458 -2321 2474 -2257
rect 2538 -2321 2554 -2257
rect 2618 -2321 2634 -2257
rect 2698 -2321 2714 -2257
rect 2778 -2321 2794 -2257
rect 2858 -2321 3000 -2257
rect 3064 -2321 3080 -2257
rect 3144 -2321 3160 -2257
rect 3224 -2321 3240 -2257
rect 3304 -2321 3320 -2257
rect 3384 -2321 3400 -2257
rect 3464 -2321 3606 -2257
rect 3670 -2321 3686 -2257
rect 3750 -2321 3766 -2257
rect 3830 -2321 3846 -2257
rect 3910 -2321 3926 -2257
rect 3990 -2321 4006 -2257
rect 4070 -2321 4212 -2257
rect 4276 -2321 4292 -2257
rect 4356 -2321 4372 -2257
rect 4436 -2321 4452 -2257
rect 4516 -2321 4532 -2257
rect 4596 -2321 4612 -2257
rect 4676 -2321 4818 -2257
rect 4882 -2321 4898 -2257
rect 4962 -2321 4978 -2257
rect 5042 -2321 5058 -2257
rect 5122 -2321 5138 -2257
rect 5202 -2321 5218 -2257
rect 5282 -2321 5386 -2257
rect 472 -2323 5386 -2321
rect 5446 -2257 6142 -2255
rect 5446 -2321 5550 -2257
rect 5614 -2321 5630 -2257
rect 5694 -2321 5710 -2257
rect 5774 -2321 5790 -2257
rect 5854 -2321 5870 -2257
rect 5934 -2321 5950 -2257
rect 6014 -2264 6142 -2257
rect 6014 -2321 6047 -2264
rect 5446 -2323 6047 -2321
rect 6016 -2328 6047 -2323
rect 6111 -2328 6142 -2264
rect 7227 -2257 12141 -2255
rect 7227 -2321 7331 -2257
rect 7395 -2321 7411 -2257
rect 7475 -2321 7491 -2257
rect 7555 -2321 7571 -2257
rect 7635 -2321 7651 -2257
rect 7715 -2321 7731 -2257
rect 7795 -2321 7937 -2257
rect 8001 -2321 8017 -2257
rect 8081 -2321 8097 -2257
rect 8161 -2321 8177 -2257
rect 8241 -2321 8257 -2257
rect 8321 -2321 8337 -2257
rect 8401 -2321 8543 -2257
rect 8607 -2321 8623 -2257
rect 8687 -2321 8703 -2257
rect 8767 -2321 8783 -2257
rect 8847 -2321 8863 -2257
rect 8927 -2321 8943 -2257
rect 9007 -2321 9149 -2257
rect 9213 -2321 9229 -2257
rect 9293 -2321 9309 -2257
rect 9373 -2321 9389 -2257
rect 9453 -2321 9469 -2257
rect 9533 -2321 9549 -2257
rect 9613 -2321 9755 -2257
rect 9819 -2321 9835 -2257
rect 9899 -2321 9915 -2257
rect 9979 -2321 9995 -2257
rect 10059 -2321 10075 -2257
rect 10139 -2321 10155 -2257
rect 10219 -2321 10361 -2257
rect 10425 -2321 10441 -2257
rect 10505 -2321 10521 -2257
rect 10585 -2321 10601 -2257
rect 10665 -2321 10681 -2257
rect 10745 -2321 10761 -2257
rect 10825 -2321 10967 -2257
rect 11031 -2321 11047 -2257
rect 11111 -2321 11127 -2257
rect 11191 -2321 11207 -2257
rect 11271 -2321 11287 -2257
rect 11351 -2321 11367 -2257
rect 11431 -2321 11573 -2257
rect 11637 -2321 11653 -2257
rect 11717 -2321 11733 -2257
rect 11797 -2321 11813 -2257
rect 11877 -2321 11893 -2257
rect 11957 -2321 11973 -2257
rect 12037 -2321 12141 -2257
rect 7227 -2323 12141 -2321
rect 12201 -2257 12897 -2255
rect 12201 -2321 12305 -2257
rect 12369 -2321 12385 -2257
rect 12449 -2321 12465 -2257
rect 12529 -2321 12545 -2257
rect 12609 -2321 12625 -2257
rect 12689 -2321 12705 -2257
rect 12769 -2264 12897 -2257
rect 12769 -2321 12802 -2264
rect 12201 -2323 12802 -2321
rect 6016 -2338 6142 -2328
rect 12771 -2328 12802 -2323
rect 12866 -2328 12897 -2264
rect 12771 -2338 12897 -2328
<< via3 >>
rect 738 3272 802 3276
rect 738 3216 742 3272
rect 742 3216 798 3272
rect 798 3216 802 3272
rect 738 3212 802 3216
rect 835 3205 899 3269
rect 915 3205 979 3269
rect 995 3205 1059 3269
rect 1075 3205 1139 3269
rect 1155 3205 1219 3269
rect 1235 3205 1299 3269
rect 1567 3205 1631 3269
rect 1647 3205 1711 3269
rect 1727 3205 1791 3269
rect 1807 3205 1871 3269
rect 1887 3205 1951 3269
rect 1967 3205 2031 3269
rect 2173 3205 2237 3269
rect 2253 3205 2317 3269
rect 2333 3205 2397 3269
rect 2413 3205 2477 3269
rect 2493 3205 2557 3269
rect 2573 3205 2637 3269
rect 2779 3205 2843 3269
rect 2859 3205 2923 3269
rect 2939 3205 3003 3269
rect 3019 3205 3083 3269
rect 3099 3205 3163 3269
rect 3179 3205 3243 3269
rect 3385 3205 3449 3269
rect 3465 3205 3529 3269
rect 3545 3205 3609 3269
rect 3625 3205 3689 3269
rect 3705 3205 3769 3269
rect 3785 3205 3849 3269
rect 3991 3205 4055 3269
rect 4071 3205 4135 3269
rect 4151 3205 4215 3269
rect 4231 3205 4295 3269
rect 4311 3205 4375 3269
rect 4391 3205 4455 3269
rect 4597 3205 4661 3269
rect 4677 3205 4741 3269
rect 4757 3205 4821 3269
rect 4837 3205 4901 3269
rect 4917 3205 4981 3269
rect 4997 3205 5061 3269
rect 5203 3205 5267 3269
rect 5283 3205 5347 3269
rect 5363 3205 5427 3269
rect 5443 3205 5507 3269
rect 5523 3205 5587 3269
rect 5603 3205 5667 3269
rect 5809 3205 5873 3269
rect 5889 3205 5953 3269
rect 5969 3205 6033 3269
rect 6049 3205 6113 3269
rect 6129 3205 6193 3269
rect 6209 3205 6273 3269
rect 7427 3272 7491 3276
rect 7427 3216 7431 3272
rect 7431 3216 7487 3272
rect 7487 3216 7491 3272
rect 7427 3212 7491 3216
rect 7524 3205 7588 3269
rect 7604 3205 7668 3269
rect 7684 3205 7748 3269
rect 7764 3205 7828 3269
rect 7844 3205 7908 3269
rect 7924 3205 7988 3269
rect 8256 3205 8320 3269
rect 8336 3205 8400 3269
rect 8416 3205 8480 3269
rect 8496 3205 8560 3269
rect 8576 3205 8640 3269
rect 8656 3205 8720 3269
rect 8862 3205 8926 3269
rect 8942 3205 9006 3269
rect 9022 3205 9086 3269
rect 9102 3205 9166 3269
rect 9182 3205 9246 3269
rect 9262 3205 9326 3269
rect 9468 3205 9532 3269
rect 9548 3205 9612 3269
rect 9628 3205 9692 3269
rect 9708 3205 9772 3269
rect 9788 3205 9852 3269
rect 9868 3205 9932 3269
rect 10074 3205 10138 3269
rect 10154 3205 10218 3269
rect 10234 3205 10298 3269
rect 10314 3205 10378 3269
rect 10394 3205 10458 3269
rect 10474 3205 10538 3269
rect 10680 3205 10744 3269
rect 10760 3205 10824 3269
rect 10840 3205 10904 3269
rect 10920 3205 10984 3269
rect 11000 3205 11064 3269
rect 11080 3205 11144 3269
rect 11286 3205 11350 3269
rect 11366 3205 11430 3269
rect 11446 3205 11510 3269
rect 11526 3205 11590 3269
rect 11606 3205 11670 3269
rect 11686 3205 11750 3269
rect 11892 3205 11956 3269
rect 11972 3205 12036 3269
rect 12052 3205 12116 3269
rect 12132 3205 12196 3269
rect 12212 3205 12276 3269
rect 12292 3205 12356 3269
rect 12498 3205 12562 3269
rect 12578 3205 12642 3269
rect 12658 3205 12722 3269
rect 12738 3205 12802 3269
rect 12818 3205 12882 3269
rect 12898 3205 12962 3269
rect 732 2985 796 3049
rect 732 2905 796 2969
rect 732 2825 796 2889
rect 732 2745 796 2809
rect 121 2667 185 2671
rect 121 2611 125 2667
rect 125 2611 181 2667
rect 181 2611 185 2667
rect 121 2607 185 2611
rect 252 2666 316 2670
rect 252 2610 256 2666
rect 256 2610 312 2666
rect 312 2610 316 2666
rect 252 2606 316 2610
rect 396 2667 460 2671
rect 396 2611 400 2667
rect 400 2611 456 2667
rect 456 2611 460 2667
rect 396 2607 460 2611
rect 732 2665 796 2729
rect 732 2585 796 2649
rect 732 2505 796 2569
rect 732 2425 796 2489
rect 732 2345 796 2409
rect 732 2265 796 2329
rect 139 2121 203 2125
rect 139 2065 143 2121
rect 143 2065 199 2121
rect 199 2065 203 2121
rect 139 2061 203 2065
rect 259 2121 323 2125
rect 259 2065 263 2121
rect 263 2065 319 2121
rect 319 2065 323 2121
rect 259 2061 323 2065
rect 402 2121 466 2125
rect 402 2065 406 2121
rect 406 2065 462 2121
rect 462 2065 466 2121
rect 402 2061 466 2065
rect 1338 2985 1402 3049
rect 1338 2905 1402 2969
rect 1338 2825 1402 2889
rect 1338 2745 1402 2809
rect 1338 2665 1402 2729
rect 1338 2585 1402 2649
rect 1338 2505 1402 2569
rect 1338 2425 1402 2489
rect 1338 2345 1402 2409
rect 1338 2265 1402 2329
rect 835 2045 899 2109
rect 915 2045 979 2109
rect 995 2045 1059 2109
rect 1075 2045 1139 2109
rect 1155 2045 1219 2109
rect 1235 2086 1299 2109
rect 1235 2045 1288 2086
rect 1288 2045 1299 2086
rect 1464 2985 1528 3049
rect 1464 2905 1528 2969
rect 1464 2825 1528 2889
rect 1464 2745 1528 2809
rect 1464 2665 1528 2729
rect 1464 2585 1528 2649
rect 1464 2505 1528 2569
rect 1464 2425 1528 2489
rect 1464 2345 1528 2409
rect 1464 2265 1528 2329
rect 2070 2985 2134 3049
rect 2070 2905 2134 2969
rect 2070 2825 2134 2889
rect 2070 2745 2134 2809
rect 2070 2665 2134 2729
rect 2070 2585 2134 2649
rect 2070 2505 2134 2569
rect 2070 2425 2134 2489
rect 2070 2345 2134 2409
rect 2070 2265 2134 2329
rect 2676 2985 2740 3049
rect 2676 2905 2740 2969
rect 2676 2825 2740 2889
rect 2676 2745 2740 2809
rect 2676 2665 2740 2729
rect 2676 2585 2740 2649
rect 2676 2505 2740 2569
rect 2676 2425 2740 2489
rect 2676 2345 2740 2409
rect 2676 2265 2740 2329
rect 3282 2985 3346 3049
rect 3282 2905 3346 2969
rect 3282 2825 3346 2889
rect 3282 2745 3346 2809
rect 3282 2665 3346 2729
rect 3282 2585 3346 2649
rect 3282 2505 3346 2569
rect 3282 2425 3346 2489
rect 3282 2345 3346 2409
rect 3282 2265 3346 2329
rect 3888 2985 3952 3049
rect 3888 2905 3952 2969
rect 3888 2825 3952 2889
rect 3888 2745 3952 2809
rect 3888 2665 3952 2729
rect 3888 2585 3952 2649
rect 3888 2505 3952 2569
rect 3888 2425 3952 2489
rect 3888 2345 3952 2409
rect 3888 2265 3952 2329
rect 4494 2985 4558 3049
rect 4494 2905 4558 2969
rect 4494 2825 4558 2889
rect 4494 2745 4558 2809
rect 4494 2665 4558 2729
rect 4494 2585 4558 2649
rect 4494 2505 4558 2569
rect 4494 2425 4558 2489
rect 4494 2345 4558 2409
rect 4494 2265 4558 2329
rect 5100 2985 5164 3049
rect 5100 2905 5164 2969
rect 5100 2825 5164 2889
rect 5100 2745 5164 2809
rect 5100 2665 5164 2729
rect 5100 2585 5164 2649
rect 5100 2505 5164 2569
rect 5100 2425 5164 2489
rect 5100 2345 5164 2409
rect 5100 2265 5164 2329
rect 5706 2985 5770 3049
rect 5706 2905 5770 2969
rect 5706 2825 5770 2889
rect 5706 2745 5770 2809
rect 5706 2665 5770 2729
rect 5706 2585 5770 2649
rect 5706 2505 5770 2569
rect 5706 2425 5770 2489
rect 5706 2345 5770 2409
rect 5706 2265 5770 2329
rect 6312 2985 6376 3049
rect 6312 2905 6376 2969
rect 6312 2825 6376 2889
rect 6312 2745 6376 2809
rect 6312 2665 6376 2729
rect 7421 2985 7485 3049
rect 7421 2905 7485 2969
rect 7421 2825 7485 2889
rect 7421 2745 7485 2809
rect 6312 2585 6376 2649
rect 6810 2667 6874 2671
rect 6810 2611 6814 2667
rect 6814 2611 6870 2667
rect 6870 2611 6874 2667
rect 6810 2607 6874 2611
rect 6941 2666 7005 2670
rect 6941 2610 6945 2666
rect 6945 2610 7001 2666
rect 7001 2610 7005 2666
rect 6941 2606 7005 2610
rect 7085 2667 7149 2671
rect 7085 2611 7089 2667
rect 7089 2611 7145 2667
rect 7145 2611 7149 2667
rect 7085 2607 7149 2611
rect 7421 2665 7485 2729
rect 6312 2505 6376 2569
rect 6312 2425 6376 2489
rect 6312 2345 6376 2409
rect 7421 2585 7485 2649
rect 7421 2505 7485 2569
rect 7421 2425 7485 2489
rect 6312 2265 6376 2329
rect 6470 2345 6534 2349
rect 6470 2289 6474 2345
rect 6474 2289 6530 2345
rect 6530 2289 6534 2345
rect 6470 2285 6534 2289
rect 7421 2345 7485 2409
rect 7421 2265 7485 2329
rect 1567 2045 1631 2109
rect 1647 2045 1711 2109
rect 1727 2045 1791 2109
rect 1807 2045 1871 2109
rect 1887 2045 1951 2109
rect 1967 2086 2031 2109
rect 1967 2045 2020 2086
rect 2020 2045 2031 2086
rect 2173 2086 2237 2109
rect 2173 2045 2184 2086
rect 2184 2045 2237 2086
rect 2253 2045 2317 2109
rect 2333 2045 2397 2109
rect 2413 2045 2477 2109
rect 2493 2045 2557 2109
rect 2573 2045 2637 2109
rect 2779 2045 2843 2109
rect 2859 2045 2923 2109
rect 2939 2045 3003 2109
rect 3019 2045 3083 2109
rect 3099 2045 3163 2109
rect 3179 2086 3243 2109
rect 3179 2045 3232 2086
rect 3232 2045 3243 2086
rect 3385 2086 3449 2109
rect 3385 2045 3396 2086
rect 3396 2045 3449 2086
rect 3465 2045 3529 2109
rect 3545 2045 3609 2109
rect 3625 2045 3689 2109
rect 3705 2045 3769 2109
rect 3785 2045 3849 2109
rect 3991 2045 4055 2109
rect 4071 2045 4135 2109
rect 4151 2045 4215 2109
rect 4231 2045 4295 2109
rect 4311 2045 4375 2109
rect 4391 2086 4455 2109
rect 4391 2045 4444 2086
rect 4444 2045 4455 2086
rect 4597 2086 4661 2109
rect 4597 2045 4608 2086
rect 4608 2045 4661 2086
rect 4677 2045 4741 2109
rect 4757 2045 4821 2109
rect 4837 2045 4901 2109
rect 4917 2045 4981 2109
rect 4997 2045 5061 2109
rect 5203 2045 5267 2109
rect 5283 2045 5347 2109
rect 5363 2045 5427 2109
rect 5443 2045 5507 2109
rect 5523 2045 5587 2109
rect 5603 2086 5667 2109
rect 5603 2045 5656 2086
rect 5656 2045 5667 2086
rect 5809 2086 5873 2109
rect 5809 2045 5820 2086
rect 5820 2045 5873 2086
rect 5889 2045 5953 2109
rect 5969 2045 6033 2109
rect 6049 2045 6113 2109
rect 6129 2045 6193 2109
rect 6209 2045 6273 2109
rect 6558 2084 6622 2088
rect 6558 2028 6562 2084
rect 6562 2028 6618 2084
rect 6618 2028 6622 2084
rect 6558 2024 6622 2028
rect 6828 2121 6892 2125
rect 6828 2065 6832 2121
rect 6832 2065 6888 2121
rect 6888 2065 6892 2121
rect 6828 2061 6892 2065
rect 6948 2121 7012 2125
rect 6948 2065 6952 2121
rect 6952 2065 7008 2121
rect 7008 2065 7012 2121
rect 6948 2061 7012 2065
rect 7091 2121 7155 2125
rect 7091 2065 7095 2121
rect 7095 2065 7151 2121
rect 7151 2065 7155 2121
rect 7091 2061 7155 2065
rect 8027 2985 8091 3049
rect 8027 2905 8091 2969
rect 8027 2825 8091 2889
rect 8027 2745 8091 2809
rect 8027 2665 8091 2729
rect 8027 2585 8091 2649
rect 8027 2505 8091 2569
rect 8027 2425 8091 2489
rect 8027 2345 8091 2409
rect 8027 2265 8091 2329
rect 7524 2045 7588 2109
rect 7604 2045 7668 2109
rect 7684 2045 7748 2109
rect 7764 2045 7828 2109
rect 7844 2045 7908 2109
rect 7924 2086 7988 2109
rect 7924 2045 7977 2086
rect 7977 2045 7988 2086
rect 8153 2985 8217 3049
rect 8153 2905 8217 2969
rect 8153 2825 8217 2889
rect 8153 2745 8217 2809
rect 8153 2665 8217 2729
rect 8153 2585 8217 2649
rect 8153 2505 8217 2569
rect 8153 2425 8217 2489
rect 8153 2345 8217 2409
rect 8153 2265 8217 2329
rect 8759 2985 8823 3049
rect 8759 2905 8823 2969
rect 8759 2825 8823 2889
rect 8759 2745 8823 2809
rect 8759 2665 8823 2729
rect 8759 2585 8823 2649
rect 8759 2505 8823 2569
rect 8759 2425 8823 2489
rect 8759 2345 8823 2409
rect 8759 2265 8823 2329
rect 9365 2985 9429 3049
rect 9365 2905 9429 2969
rect 9365 2825 9429 2889
rect 9365 2745 9429 2809
rect 9365 2665 9429 2729
rect 9365 2585 9429 2649
rect 9365 2505 9429 2569
rect 9365 2425 9429 2489
rect 9365 2345 9429 2409
rect 9365 2265 9429 2329
rect 9971 2985 10035 3049
rect 9971 2905 10035 2969
rect 9971 2825 10035 2889
rect 9971 2745 10035 2809
rect 9971 2665 10035 2729
rect 9971 2585 10035 2649
rect 9971 2505 10035 2569
rect 9971 2425 10035 2489
rect 9971 2345 10035 2409
rect 9971 2265 10035 2329
rect 10577 2985 10641 3049
rect 10577 2905 10641 2969
rect 10577 2825 10641 2889
rect 10577 2745 10641 2809
rect 10577 2665 10641 2729
rect 10577 2585 10641 2649
rect 10577 2505 10641 2569
rect 10577 2425 10641 2489
rect 10577 2345 10641 2409
rect 10577 2265 10641 2329
rect 11183 2985 11247 3049
rect 11183 2905 11247 2969
rect 11183 2825 11247 2889
rect 11183 2745 11247 2809
rect 11183 2665 11247 2729
rect 11183 2585 11247 2649
rect 11183 2505 11247 2569
rect 11183 2425 11247 2489
rect 11183 2345 11247 2409
rect 11183 2265 11247 2329
rect 11789 2985 11853 3049
rect 11789 2905 11853 2969
rect 11789 2825 11853 2889
rect 11789 2745 11853 2809
rect 11789 2665 11853 2729
rect 11789 2585 11853 2649
rect 11789 2505 11853 2569
rect 11789 2425 11853 2489
rect 11789 2345 11853 2409
rect 11789 2265 11853 2329
rect 12395 2985 12459 3049
rect 12395 2905 12459 2969
rect 12395 2825 12459 2889
rect 12395 2745 12459 2809
rect 12395 2665 12459 2729
rect 12395 2585 12459 2649
rect 12395 2505 12459 2569
rect 12395 2425 12459 2489
rect 12395 2345 12459 2409
rect 12395 2265 12459 2329
rect 13001 2985 13065 3049
rect 13001 2905 13065 2969
rect 13001 2825 13065 2889
rect 13001 2745 13065 2809
rect 13001 2665 13065 2729
rect 13001 2585 13065 2649
rect 13001 2505 13065 2569
rect 13001 2425 13065 2489
rect 13001 2345 13065 2409
rect 13001 2265 13065 2329
rect 13159 2345 13223 2349
rect 13159 2289 13163 2345
rect 13163 2289 13219 2345
rect 13219 2289 13223 2345
rect 13159 2285 13223 2289
rect 8256 2045 8320 2109
rect 8336 2045 8400 2109
rect 8416 2045 8480 2109
rect 8496 2045 8560 2109
rect 8576 2045 8640 2109
rect 8656 2086 8720 2109
rect 8656 2045 8709 2086
rect 8709 2045 8720 2086
rect 8862 2086 8926 2109
rect 8862 2045 8873 2086
rect 8873 2045 8926 2086
rect 8942 2045 9006 2109
rect 9022 2045 9086 2109
rect 9102 2045 9166 2109
rect 9182 2045 9246 2109
rect 9262 2045 9326 2109
rect 9468 2045 9532 2109
rect 9548 2045 9612 2109
rect 9628 2045 9692 2109
rect 9708 2045 9772 2109
rect 9788 2045 9852 2109
rect 9868 2086 9932 2109
rect 9868 2045 9921 2086
rect 9921 2045 9932 2086
rect 10074 2086 10138 2109
rect 10074 2045 10085 2086
rect 10085 2045 10138 2086
rect 10154 2045 10218 2109
rect 10234 2045 10298 2109
rect 10314 2045 10378 2109
rect 10394 2045 10458 2109
rect 10474 2045 10538 2109
rect 10680 2045 10744 2109
rect 10760 2045 10824 2109
rect 10840 2045 10904 2109
rect 10920 2045 10984 2109
rect 11000 2045 11064 2109
rect 11080 2086 11144 2109
rect 11080 2045 11133 2086
rect 11133 2045 11144 2086
rect 11286 2086 11350 2109
rect 11286 2045 11297 2086
rect 11297 2045 11350 2086
rect 11366 2045 11430 2109
rect 11446 2045 11510 2109
rect 11526 2045 11590 2109
rect 11606 2045 11670 2109
rect 11686 2045 11750 2109
rect 11892 2045 11956 2109
rect 11972 2045 12036 2109
rect 12052 2045 12116 2109
rect 12132 2045 12196 2109
rect 12212 2045 12276 2109
rect 12292 2086 12356 2109
rect 12292 2045 12345 2086
rect 12345 2045 12356 2086
rect 12498 2086 12562 2109
rect 12498 2045 12509 2086
rect 12509 2045 12562 2086
rect 12578 2045 12642 2109
rect 12658 2045 12722 2109
rect 12738 2045 12802 2109
rect 12818 2045 12882 2109
rect 12898 2045 12962 2109
rect 13247 2084 13311 2088
rect 13247 2028 13251 2084
rect 13251 2028 13307 2084
rect 13307 2028 13311 2084
rect 13247 2024 13311 2028
rect 1189 1796 1253 1860
rect 1269 1796 1333 1860
rect 1349 1796 1413 1860
rect 1429 1796 1493 1860
rect 1509 1796 1573 1860
rect 1589 1820 1646 1860
rect 1646 1820 1653 1860
rect 1589 1796 1653 1820
rect 1086 1576 1150 1640
rect 1086 1496 1150 1560
rect 1086 1416 1150 1480
rect 1086 1336 1150 1400
rect 1086 1256 1150 1320
rect 1086 1176 1150 1240
rect 1086 1096 1150 1160
rect 1086 1016 1150 1080
rect 1086 936 1150 1000
rect 1086 856 1150 920
rect 1692 1576 1756 1640
rect 1692 1496 1756 1560
rect 1692 1416 1756 1480
rect 1692 1336 1756 1400
rect 1692 1256 1756 1320
rect 1692 1176 1756 1240
rect 1692 1096 1756 1160
rect 1692 1016 1756 1080
rect 1692 936 1756 1000
rect 1692 856 1756 920
rect 1921 1796 1985 1860
rect 2001 1796 2065 1860
rect 2081 1796 2145 1860
rect 2161 1796 2225 1860
rect 2241 1796 2305 1860
rect 2321 1820 2378 1860
rect 2378 1820 2385 1860
rect 2321 1796 2385 1820
rect 2527 1820 2534 1860
rect 2534 1820 2591 1860
rect 2527 1796 2591 1820
rect 2607 1796 2671 1860
rect 2687 1796 2751 1860
rect 2767 1796 2831 1860
rect 2847 1796 2911 1860
rect 2927 1796 2991 1860
rect 3133 1796 3197 1860
rect 3213 1796 3277 1860
rect 3293 1796 3357 1860
rect 3373 1796 3437 1860
rect 3453 1796 3517 1860
rect 3533 1820 3590 1860
rect 3590 1820 3597 1860
rect 3533 1796 3597 1820
rect 3739 1820 3746 1860
rect 3746 1820 3803 1860
rect 3739 1796 3803 1820
rect 3819 1796 3883 1860
rect 3899 1796 3963 1860
rect 3979 1796 4043 1860
rect 4059 1796 4123 1860
rect 4139 1796 4203 1860
rect 1818 1576 1882 1640
rect 1818 1496 1882 1560
rect 1818 1416 1882 1480
rect 1818 1336 1882 1400
rect 1818 1256 1882 1320
rect 1818 1176 1882 1240
rect 1818 1096 1882 1160
rect 1818 1016 1882 1080
rect 1818 936 1882 1000
rect 1818 856 1882 920
rect 2424 1576 2488 1640
rect 2424 1496 2488 1560
rect 2424 1416 2488 1480
rect 2424 1336 2488 1400
rect 2424 1256 2488 1320
rect 2424 1176 2488 1240
rect 2424 1096 2488 1160
rect 2424 1016 2488 1080
rect 2424 936 2488 1000
rect 2424 856 2488 920
rect 3030 1576 3094 1640
rect 3030 1496 3094 1560
rect 3030 1416 3094 1480
rect 3030 1336 3094 1400
rect 3030 1256 3094 1320
rect 3030 1176 3094 1240
rect 3030 1096 3094 1160
rect 3030 1016 3094 1080
rect 3030 936 3094 1000
rect 3030 856 3094 920
rect 3636 1576 3700 1640
rect 3636 1496 3700 1560
rect 3636 1416 3700 1480
rect 3636 1336 3700 1400
rect 3636 1256 3700 1320
rect 3636 1176 3700 1240
rect 3636 1096 3700 1160
rect 3636 1016 3700 1080
rect 3636 936 3700 1000
rect 3636 856 3700 920
rect 4242 1576 4306 1640
rect 4242 1496 4306 1560
rect 4242 1416 4306 1480
rect 4242 1336 4306 1400
rect 4242 1256 4306 1320
rect 4242 1176 4306 1240
rect 4242 1096 4306 1160
rect 4242 1016 4306 1080
rect 4242 936 4306 1000
rect 4242 856 4306 920
rect 4471 1796 4535 1860
rect 4551 1796 4615 1860
rect 4631 1796 4695 1860
rect 4711 1796 4775 1860
rect 4791 1796 4855 1860
rect 4871 1820 4928 1860
rect 4928 1820 4935 1860
rect 4871 1796 4935 1820
rect 5077 1820 5084 1860
rect 5084 1820 5141 1860
rect 5077 1796 5141 1820
rect 5157 1796 5221 1860
rect 5237 1796 5301 1860
rect 5317 1796 5381 1860
rect 5397 1796 5461 1860
rect 5477 1796 5541 1860
rect 4368 1576 4432 1640
rect 4368 1496 4432 1560
rect 4368 1416 4432 1480
rect 4368 1336 4432 1400
rect 4368 1256 4432 1320
rect 4368 1176 4432 1240
rect 4368 1096 4432 1160
rect 4368 1016 4432 1080
rect 4368 936 4432 1000
rect 4368 856 4432 920
rect 4974 1576 5038 1640
rect 4974 1496 5038 1560
rect 4974 1416 5038 1480
rect 4974 1336 5038 1400
rect 4974 1256 5038 1320
rect 4974 1176 5038 1240
rect 4974 1096 5038 1160
rect 4974 1016 5038 1080
rect 4974 936 5038 1000
rect 4974 856 5038 920
rect 5580 1576 5644 1640
rect 5580 1496 5644 1560
rect 5580 1416 5644 1480
rect 5580 1336 5644 1400
rect 5580 1256 5644 1320
rect 5580 1176 5644 1240
rect 5580 1096 5644 1160
rect 5580 1016 5644 1080
rect 5580 936 5644 1000
rect 5580 856 5644 920
rect 5809 1820 5816 1860
rect 5816 1820 5873 1860
rect 5809 1796 5873 1820
rect 5889 1796 5953 1860
rect 5969 1796 6033 1860
rect 6049 1796 6113 1860
rect 6129 1796 6193 1860
rect 6209 1796 6273 1860
rect 6558 1881 6622 1885
rect 6558 1825 6562 1881
rect 6562 1825 6618 1881
rect 6618 1825 6622 1881
rect 6558 1821 6622 1825
rect 5706 1576 5770 1640
rect 5706 1496 5770 1560
rect 5706 1416 5770 1480
rect 5706 1336 5770 1400
rect 5706 1256 5770 1320
rect 5706 1176 5770 1240
rect 5706 1096 5770 1160
rect 5706 1016 5770 1080
rect 5706 936 5770 1000
rect 5706 856 5770 920
rect 6312 1576 6376 1640
rect 7878 1796 7942 1860
rect 7958 1796 8022 1860
rect 8038 1796 8102 1860
rect 8118 1796 8182 1860
rect 8198 1796 8262 1860
rect 8278 1820 8335 1860
rect 8335 1820 8342 1860
rect 8278 1796 8342 1820
rect 6312 1496 6376 1560
rect 6467 1619 6531 1623
rect 6467 1563 6471 1619
rect 6471 1563 6527 1619
rect 6527 1563 6531 1619
rect 6467 1559 6531 1563
rect 7775 1576 7839 1640
rect 6312 1416 6376 1480
rect 6312 1336 6376 1400
rect 6312 1256 6376 1320
rect 6312 1176 6376 1240
rect 6312 1096 6376 1160
rect 6312 1016 6376 1080
rect 6312 936 6376 1000
rect 6312 856 6376 920
rect 7775 1496 7839 1560
rect 7775 1416 7839 1480
rect 7775 1336 7839 1400
rect 7775 1256 7839 1320
rect 7775 1176 7839 1240
rect 7775 1096 7839 1160
rect 7775 1016 7839 1080
rect 7775 936 7839 1000
rect 7775 856 7839 920
rect 724 694 788 698
rect 724 638 728 694
rect 728 638 784 694
rect 784 638 788 694
rect 724 634 788 638
rect 1189 636 1253 700
rect 1269 636 1333 700
rect 1349 636 1413 700
rect 1429 636 1493 700
rect 1509 636 1573 700
rect 1589 636 1653 700
rect 1921 636 1985 700
rect 2001 636 2065 700
rect 2081 636 2145 700
rect 2161 636 2225 700
rect 2241 636 2305 700
rect 2321 636 2385 700
rect 2527 636 2591 700
rect 2607 636 2671 700
rect 2687 636 2751 700
rect 2767 636 2831 700
rect 2847 636 2911 700
rect 2927 636 2991 700
rect 3133 636 3197 700
rect 3213 636 3277 700
rect 3293 636 3357 700
rect 3373 636 3437 700
rect 3453 636 3517 700
rect 3533 636 3597 700
rect 3739 636 3803 700
rect 3819 636 3883 700
rect 3899 636 3963 700
rect 3979 636 4043 700
rect 4059 636 4123 700
rect 4139 636 4203 700
rect 4471 636 4535 700
rect 4551 636 4615 700
rect 4631 636 4695 700
rect 4711 636 4775 700
rect 4791 636 4855 700
rect 4871 636 4935 700
rect 5077 636 5141 700
rect 5157 636 5221 700
rect 5237 636 5301 700
rect 5317 636 5381 700
rect 5397 636 5461 700
rect 5477 636 5541 700
rect 5809 636 5873 700
rect 5889 636 5953 700
rect 5969 636 6033 700
rect 6049 636 6113 700
rect 6129 636 6193 700
rect 6209 636 6273 700
rect 8381 1576 8445 1640
rect 8381 1496 8445 1560
rect 8381 1416 8445 1480
rect 8381 1336 8445 1400
rect 8381 1256 8445 1320
rect 8381 1176 8445 1240
rect 8381 1096 8445 1160
rect 8381 1016 8445 1080
rect 8381 936 8445 1000
rect 8381 856 8445 920
rect 8610 1796 8674 1860
rect 8690 1796 8754 1860
rect 8770 1796 8834 1860
rect 8850 1796 8914 1860
rect 8930 1796 8994 1860
rect 9010 1820 9067 1860
rect 9067 1820 9074 1860
rect 9010 1796 9074 1820
rect 9216 1820 9223 1860
rect 9223 1820 9280 1860
rect 9216 1796 9280 1820
rect 9296 1796 9360 1860
rect 9376 1796 9440 1860
rect 9456 1796 9520 1860
rect 9536 1796 9600 1860
rect 9616 1796 9680 1860
rect 9822 1796 9886 1860
rect 9902 1796 9966 1860
rect 9982 1796 10046 1860
rect 10062 1796 10126 1860
rect 10142 1796 10206 1860
rect 10222 1820 10279 1860
rect 10279 1820 10286 1860
rect 10222 1796 10286 1820
rect 10428 1820 10435 1860
rect 10435 1820 10492 1860
rect 10428 1796 10492 1820
rect 10508 1796 10572 1860
rect 10588 1796 10652 1860
rect 10668 1796 10732 1860
rect 10748 1796 10812 1860
rect 10828 1796 10892 1860
rect 8507 1576 8571 1640
rect 8507 1496 8571 1560
rect 8507 1416 8571 1480
rect 8507 1336 8571 1400
rect 8507 1256 8571 1320
rect 8507 1176 8571 1240
rect 8507 1096 8571 1160
rect 8507 1016 8571 1080
rect 8507 936 8571 1000
rect 8507 856 8571 920
rect 9113 1576 9177 1640
rect 9113 1496 9177 1560
rect 9113 1416 9177 1480
rect 9113 1336 9177 1400
rect 9113 1256 9177 1320
rect 9113 1176 9177 1240
rect 9113 1096 9177 1160
rect 9113 1016 9177 1080
rect 9113 936 9177 1000
rect 9113 856 9177 920
rect 9719 1576 9783 1640
rect 9719 1496 9783 1560
rect 9719 1416 9783 1480
rect 9719 1336 9783 1400
rect 9719 1256 9783 1320
rect 9719 1176 9783 1240
rect 9719 1096 9783 1160
rect 9719 1016 9783 1080
rect 9719 936 9783 1000
rect 9719 856 9783 920
rect 10325 1576 10389 1640
rect 10325 1496 10389 1560
rect 10325 1416 10389 1480
rect 10325 1336 10389 1400
rect 10325 1256 10389 1320
rect 10325 1176 10389 1240
rect 10325 1096 10389 1160
rect 10325 1016 10389 1080
rect 10325 936 10389 1000
rect 10325 856 10389 920
rect 10931 1576 10995 1640
rect 10931 1496 10995 1560
rect 10931 1416 10995 1480
rect 10931 1336 10995 1400
rect 10931 1256 10995 1320
rect 10931 1176 10995 1240
rect 10931 1096 10995 1160
rect 10931 1016 10995 1080
rect 10931 936 10995 1000
rect 10931 856 10995 920
rect 11160 1796 11224 1860
rect 11240 1796 11304 1860
rect 11320 1796 11384 1860
rect 11400 1796 11464 1860
rect 11480 1796 11544 1860
rect 11560 1820 11617 1860
rect 11617 1820 11624 1860
rect 11560 1796 11624 1820
rect 11766 1820 11773 1860
rect 11773 1820 11830 1860
rect 11766 1796 11830 1820
rect 11846 1796 11910 1860
rect 11926 1796 11990 1860
rect 12006 1796 12070 1860
rect 12086 1796 12150 1860
rect 12166 1796 12230 1860
rect 11057 1576 11121 1640
rect 11057 1496 11121 1560
rect 11057 1416 11121 1480
rect 11057 1336 11121 1400
rect 11057 1256 11121 1320
rect 11057 1176 11121 1240
rect 11057 1096 11121 1160
rect 11057 1016 11121 1080
rect 11057 936 11121 1000
rect 11057 856 11121 920
rect 11663 1576 11727 1640
rect 11663 1496 11727 1560
rect 11663 1416 11727 1480
rect 11663 1336 11727 1400
rect 11663 1256 11727 1320
rect 11663 1176 11727 1240
rect 11663 1096 11727 1160
rect 11663 1016 11727 1080
rect 11663 936 11727 1000
rect 11663 856 11727 920
rect 12269 1576 12333 1640
rect 12269 1496 12333 1560
rect 12269 1416 12333 1480
rect 12269 1336 12333 1400
rect 12269 1256 12333 1320
rect 12269 1176 12333 1240
rect 12269 1096 12333 1160
rect 12269 1016 12333 1080
rect 12269 936 12333 1000
rect 12269 856 12333 920
rect 12498 1820 12505 1860
rect 12505 1820 12562 1860
rect 12498 1796 12562 1820
rect 12578 1796 12642 1860
rect 12658 1796 12722 1860
rect 12738 1796 12802 1860
rect 12818 1796 12882 1860
rect 12898 1796 12962 1860
rect 13247 1881 13311 1885
rect 13247 1825 13251 1881
rect 13251 1825 13307 1881
rect 13307 1825 13311 1881
rect 13247 1821 13311 1825
rect 12395 1576 12459 1640
rect 12395 1496 12459 1560
rect 12395 1416 12459 1480
rect 12395 1336 12459 1400
rect 12395 1256 12459 1320
rect 12395 1176 12459 1240
rect 12395 1096 12459 1160
rect 12395 1016 12459 1080
rect 12395 936 12459 1000
rect 12395 856 12459 920
rect 13001 1576 13065 1640
rect 13001 1496 13065 1560
rect 13156 1619 13220 1623
rect 13156 1563 13160 1619
rect 13160 1563 13216 1619
rect 13216 1563 13220 1619
rect 13156 1559 13220 1563
rect 13001 1416 13065 1480
rect 13001 1336 13065 1400
rect 13001 1256 13065 1320
rect 13001 1176 13065 1240
rect 13001 1096 13065 1160
rect 13001 1016 13065 1080
rect 13001 936 13065 1000
rect 13001 856 13065 920
rect 7413 694 7477 698
rect 7413 638 7417 694
rect 7417 638 7473 694
rect 7473 638 7477 694
rect 7413 634 7477 638
rect 7878 636 7942 700
rect 7958 636 8022 700
rect 8038 636 8102 700
rect 8118 636 8182 700
rect 8198 636 8262 700
rect 8278 636 8342 700
rect 8610 636 8674 700
rect 8690 636 8754 700
rect 8770 636 8834 700
rect 8850 636 8914 700
rect 8930 636 8994 700
rect 9010 636 9074 700
rect 9216 636 9280 700
rect 9296 636 9360 700
rect 9376 636 9440 700
rect 9456 636 9520 700
rect 9536 636 9600 700
rect 9616 636 9680 700
rect 9822 636 9886 700
rect 9902 636 9966 700
rect 9982 636 10046 700
rect 10062 636 10126 700
rect 10142 636 10206 700
rect 10222 636 10286 700
rect 10428 636 10492 700
rect 10508 636 10572 700
rect 10588 636 10652 700
rect 10668 636 10732 700
rect 10748 636 10812 700
rect 10828 636 10892 700
rect 11160 636 11224 700
rect 11240 636 11304 700
rect 11320 636 11384 700
rect 11400 636 11464 700
rect 11480 636 11544 700
rect 11560 636 11624 700
rect 11766 636 11830 700
rect 11846 636 11910 700
rect 11926 636 11990 700
rect 12006 636 12070 700
rect 12086 636 12150 700
rect 12166 636 12230 700
rect 12498 636 12562 700
rect 12578 636 12642 700
rect 12658 636 12722 700
rect 12738 636 12802 700
rect 12818 636 12882 700
rect 12898 636 12962 700
rect 576 248 640 312
rect 656 248 720 312
rect 736 248 800 312
rect 816 248 880 312
rect 896 248 960 312
rect 976 248 1040 312
rect 1308 248 1372 312
rect 1388 248 1452 312
rect 1468 248 1532 312
rect 1548 248 1612 312
rect 1628 248 1692 312
rect 1708 248 1772 312
rect 1914 248 1978 312
rect 1994 248 2058 312
rect 2074 248 2138 312
rect 2154 248 2218 312
rect 2234 248 2298 312
rect 2314 248 2378 312
rect 2646 248 2710 312
rect 2726 248 2790 312
rect 2806 248 2870 312
rect 2886 248 2950 312
rect 2966 248 3030 312
rect 3046 248 3110 312
rect 3252 248 3316 312
rect 3332 248 3396 312
rect 3412 248 3476 312
rect 3492 248 3556 312
rect 3572 248 3636 312
rect 3652 248 3716 312
rect 3858 248 3922 312
rect 3938 248 4002 312
rect 4018 248 4082 312
rect 4098 248 4162 312
rect 4178 248 4242 312
rect 4258 248 4322 312
rect 4464 248 4528 312
rect 4544 248 4608 312
rect 4624 248 4688 312
rect 4704 248 4768 312
rect 4784 248 4848 312
rect 4864 248 4928 312
rect 5196 248 5260 312
rect 5276 248 5340 312
rect 5356 248 5420 312
rect 5436 248 5500 312
rect 5516 248 5580 312
rect 5596 248 5660 312
rect 6061 310 6125 314
rect 6061 254 6065 310
rect 6065 254 6121 310
rect 6121 254 6125 310
rect 6061 250 6125 254
rect 473 28 537 92
rect 473 -52 537 12
rect 473 -132 537 -68
rect 473 -212 537 -148
rect 473 -292 537 -228
rect 473 -372 537 -308
rect 473 -452 537 -388
rect 473 -532 537 -468
rect 318 -615 382 -611
rect 318 -671 322 -615
rect 322 -671 378 -615
rect 378 -671 382 -615
rect 318 -675 382 -671
rect 473 -612 537 -548
rect 473 -692 537 -628
rect 1079 28 1143 92
rect 1079 -52 1143 12
rect 1079 -132 1143 -68
rect 1079 -212 1143 -148
rect 1079 -292 1143 -228
rect 1079 -372 1143 -308
rect 1079 -452 1143 -388
rect 1079 -532 1143 -468
rect 1079 -612 1143 -548
rect 1079 -692 1143 -628
rect 227 -877 291 -873
rect 227 -933 231 -877
rect 231 -933 287 -877
rect 287 -933 291 -877
rect 227 -937 291 -933
rect 576 -912 640 -848
rect 656 -912 720 -848
rect 736 -912 800 -848
rect 816 -912 880 -848
rect 896 -912 960 -848
rect 976 -872 1040 -848
rect 976 -912 1033 -872
rect 1033 -912 1040 -872
rect 1205 28 1269 92
rect 1205 -52 1269 12
rect 1205 -132 1269 -68
rect 1205 -212 1269 -148
rect 1205 -292 1269 -228
rect 1205 -372 1269 -308
rect 1205 -452 1269 -388
rect 1205 -532 1269 -468
rect 1205 -612 1269 -548
rect 1205 -692 1269 -628
rect 1811 28 1875 92
rect 1811 -52 1875 12
rect 1811 -132 1875 -68
rect 1811 -212 1875 -148
rect 1811 -292 1875 -228
rect 1811 -372 1875 -308
rect 1811 -452 1875 -388
rect 1811 -532 1875 -468
rect 1811 -612 1875 -548
rect 1811 -692 1875 -628
rect 2417 28 2481 92
rect 2417 -52 2481 12
rect 2417 -132 2481 -68
rect 2417 -212 2481 -148
rect 2417 -292 2481 -228
rect 2417 -372 2481 -308
rect 2417 -452 2481 -388
rect 2417 -532 2481 -468
rect 2417 -612 2481 -548
rect 2417 -692 2481 -628
rect 1308 -912 1372 -848
rect 1388 -912 1452 -848
rect 1468 -912 1532 -848
rect 1548 -912 1612 -848
rect 1628 -912 1692 -848
rect 1708 -872 1772 -848
rect 1708 -912 1765 -872
rect 1765 -912 1772 -872
rect 1914 -872 1978 -848
rect 1914 -912 1921 -872
rect 1921 -912 1978 -872
rect 1994 -912 2058 -848
rect 2074 -912 2138 -848
rect 2154 -912 2218 -848
rect 2234 -912 2298 -848
rect 2314 -912 2378 -848
rect 2543 28 2607 92
rect 2543 -52 2607 12
rect 2543 -132 2607 -68
rect 2543 -212 2607 -148
rect 2543 -292 2607 -228
rect 2543 -372 2607 -308
rect 2543 -452 2607 -388
rect 2543 -532 2607 -468
rect 2543 -612 2607 -548
rect 2543 -692 2607 -628
rect 3149 28 3213 92
rect 3149 -52 3213 12
rect 3149 -132 3213 -68
rect 3149 -212 3213 -148
rect 3149 -292 3213 -228
rect 3149 -372 3213 -308
rect 3149 -452 3213 -388
rect 3149 -532 3213 -468
rect 3149 -612 3213 -548
rect 3149 -692 3213 -628
rect 3755 28 3819 92
rect 3755 -52 3819 12
rect 3755 -132 3819 -68
rect 3755 -212 3819 -148
rect 3755 -292 3819 -228
rect 3755 -372 3819 -308
rect 3755 -452 3819 -388
rect 3755 -532 3819 -468
rect 3755 -612 3819 -548
rect 3755 -692 3819 -628
rect 4361 28 4425 92
rect 4361 -52 4425 12
rect 4361 -132 4425 -68
rect 4361 -212 4425 -148
rect 4361 -292 4425 -228
rect 4361 -372 4425 -308
rect 4361 -452 4425 -388
rect 4361 -532 4425 -468
rect 4361 -612 4425 -548
rect 4361 -692 4425 -628
rect 4967 28 5031 92
rect 4967 -52 5031 12
rect 4967 -132 5031 -68
rect 4967 -212 5031 -148
rect 4967 -292 5031 -228
rect 4967 -372 5031 -308
rect 4967 -452 5031 -388
rect 4967 -532 5031 -468
rect 4967 -612 5031 -548
rect 4967 -692 5031 -628
rect 2646 -912 2710 -848
rect 2726 -912 2790 -848
rect 2806 -912 2870 -848
rect 2886 -912 2950 -848
rect 2966 -912 3030 -848
rect 3046 -872 3110 -848
rect 3046 -912 3103 -872
rect 3103 -912 3110 -872
rect 3252 -872 3316 -848
rect 3252 -912 3259 -872
rect 3259 -912 3316 -872
rect 3332 -912 3396 -848
rect 3412 -912 3476 -848
rect 3492 -912 3556 -848
rect 3572 -912 3636 -848
rect 3652 -912 3716 -848
rect 3858 -912 3922 -848
rect 3938 -912 4002 -848
rect 4018 -912 4082 -848
rect 4098 -912 4162 -848
rect 4178 -912 4242 -848
rect 4258 -872 4322 -848
rect 4258 -912 4315 -872
rect 4315 -912 4322 -872
rect 4464 -872 4528 -848
rect 4464 -912 4471 -872
rect 4471 -912 4528 -872
rect 4544 -912 4608 -848
rect 4624 -912 4688 -848
rect 4704 -912 4768 -848
rect 4784 -912 4848 -848
rect 4864 -912 4928 -848
rect 5093 28 5157 92
rect 5093 -52 5157 12
rect 5093 -132 5157 -68
rect 5093 -212 5157 -148
rect 5093 -292 5157 -228
rect 5093 -372 5157 -308
rect 5093 -452 5157 -388
rect 5093 -532 5157 -468
rect 5093 -612 5157 -548
rect 5093 -692 5157 -628
rect 7331 248 7395 312
rect 7411 248 7475 312
rect 7491 248 7555 312
rect 7571 248 7635 312
rect 7651 248 7715 312
rect 7731 248 7795 312
rect 8063 248 8127 312
rect 8143 248 8207 312
rect 8223 248 8287 312
rect 8303 248 8367 312
rect 8383 248 8447 312
rect 8463 248 8527 312
rect 8669 248 8733 312
rect 8749 248 8813 312
rect 8829 248 8893 312
rect 8909 248 8973 312
rect 8989 248 9053 312
rect 9069 248 9133 312
rect 9401 248 9465 312
rect 9481 248 9545 312
rect 9561 248 9625 312
rect 9641 248 9705 312
rect 9721 248 9785 312
rect 9801 248 9865 312
rect 10007 248 10071 312
rect 10087 248 10151 312
rect 10167 248 10231 312
rect 10247 248 10311 312
rect 10327 248 10391 312
rect 10407 248 10471 312
rect 10613 248 10677 312
rect 10693 248 10757 312
rect 10773 248 10837 312
rect 10853 248 10917 312
rect 10933 248 10997 312
rect 11013 248 11077 312
rect 11219 248 11283 312
rect 11299 248 11363 312
rect 11379 248 11443 312
rect 11459 248 11523 312
rect 11539 248 11603 312
rect 11619 248 11683 312
rect 11951 248 12015 312
rect 12031 248 12095 312
rect 12111 248 12175 312
rect 12191 248 12255 312
rect 12271 248 12335 312
rect 12351 248 12415 312
rect 12816 310 12880 314
rect 12816 254 12820 310
rect 12820 254 12876 310
rect 12876 254 12880 310
rect 12816 250 12880 254
rect 5699 28 5763 92
rect 5699 -52 5763 12
rect 5699 -132 5763 -68
rect 5699 -212 5763 -148
rect 5699 -292 5763 -228
rect 5699 -372 5763 -308
rect 5699 -452 5763 -388
rect 5699 -532 5763 -468
rect 5699 -612 5763 -548
rect 7228 28 7292 92
rect 7228 -52 7292 12
rect 7228 -132 7292 -68
rect 7228 -212 7292 -148
rect 7228 -292 7292 -228
rect 7228 -372 7292 -308
rect 7228 -452 7292 -388
rect 7228 -532 7292 -468
rect 5699 -692 5763 -628
rect 7073 -615 7137 -611
rect 7073 -671 7077 -615
rect 7077 -671 7133 -615
rect 7133 -671 7137 -615
rect 7073 -675 7137 -671
rect 7228 -612 7292 -548
rect 5196 -872 5260 -848
rect 5196 -912 5203 -872
rect 5203 -912 5260 -872
rect 5276 -912 5340 -848
rect 5356 -912 5420 -848
rect 5436 -912 5500 -848
rect 5516 -912 5580 -848
rect 5596 -912 5660 -848
rect 7228 -692 7292 -628
rect 7834 28 7898 92
rect 7834 -52 7898 12
rect 7834 -132 7898 -68
rect 7834 -212 7898 -148
rect 7834 -292 7898 -228
rect 7834 -372 7898 -308
rect 7834 -452 7898 -388
rect 7834 -532 7898 -468
rect 7834 -612 7898 -548
rect 7834 -692 7898 -628
rect 6982 -877 7046 -873
rect 6982 -933 6986 -877
rect 6986 -933 7042 -877
rect 7042 -933 7046 -877
rect 6982 -937 7046 -933
rect 7331 -912 7395 -848
rect 7411 -912 7475 -848
rect 7491 -912 7555 -848
rect 7571 -912 7635 -848
rect 7651 -912 7715 -848
rect 7731 -872 7795 -848
rect 7731 -912 7788 -872
rect 7788 -912 7795 -872
rect 7960 28 8024 92
rect 7960 -52 8024 12
rect 7960 -132 8024 -68
rect 7960 -212 8024 -148
rect 7960 -292 8024 -228
rect 7960 -372 8024 -308
rect 7960 -452 8024 -388
rect 7960 -532 8024 -468
rect 7960 -612 8024 -548
rect 7960 -692 8024 -628
rect 8566 28 8630 92
rect 8566 -52 8630 12
rect 8566 -132 8630 -68
rect 8566 -212 8630 -148
rect 8566 -292 8630 -228
rect 8566 -372 8630 -308
rect 8566 -452 8630 -388
rect 8566 -532 8630 -468
rect 8566 -612 8630 -548
rect 8566 -692 8630 -628
rect 9172 28 9236 92
rect 9172 -52 9236 12
rect 9172 -132 9236 -68
rect 9172 -212 9236 -148
rect 9172 -292 9236 -228
rect 9172 -372 9236 -308
rect 9172 -452 9236 -388
rect 9172 -532 9236 -468
rect 9172 -612 9236 -548
rect 9172 -692 9236 -628
rect 8063 -912 8127 -848
rect 8143 -912 8207 -848
rect 8223 -912 8287 -848
rect 8303 -912 8367 -848
rect 8383 -912 8447 -848
rect 8463 -872 8527 -848
rect 8463 -912 8520 -872
rect 8520 -912 8527 -872
rect 8669 -872 8733 -848
rect 8669 -912 8676 -872
rect 8676 -912 8733 -872
rect 8749 -912 8813 -848
rect 8829 -912 8893 -848
rect 8909 -912 8973 -848
rect 8989 -912 9053 -848
rect 9069 -912 9133 -848
rect 9298 28 9362 92
rect 9298 -52 9362 12
rect 9298 -132 9362 -68
rect 9298 -212 9362 -148
rect 9298 -292 9362 -228
rect 9298 -372 9362 -308
rect 9298 -452 9362 -388
rect 9298 -532 9362 -468
rect 9298 -612 9362 -548
rect 9298 -692 9362 -628
rect 9904 28 9968 92
rect 9904 -52 9968 12
rect 9904 -132 9968 -68
rect 9904 -212 9968 -148
rect 9904 -292 9968 -228
rect 9904 -372 9968 -308
rect 9904 -452 9968 -388
rect 9904 -532 9968 -468
rect 9904 -612 9968 -548
rect 9904 -692 9968 -628
rect 10510 28 10574 92
rect 10510 -52 10574 12
rect 10510 -132 10574 -68
rect 10510 -212 10574 -148
rect 10510 -292 10574 -228
rect 10510 -372 10574 -308
rect 10510 -452 10574 -388
rect 10510 -532 10574 -468
rect 10510 -612 10574 -548
rect 10510 -692 10574 -628
rect 11116 28 11180 92
rect 11116 -52 11180 12
rect 11116 -132 11180 -68
rect 11116 -212 11180 -148
rect 11116 -292 11180 -228
rect 11116 -372 11180 -308
rect 11116 -452 11180 -388
rect 11116 -532 11180 -468
rect 11116 -612 11180 -548
rect 11116 -692 11180 -628
rect 11722 28 11786 92
rect 11722 -52 11786 12
rect 11722 -132 11786 -68
rect 11722 -212 11786 -148
rect 11722 -292 11786 -228
rect 11722 -372 11786 -308
rect 11722 -452 11786 -388
rect 11722 -532 11786 -468
rect 11722 -612 11786 -548
rect 11722 -692 11786 -628
rect 9401 -912 9465 -848
rect 9481 -912 9545 -848
rect 9561 -912 9625 -848
rect 9641 -912 9705 -848
rect 9721 -912 9785 -848
rect 9801 -872 9865 -848
rect 9801 -912 9858 -872
rect 9858 -912 9865 -872
rect 10007 -872 10071 -848
rect 10007 -912 10014 -872
rect 10014 -912 10071 -872
rect 10087 -912 10151 -848
rect 10167 -912 10231 -848
rect 10247 -912 10311 -848
rect 10327 -912 10391 -848
rect 10407 -912 10471 -848
rect 10613 -912 10677 -848
rect 10693 -912 10757 -848
rect 10773 -912 10837 -848
rect 10853 -912 10917 -848
rect 10933 -912 10997 -848
rect 11013 -872 11077 -848
rect 11013 -912 11070 -872
rect 11070 -912 11077 -872
rect 11219 -872 11283 -848
rect 11219 -912 11226 -872
rect 11226 -912 11283 -872
rect 11299 -912 11363 -848
rect 11379 -912 11443 -848
rect 11459 -912 11523 -848
rect 11539 -912 11603 -848
rect 11619 -912 11683 -848
rect 11848 28 11912 92
rect 11848 -52 11912 12
rect 11848 -132 11912 -68
rect 11848 -212 11912 -148
rect 11848 -292 11912 -228
rect 11848 -372 11912 -308
rect 11848 -452 11912 -388
rect 11848 -532 11912 -468
rect 11848 -612 11912 -548
rect 11848 -692 11912 -628
rect 12454 28 12518 92
rect 12454 -52 12518 12
rect 12454 -132 12518 -68
rect 12454 -212 12518 -148
rect 12454 -292 12518 -228
rect 12454 -372 12518 -308
rect 12454 -452 12518 -388
rect 12454 -532 12518 -468
rect 12454 -612 12518 -548
rect 12454 -692 12518 -628
rect 11951 -872 12015 -848
rect 11951 -912 11958 -872
rect 11958 -912 12015 -872
rect 12031 -912 12095 -848
rect 12111 -912 12175 -848
rect 12191 -912 12255 -848
rect 12271 -912 12335 -848
rect 12351 -912 12415 -848
rect 227 -1080 291 -1076
rect 227 -1136 231 -1080
rect 231 -1136 287 -1080
rect 287 -1136 291 -1080
rect 227 -1140 291 -1136
rect 576 -1161 640 -1097
rect 656 -1161 720 -1097
rect 736 -1161 800 -1097
rect 816 -1161 880 -1097
rect 896 -1161 960 -1097
rect 976 -1138 1029 -1097
rect 1029 -1138 1040 -1097
rect 976 -1161 1040 -1138
rect 1182 -1138 1193 -1097
rect 1193 -1138 1246 -1097
rect 1182 -1161 1246 -1138
rect 1262 -1161 1326 -1097
rect 1342 -1161 1406 -1097
rect 1422 -1161 1486 -1097
rect 1502 -1161 1566 -1097
rect 1582 -1161 1646 -1097
rect 1788 -1161 1852 -1097
rect 1868 -1161 1932 -1097
rect 1948 -1161 2012 -1097
rect 2028 -1161 2092 -1097
rect 2108 -1161 2172 -1097
rect 2188 -1138 2241 -1097
rect 2241 -1138 2252 -1097
rect 2188 -1161 2252 -1138
rect 2394 -1138 2405 -1097
rect 2405 -1138 2458 -1097
rect 2394 -1161 2458 -1138
rect 2474 -1161 2538 -1097
rect 2554 -1161 2618 -1097
rect 2634 -1161 2698 -1097
rect 2714 -1161 2778 -1097
rect 2794 -1161 2858 -1097
rect 3000 -1161 3064 -1097
rect 3080 -1161 3144 -1097
rect 3160 -1161 3224 -1097
rect 3240 -1161 3304 -1097
rect 3320 -1161 3384 -1097
rect 3400 -1138 3453 -1097
rect 3453 -1138 3464 -1097
rect 3400 -1161 3464 -1138
rect 3606 -1138 3617 -1097
rect 3617 -1138 3670 -1097
rect 3606 -1161 3670 -1138
rect 3686 -1161 3750 -1097
rect 3766 -1161 3830 -1097
rect 3846 -1161 3910 -1097
rect 3926 -1161 3990 -1097
rect 4006 -1161 4070 -1097
rect 4212 -1161 4276 -1097
rect 4292 -1161 4356 -1097
rect 4372 -1161 4436 -1097
rect 4452 -1161 4516 -1097
rect 4532 -1161 4596 -1097
rect 4612 -1138 4665 -1097
rect 4665 -1138 4676 -1097
rect 4612 -1161 4676 -1138
rect 4818 -1138 4829 -1097
rect 4829 -1138 4882 -1097
rect 4818 -1161 4882 -1138
rect 4898 -1161 4962 -1097
rect 4978 -1161 5042 -1097
rect 5058 -1161 5122 -1097
rect 5138 -1161 5202 -1097
rect 5218 -1161 5282 -1097
rect 315 -1341 379 -1337
rect 315 -1397 319 -1341
rect 319 -1397 375 -1341
rect 375 -1397 379 -1341
rect 315 -1401 379 -1397
rect 473 -1381 537 -1317
rect 473 -1461 537 -1397
rect 473 -1541 537 -1477
rect 473 -1621 537 -1557
rect 473 -1701 537 -1637
rect 473 -1781 537 -1717
rect 473 -1861 537 -1797
rect 473 -1941 537 -1877
rect 473 -2021 537 -1957
rect 473 -2101 537 -2037
rect 1079 -1381 1143 -1317
rect 1079 -1461 1143 -1397
rect 1079 -1541 1143 -1477
rect 1079 -1621 1143 -1557
rect 1079 -1701 1143 -1637
rect 1079 -1781 1143 -1717
rect 1079 -1861 1143 -1797
rect 1079 -1941 1143 -1877
rect 1079 -2021 1143 -1957
rect 1079 -2101 1143 -2037
rect 1685 -1381 1749 -1317
rect 1685 -1461 1749 -1397
rect 1685 -1541 1749 -1477
rect 1685 -1621 1749 -1557
rect 1685 -1701 1749 -1637
rect 1685 -1781 1749 -1717
rect 1685 -1861 1749 -1797
rect 1685 -1941 1749 -1877
rect 1685 -2021 1749 -1957
rect 1685 -2101 1749 -2037
rect 2291 -1381 2355 -1317
rect 2291 -1461 2355 -1397
rect 2291 -1541 2355 -1477
rect 2291 -1621 2355 -1557
rect 2291 -1701 2355 -1637
rect 2291 -1781 2355 -1717
rect 2291 -1861 2355 -1797
rect 2291 -1941 2355 -1877
rect 2291 -2021 2355 -1957
rect 2291 -2101 2355 -2037
rect 2897 -1381 2961 -1317
rect 2897 -1461 2961 -1397
rect 2897 -1541 2961 -1477
rect 2897 -1621 2961 -1557
rect 2897 -1701 2961 -1637
rect 2897 -1781 2961 -1717
rect 2897 -1861 2961 -1797
rect 2897 -1941 2961 -1877
rect 2897 -2021 2961 -1957
rect 2897 -2101 2961 -2037
rect 3503 -1381 3567 -1317
rect 3503 -1461 3567 -1397
rect 3503 -1541 3567 -1477
rect 3503 -1621 3567 -1557
rect 3503 -1701 3567 -1637
rect 3503 -1781 3567 -1717
rect 3503 -1861 3567 -1797
rect 3503 -1941 3567 -1877
rect 3503 -2021 3567 -1957
rect 3503 -2101 3567 -2037
rect 4109 -1381 4173 -1317
rect 4109 -1461 4173 -1397
rect 4109 -1541 4173 -1477
rect 4109 -1621 4173 -1557
rect 4109 -1701 4173 -1637
rect 4109 -1781 4173 -1717
rect 4109 -1861 4173 -1797
rect 4109 -1941 4173 -1877
rect 4109 -2021 4173 -1957
rect 4109 -2101 4173 -2037
rect 4715 -1381 4779 -1317
rect 4715 -1461 4779 -1397
rect 4715 -1541 4779 -1477
rect 4715 -1621 4779 -1557
rect 4715 -1701 4779 -1637
rect 4715 -1781 4779 -1717
rect 4715 -1861 4779 -1797
rect 4715 -1941 4779 -1877
rect 4715 -2021 4779 -1957
rect 4715 -2101 4779 -2037
rect 5321 -1381 5385 -1317
rect 5321 -1461 5385 -1397
rect 5321 -1541 5385 -1477
rect 5321 -1621 5385 -1557
rect 5321 -1701 5385 -1637
rect 5321 -1781 5385 -1717
rect 5321 -1861 5385 -1797
rect 5321 -1941 5385 -1877
rect 5321 -2021 5385 -1957
rect 5321 -2101 5385 -2037
rect 5550 -1138 5561 -1097
rect 5561 -1138 5614 -1097
rect 5550 -1161 5614 -1138
rect 5630 -1161 5694 -1097
rect 5710 -1161 5774 -1097
rect 5790 -1161 5854 -1097
rect 5870 -1161 5934 -1097
rect 5950 -1161 6014 -1097
rect 5447 -1381 5511 -1317
rect 5447 -1461 5511 -1397
rect 5447 -1541 5511 -1477
rect 5447 -1621 5511 -1557
rect 5447 -1701 5511 -1637
rect 5447 -1781 5511 -1717
rect 5447 -1861 5511 -1797
rect 5447 -1941 5511 -1877
rect 5447 -2021 5511 -1957
rect 5447 -2101 5511 -2037
rect 6383 -1117 6447 -1113
rect 6383 -1173 6387 -1117
rect 6387 -1173 6443 -1117
rect 6443 -1173 6447 -1117
rect 6383 -1177 6447 -1173
rect 6526 -1117 6590 -1113
rect 6526 -1173 6530 -1117
rect 6530 -1173 6586 -1117
rect 6586 -1173 6590 -1117
rect 6526 -1177 6590 -1173
rect 6646 -1117 6710 -1113
rect 6646 -1173 6650 -1117
rect 6650 -1173 6706 -1117
rect 6706 -1173 6710 -1117
rect 6646 -1177 6710 -1173
rect 6982 -1080 7046 -1076
rect 6982 -1136 6986 -1080
rect 6986 -1136 7042 -1080
rect 7042 -1136 7046 -1080
rect 6982 -1140 7046 -1136
rect 7331 -1161 7395 -1097
rect 7411 -1161 7475 -1097
rect 7491 -1161 7555 -1097
rect 7571 -1161 7635 -1097
rect 7651 -1161 7715 -1097
rect 7731 -1138 7784 -1097
rect 7784 -1138 7795 -1097
rect 7731 -1161 7795 -1138
rect 7937 -1138 7948 -1097
rect 7948 -1138 8001 -1097
rect 7937 -1161 8001 -1138
rect 8017 -1161 8081 -1097
rect 8097 -1161 8161 -1097
rect 8177 -1161 8241 -1097
rect 8257 -1161 8321 -1097
rect 8337 -1161 8401 -1097
rect 8543 -1161 8607 -1097
rect 8623 -1161 8687 -1097
rect 8703 -1161 8767 -1097
rect 8783 -1161 8847 -1097
rect 8863 -1161 8927 -1097
rect 8943 -1138 8996 -1097
rect 8996 -1138 9007 -1097
rect 8943 -1161 9007 -1138
rect 9149 -1138 9160 -1097
rect 9160 -1138 9213 -1097
rect 9149 -1161 9213 -1138
rect 9229 -1161 9293 -1097
rect 9309 -1161 9373 -1097
rect 9389 -1161 9453 -1097
rect 9469 -1161 9533 -1097
rect 9549 -1161 9613 -1097
rect 9755 -1161 9819 -1097
rect 9835 -1161 9899 -1097
rect 9915 -1161 9979 -1097
rect 9995 -1161 10059 -1097
rect 10075 -1161 10139 -1097
rect 10155 -1138 10208 -1097
rect 10208 -1138 10219 -1097
rect 10155 -1161 10219 -1138
rect 10361 -1138 10372 -1097
rect 10372 -1138 10425 -1097
rect 10361 -1161 10425 -1138
rect 10441 -1161 10505 -1097
rect 10521 -1161 10585 -1097
rect 10601 -1161 10665 -1097
rect 10681 -1161 10745 -1097
rect 10761 -1161 10825 -1097
rect 10967 -1161 11031 -1097
rect 11047 -1161 11111 -1097
rect 11127 -1161 11191 -1097
rect 11207 -1161 11271 -1097
rect 11287 -1161 11351 -1097
rect 11367 -1138 11420 -1097
rect 11420 -1138 11431 -1097
rect 11367 -1161 11431 -1138
rect 11573 -1138 11584 -1097
rect 11584 -1138 11637 -1097
rect 11573 -1161 11637 -1138
rect 11653 -1161 11717 -1097
rect 11733 -1161 11797 -1097
rect 11813 -1161 11877 -1097
rect 11893 -1161 11957 -1097
rect 11973 -1161 12037 -1097
rect 6053 -1381 6117 -1317
rect 6053 -1461 6117 -1397
rect 7070 -1341 7134 -1337
rect 7070 -1397 7074 -1341
rect 7074 -1397 7130 -1341
rect 7130 -1397 7134 -1341
rect 7070 -1401 7134 -1397
rect 7228 -1381 7292 -1317
rect 6053 -1541 6117 -1477
rect 6053 -1621 6117 -1557
rect 6053 -1701 6117 -1637
rect 7228 -1461 7292 -1397
rect 7228 -1541 7292 -1477
rect 7228 -1621 7292 -1557
rect 6053 -1781 6117 -1717
rect 6389 -1663 6453 -1659
rect 6389 -1719 6393 -1663
rect 6393 -1719 6449 -1663
rect 6449 -1719 6453 -1663
rect 6389 -1723 6453 -1719
rect 6533 -1662 6597 -1658
rect 6533 -1718 6537 -1662
rect 6537 -1718 6593 -1662
rect 6593 -1718 6597 -1662
rect 6533 -1722 6597 -1718
rect 6664 -1663 6728 -1659
rect 6664 -1719 6668 -1663
rect 6668 -1719 6724 -1663
rect 6724 -1719 6728 -1663
rect 6664 -1723 6728 -1719
rect 7228 -1701 7292 -1637
rect 6053 -1861 6117 -1797
rect 6053 -1941 6117 -1877
rect 6053 -2021 6117 -1957
rect 6053 -2101 6117 -2037
rect 7228 -1781 7292 -1717
rect 7228 -1861 7292 -1797
rect 7228 -1941 7292 -1877
rect 7228 -2021 7292 -1957
rect 7228 -2101 7292 -2037
rect 7834 -1381 7898 -1317
rect 7834 -1461 7898 -1397
rect 7834 -1541 7898 -1477
rect 7834 -1621 7898 -1557
rect 7834 -1701 7898 -1637
rect 7834 -1781 7898 -1717
rect 7834 -1861 7898 -1797
rect 7834 -1941 7898 -1877
rect 7834 -2021 7898 -1957
rect 7834 -2101 7898 -2037
rect 8440 -1381 8504 -1317
rect 8440 -1461 8504 -1397
rect 8440 -1541 8504 -1477
rect 8440 -1621 8504 -1557
rect 8440 -1701 8504 -1637
rect 8440 -1781 8504 -1717
rect 8440 -1861 8504 -1797
rect 8440 -1941 8504 -1877
rect 8440 -2021 8504 -1957
rect 8440 -2101 8504 -2037
rect 9046 -1381 9110 -1317
rect 9046 -1461 9110 -1397
rect 9046 -1541 9110 -1477
rect 9046 -1621 9110 -1557
rect 9046 -1701 9110 -1637
rect 9046 -1781 9110 -1717
rect 9046 -1861 9110 -1797
rect 9046 -1941 9110 -1877
rect 9046 -2021 9110 -1957
rect 9046 -2101 9110 -2037
rect 9652 -1381 9716 -1317
rect 9652 -1461 9716 -1397
rect 9652 -1541 9716 -1477
rect 9652 -1621 9716 -1557
rect 9652 -1701 9716 -1637
rect 9652 -1781 9716 -1717
rect 9652 -1861 9716 -1797
rect 9652 -1941 9716 -1877
rect 9652 -2021 9716 -1957
rect 9652 -2101 9716 -2037
rect 10258 -1381 10322 -1317
rect 10258 -1461 10322 -1397
rect 10258 -1541 10322 -1477
rect 10258 -1621 10322 -1557
rect 10258 -1701 10322 -1637
rect 10258 -1781 10322 -1717
rect 10258 -1861 10322 -1797
rect 10258 -1941 10322 -1877
rect 10258 -2021 10322 -1957
rect 10258 -2101 10322 -2037
rect 10864 -1381 10928 -1317
rect 10864 -1461 10928 -1397
rect 10864 -1541 10928 -1477
rect 10864 -1621 10928 -1557
rect 10864 -1701 10928 -1637
rect 10864 -1781 10928 -1717
rect 10864 -1861 10928 -1797
rect 10864 -1941 10928 -1877
rect 10864 -2021 10928 -1957
rect 10864 -2101 10928 -2037
rect 11470 -1381 11534 -1317
rect 11470 -1461 11534 -1397
rect 11470 -1541 11534 -1477
rect 11470 -1621 11534 -1557
rect 11470 -1701 11534 -1637
rect 11470 -1781 11534 -1717
rect 11470 -1861 11534 -1797
rect 11470 -1941 11534 -1877
rect 11470 -2021 11534 -1957
rect 11470 -2101 11534 -2037
rect 12076 -1381 12140 -1317
rect 12076 -1461 12140 -1397
rect 12076 -1541 12140 -1477
rect 12076 -1621 12140 -1557
rect 12076 -1701 12140 -1637
rect 12076 -1781 12140 -1717
rect 12076 -1861 12140 -1797
rect 12076 -1941 12140 -1877
rect 12076 -2021 12140 -1957
rect 12076 -2101 12140 -2037
rect 12305 -1138 12316 -1097
rect 12316 -1138 12369 -1097
rect 12305 -1161 12369 -1138
rect 12385 -1161 12449 -1097
rect 12465 -1161 12529 -1097
rect 12545 -1161 12609 -1097
rect 12625 -1161 12689 -1097
rect 12705 -1161 12769 -1097
rect 12202 -1381 12266 -1317
rect 12202 -1461 12266 -1397
rect 12202 -1541 12266 -1477
rect 12202 -1621 12266 -1557
rect 12202 -1701 12266 -1637
rect 12202 -1781 12266 -1717
rect 12202 -1861 12266 -1797
rect 12202 -1941 12266 -1877
rect 12202 -2021 12266 -1957
rect 12202 -2101 12266 -2037
rect 13138 -1117 13202 -1113
rect 13138 -1173 13142 -1117
rect 13142 -1173 13198 -1117
rect 13198 -1173 13202 -1117
rect 13138 -1177 13202 -1173
rect 13281 -1117 13345 -1113
rect 13281 -1173 13285 -1117
rect 13285 -1173 13341 -1117
rect 13341 -1173 13345 -1117
rect 13281 -1177 13345 -1173
rect 13401 -1117 13465 -1113
rect 13401 -1173 13405 -1117
rect 13405 -1173 13461 -1117
rect 13461 -1173 13465 -1117
rect 13401 -1177 13465 -1173
rect 12808 -1381 12872 -1317
rect 12808 -1461 12872 -1397
rect 12808 -1541 12872 -1477
rect 12808 -1621 12872 -1557
rect 12808 -1701 12872 -1637
rect 12808 -1781 12872 -1717
rect 13144 -1663 13208 -1659
rect 13144 -1719 13148 -1663
rect 13148 -1719 13204 -1663
rect 13204 -1719 13208 -1663
rect 13144 -1723 13208 -1719
rect 13288 -1662 13352 -1658
rect 13288 -1718 13292 -1662
rect 13292 -1718 13348 -1662
rect 13348 -1718 13352 -1662
rect 13288 -1722 13352 -1718
rect 13419 -1663 13483 -1659
rect 13419 -1719 13423 -1663
rect 13423 -1719 13479 -1663
rect 13479 -1719 13483 -1663
rect 13419 -1723 13483 -1719
rect 12808 -1861 12872 -1797
rect 12808 -1941 12872 -1877
rect 12808 -2021 12872 -1957
rect 12808 -2101 12872 -2037
rect 576 -2321 640 -2257
rect 656 -2321 720 -2257
rect 736 -2321 800 -2257
rect 816 -2321 880 -2257
rect 896 -2321 960 -2257
rect 976 -2321 1040 -2257
rect 1182 -2321 1246 -2257
rect 1262 -2321 1326 -2257
rect 1342 -2321 1406 -2257
rect 1422 -2321 1486 -2257
rect 1502 -2321 1566 -2257
rect 1582 -2321 1646 -2257
rect 1788 -2321 1852 -2257
rect 1868 -2321 1932 -2257
rect 1948 -2321 2012 -2257
rect 2028 -2321 2092 -2257
rect 2108 -2321 2172 -2257
rect 2188 -2321 2252 -2257
rect 2394 -2321 2458 -2257
rect 2474 -2321 2538 -2257
rect 2554 -2321 2618 -2257
rect 2634 -2321 2698 -2257
rect 2714 -2321 2778 -2257
rect 2794 -2321 2858 -2257
rect 3000 -2321 3064 -2257
rect 3080 -2321 3144 -2257
rect 3160 -2321 3224 -2257
rect 3240 -2321 3304 -2257
rect 3320 -2321 3384 -2257
rect 3400 -2321 3464 -2257
rect 3606 -2321 3670 -2257
rect 3686 -2321 3750 -2257
rect 3766 -2321 3830 -2257
rect 3846 -2321 3910 -2257
rect 3926 -2321 3990 -2257
rect 4006 -2321 4070 -2257
rect 4212 -2321 4276 -2257
rect 4292 -2321 4356 -2257
rect 4372 -2321 4436 -2257
rect 4452 -2321 4516 -2257
rect 4532 -2321 4596 -2257
rect 4612 -2321 4676 -2257
rect 4818 -2321 4882 -2257
rect 4898 -2321 4962 -2257
rect 4978 -2321 5042 -2257
rect 5058 -2321 5122 -2257
rect 5138 -2321 5202 -2257
rect 5218 -2321 5282 -2257
rect 5550 -2321 5614 -2257
rect 5630 -2321 5694 -2257
rect 5710 -2321 5774 -2257
rect 5790 -2321 5854 -2257
rect 5870 -2321 5934 -2257
rect 5950 -2321 6014 -2257
rect 6047 -2268 6111 -2264
rect 6047 -2324 6051 -2268
rect 6051 -2324 6107 -2268
rect 6107 -2324 6111 -2268
rect 6047 -2328 6111 -2324
rect 7331 -2321 7395 -2257
rect 7411 -2321 7475 -2257
rect 7491 -2321 7555 -2257
rect 7571 -2321 7635 -2257
rect 7651 -2321 7715 -2257
rect 7731 -2321 7795 -2257
rect 7937 -2321 8001 -2257
rect 8017 -2321 8081 -2257
rect 8097 -2321 8161 -2257
rect 8177 -2321 8241 -2257
rect 8257 -2321 8321 -2257
rect 8337 -2321 8401 -2257
rect 8543 -2321 8607 -2257
rect 8623 -2321 8687 -2257
rect 8703 -2321 8767 -2257
rect 8783 -2321 8847 -2257
rect 8863 -2321 8927 -2257
rect 8943 -2321 9007 -2257
rect 9149 -2321 9213 -2257
rect 9229 -2321 9293 -2257
rect 9309 -2321 9373 -2257
rect 9389 -2321 9453 -2257
rect 9469 -2321 9533 -2257
rect 9549 -2321 9613 -2257
rect 9755 -2321 9819 -2257
rect 9835 -2321 9899 -2257
rect 9915 -2321 9979 -2257
rect 9995 -2321 10059 -2257
rect 10075 -2321 10139 -2257
rect 10155 -2321 10219 -2257
rect 10361 -2321 10425 -2257
rect 10441 -2321 10505 -2257
rect 10521 -2321 10585 -2257
rect 10601 -2321 10665 -2257
rect 10681 -2321 10745 -2257
rect 10761 -2321 10825 -2257
rect 10967 -2321 11031 -2257
rect 11047 -2321 11111 -2257
rect 11127 -2321 11191 -2257
rect 11207 -2321 11271 -2257
rect 11287 -2321 11351 -2257
rect 11367 -2321 11431 -2257
rect 11573 -2321 11637 -2257
rect 11653 -2321 11717 -2257
rect 11733 -2321 11797 -2257
rect 11813 -2321 11877 -2257
rect 11893 -2321 11957 -2257
rect 11973 -2321 12037 -2257
rect 12305 -2321 12369 -2257
rect 12385 -2321 12449 -2257
rect 12465 -2321 12529 -2257
rect 12545 -2321 12609 -2257
rect 12625 -2321 12689 -2257
rect 12705 -2321 12769 -2257
rect 12802 -2268 12866 -2264
rect 12802 -2324 12806 -2268
rect 12806 -2324 12862 -2268
rect 12862 -2324 12866 -2268
rect 12802 -2328 12866 -2324
<< metal4 >>
rect 707 3281 833 3286
rect 7396 3281 7522 3286
rect 61 3276 13444 3281
rect 61 3212 738 3276
rect 802 3269 7427 3276
rect 802 3212 835 3269
rect 61 3205 835 3212
rect 899 3205 915 3269
rect 979 3205 995 3269
rect 1059 3205 1075 3269
rect 1139 3205 1155 3269
rect 1219 3205 1235 3269
rect 1299 3205 1567 3269
rect 1631 3205 1647 3269
rect 1711 3205 1727 3269
rect 1791 3205 1807 3269
rect 1871 3205 1887 3269
rect 1951 3205 1967 3269
rect 2031 3205 2173 3269
rect 2237 3205 2253 3269
rect 2317 3205 2333 3269
rect 2397 3205 2413 3269
rect 2477 3205 2493 3269
rect 2557 3205 2573 3269
rect 2637 3205 2779 3269
rect 2843 3205 2859 3269
rect 2923 3205 2939 3269
rect 3003 3205 3019 3269
rect 3083 3205 3099 3269
rect 3163 3205 3179 3269
rect 3243 3205 3385 3269
rect 3449 3205 3465 3269
rect 3529 3205 3545 3269
rect 3609 3205 3625 3269
rect 3689 3205 3705 3269
rect 3769 3205 3785 3269
rect 3849 3205 3991 3269
rect 4055 3205 4071 3269
rect 4135 3205 4151 3269
rect 4215 3205 4231 3269
rect 4295 3205 4311 3269
rect 4375 3205 4391 3269
rect 4455 3205 4597 3269
rect 4661 3205 4677 3269
rect 4741 3205 4757 3269
rect 4821 3205 4837 3269
rect 4901 3205 4917 3269
rect 4981 3205 4997 3269
rect 5061 3205 5203 3269
rect 5267 3205 5283 3269
rect 5347 3205 5363 3269
rect 5427 3205 5443 3269
rect 5507 3205 5523 3269
rect 5587 3205 5603 3269
rect 5667 3205 5809 3269
rect 5873 3205 5889 3269
rect 5953 3205 5969 3269
rect 6033 3205 6049 3269
rect 6113 3205 6129 3269
rect 6193 3205 6209 3269
rect 6273 3212 7427 3269
rect 7491 3269 13444 3276
rect 7491 3212 7524 3269
rect 6273 3205 7524 3212
rect 7588 3205 7604 3269
rect 7668 3205 7684 3269
rect 7748 3205 7764 3269
rect 7828 3205 7844 3269
rect 7908 3205 7924 3269
rect 7988 3205 8256 3269
rect 8320 3205 8336 3269
rect 8400 3205 8416 3269
rect 8480 3205 8496 3269
rect 8560 3205 8576 3269
rect 8640 3205 8656 3269
rect 8720 3205 8862 3269
rect 8926 3205 8942 3269
rect 9006 3205 9022 3269
rect 9086 3205 9102 3269
rect 9166 3205 9182 3269
rect 9246 3205 9262 3269
rect 9326 3205 9468 3269
rect 9532 3205 9548 3269
rect 9612 3205 9628 3269
rect 9692 3205 9708 3269
rect 9772 3205 9788 3269
rect 9852 3205 9868 3269
rect 9932 3205 10074 3269
rect 10138 3205 10154 3269
rect 10218 3205 10234 3269
rect 10298 3205 10314 3269
rect 10378 3205 10394 3269
rect 10458 3205 10474 3269
rect 10538 3205 10680 3269
rect 10744 3205 10760 3269
rect 10824 3205 10840 3269
rect 10904 3205 10920 3269
rect 10984 3205 11000 3269
rect 11064 3205 11080 3269
rect 11144 3205 11286 3269
rect 11350 3205 11366 3269
rect 11430 3205 11446 3269
rect 11510 3205 11526 3269
rect 11590 3205 11606 3269
rect 11670 3205 11686 3269
rect 11750 3205 11892 3269
rect 11956 3205 11972 3269
rect 12036 3205 12052 3269
rect 12116 3205 12132 3269
rect 12196 3205 12212 3269
rect 12276 3205 12292 3269
rect 12356 3205 12498 3269
rect 12562 3205 12578 3269
rect 12642 3205 12658 3269
rect 12722 3205 12738 3269
rect 12802 3205 12818 3269
rect 12882 3205 12898 3269
rect 12962 3205 13444 3269
rect 61 3203 13444 3205
rect 61 2671 523 3203
rect 61 2607 121 2671
rect 185 2670 396 2671
rect 185 2607 252 2670
rect 61 2606 252 2607
rect 316 2607 396 2670
rect 460 2607 523 2671
rect 316 2606 523 2607
rect 61 2588 523 2606
rect 731 3049 797 3139
rect 731 2985 732 3049
rect 796 2985 797 3049
rect 731 2969 797 2985
rect 731 2905 732 2969
rect 796 2905 797 2969
rect 731 2889 797 2905
rect 731 2825 732 2889
rect 796 2825 797 2889
rect 731 2809 797 2825
rect 731 2745 732 2809
rect 796 2745 797 2809
rect 731 2729 797 2745
rect 731 2665 732 2729
rect 796 2665 797 2729
rect 731 2649 797 2665
rect 731 2585 732 2649
rect 796 2585 797 2649
rect 731 2569 797 2585
rect 731 2505 732 2569
rect 796 2505 797 2569
rect 731 2489 797 2505
rect 731 2425 732 2489
rect 796 2425 797 2489
rect 731 2409 797 2425
rect 731 2345 732 2409
rect 796 2345 797 2409
rect 731 2329 797 2345
rect 731 2265 732 2329
rect 796 2265 797 2329
rect 78 2125 509 2140
rect 78 2061 139 2125
rect 203 2061 259 2125
rect 323 2061 402 2125
rect 466 2061 509 2125
rect 78 2046 509 2061
rect 79 702 509 2046
rect 731 2111 797 2265
rect 857 2173 917 3203
rect 977 2111 1037 3143
rect 1097 2173 1157 3203
rect 1217 2111 1277 3143
rect 1337 3049 1403 3139
rect 1337 2985 1338 3049
rect 1402 2985 1403 3049
rect 1337 2969 1403 2985
rect 1337 2905 1338 2969
rect 1402 2905 1403 2969
rect 1337 2889 1403 2905
rect 1337 2825 1338 2889
rect 1402 2825 1403 2889
rect 1337 2809 1403 2825
rect 1337 2745 1338 2809
rect 1402 2745 1403 2809
rect 1337 2729 1403 2745
rect 1337 2665 1338 2729
rect 1402 2665 1403 2729
rect 1337 2649 1403 2665
rect 1337 2585 1338 2649
rect 1402 2585 1403 2649
rect 1337 2569 1403 2585
rect 1337 2505 1338 2569
rect 1402 2505 1403 2569
rect 1337 2489 1403 2505
rect 1337 2425 1338 2489
rect 1402 2425 1403 2489
rect 1337 2409 1403 2425
rect 1337 2345 1338 2409
rect 1402 2345 1403 2409
rect 1337 2329 1403 2345
rect 1337 2265 1338 2329
rect 1402 2265 1403 2329
rect 1337 2111 1403 2265
rect 731 2109 1403 2111
rect 731 2045 835 2109
rect 899 2045 915 2109
rect 979 2045 995 2109
rect 1059 2045 1075 2109
rect 1139 2045 1155 2109
rect 1219 2045 1235 2109
rect 1299 2045 1403 2109
rect 731 2043 1403 2045
rect 1463 3049 1529 3139
rect 1463 2985 1464 3049
rect 1528 2985 1529 3049
rect 1463 2969 1529 2985
rect 1463 2905 1464 2969
rect 1528 2905 1529 2969
rect 1463 2889 1529 2905
rect 1463 2825 1464 2889
rect 1528 2825 1529 2889
rect 1463 2809 1529 2825
rect 1463 2745 1464 2809
rect 1528 2745 1529 2809
rect 1463 2729 1529 2745
rect 1463 2665 1464 2729
rect 1528 2665 1529 2729
rect 1463 2649 1529 2665
rect 1463 2585 1464 2649
rect 1528 2585 1529 2649
rect 1463 2569 1529 2585
rect 1463 2505 1464 2569
rect 1528 2505 1529 2569
rect 1463 2489 1529 2505
rect 1463 2425 1464 2489
rect 1528 2425 1529 2489
rect 1463 2409 1529 2425
rect 1463 2345 1464 2409
rect 1528 2345 1529 2409
rect 1463 2329 1529 2345
rect 1463 2265 1464 2329
rect 1528 2265 1529 2329
rect 1463 2111 1529 2265
rect 1589 2173 1649 3203
rect 1709 2111 1769 3143
rect 1829 2173 1889 3203
rect 1949 2111 2009 3143
rect 2069 3049 2135 3139
rect 2069 2985 2070 3049
rect 2134 2985 2135 3049
rect 2069 2969 2135 2985
rect 2069 2905 2070 2969
rect 2134 2905 2135 2969
rect 2069 2889 2135 2905
rect 2069 2825 2070 2889
rect 2134 2825 2135 2889
rect 2069 2809 2135 2825
rect 2069 2745 2070 2809
rect 2134 2745 2135 2809
rect 2069 2729 2135 2745
rect 2069 2665 2070 2729
rect 2134 2665 2135 2729
rect 2069 2649 2135 2665
rect 2069 2585 2070 2649
rect 2134 2585 2135 2649
rect 2069 2569 2135 2585
rect 2069 2505 2070 2569
rect 2134 2505 2135 2569
rect 2069 2489 2135 2505
rect 2069 2425 2070 2489
rect 2134 2425 2135 2489
rect 2069 2409 2135 2425
rect 2069 2345 2070 2409
rect 2134 2345 2135 2409
rect 2069 2329 2135 2345
rect 2069 2265 2070 2329
rect 2134 2265 2135 2329
rect 2069 2111 2135 2265
rect 2195 2111 2255 3143
rect 2315 2173 2375 3203
rect 2435 2111 2495 3143
rect 2555 2173 2615 3203
rect 2675 3049 2741 3139
rect 2675 2985 2676 3049
rect 2740 2985 2741 3049
rect 2675 2969 2741 2985
rect 2675 2905 2676 2969
rect 2740 2905 2741 2969
rect 2675 2889 2741 2905
rect 2675 2825 2676 2889
rect 2740 2825 2741 2889
rect 2675 2809 2741 2825
rect 2675 2745 2676 2809
rect 2740 2745 2741 2809
rect 2675 2729 2741 2745
rect 2675 2665 2676 2729
rect 2740 2665 2741 2729
rect 2675 2649 2741 2665
rect 2675 2585 2676 2649
rect 2740 2585 2741 2649
rect 2675 2569 2741 2585
rect 2675 2505 2676 2569
rect 2740 2505 2741 2569
rect 2675 2489 2741 2505
rect 2675 2425 2676 2489
rect 2740 2425 2741 2489
rect 2675 2409 2741 2425
rect 2675 2345 2676 2409
rect 2740 2345 2741 2409
rect 2675 2329 2741 2345
rect 2675 2265 2676 2329
rect 2740 2265 2741 2329
rect 2675 2111 2741 2265
rect 2801 2173 2861 3203
rect 2921 2111 2981 3143
rect 3041 2173 3101 3203
rect 3161 2111 3221 3143
rect 3281 3049 3347 3139
rect 3281 2985 3282 3049
rect 3346 2985 3347 3049
rect 3281 2969 3347 2985
rect 3281 2905 3282 2969
rect 3346 2905 3347 2969
rect 3281 2889 3347 2905
rect 3281 2825 3282 2889
rect 3346 2825 3347 2889
rect 3281 2809 3347 2825
rect 3281 2745 3282 2809
rect 3346 2745 3347 2809
rect 3281 2729 3347 2745
rect 3281 2665 3282 2729
rect 3346 2665 3347 2729
rect 3281 2649 3347 2665
rect 3281 2585 3282 2649
rect 3346 2585 3347 2649
rect 3281 2569 3347 2585
rect 3281 2505 3282 2569
rect 3346 2505 3347 2569
rect 3281 2489 3347 2505
rect 3281 2425 3282 2489
rect 3346 2425 3347 2489
rect 3281 2409 3347 2425
rect 3281 2345 3282 2409
rect 3346 2345 3347 2409
rect 3281 2329 3347 2345
rect 3281 2265 3282 2329
rect 3346 2265 3347 2329
rect 3281 2111 3347 2265
rect 3407 2111 3467 3143
rect 3527 2173 3587 3203
rect 3647 2111 3707 3143
rect 3767 2173 3827 3203
rect 3887 3049 3953 3139
rect 3887 2985 3888 3049
rect 3952 2985 3953 3049
rect 3887 2969 3953 2985
rect 3887 2905 3888 2969
rect 3952 2905 3953 2969
rect 3887 2889 3953 2905
rect 3887 2825 3888 2889
rect 3952 2825 3953 2889
rect 3887 2809 3953 2825
rect 3887 2745 3888 2809
rect 3952 2745 3953 2809
rect 3887 2729 3953 2745
rect 3887 2665 3888 2729
rect 3952 2665 3953 2729
rect 3887 2649 3953 2665
rect 3887 2585 3888 2649
rect 3952 2585 3953 2649
rect 3887 2569 3953 2585
rect 3887 2505 3888 2569
rect 3952 2505 3953 2569
rect 3887 2489 3953 2505
rect 3887 2425 3888 2489
rect 3952 2425 3953 2489
rect 3887 2409 3953 2425
rect 3887 2345 3888 2409
rect 3952 2345 3953 2409
rect 3887 2329 3953 2345
rect 3887 2265 3888 2329
rect 3952 2265 3953 2329
rect 3887 2111 3953 2265
rect 4013 2173 4073 3203
rect 4133 2111 4193 3143
rect 4253 2173 4313 3203
rect 4373 2111 4433 3143
rect 4493 3049 4559 3139
rect 4493 2985 4494 3049
rect 4558 2985 4559 3049
rect 4493 2969 4559 2985
rect 4493 2905 4494 2969
rect 4558 2905 4559 2969
rect 4493 2889 4559 2905
rect 4493 2825 4494 2889
rect 4558 2825 4559 2889
rect 4493 2809 4559 2825
rect 4493 2745 4494 2809
rect 4558 2745 4559 2809
rect 4493 2729 4559 2745
rect 4493 2665 4494 2729
rect 4558 2665 4559 2729
rect 4493 2649 4559 2665
rect 4493 2585 4494 2649
rect 4558 2585 4559 2649
rect 4493 2569 4559 2585
rect 4493 2505 4494 2569
rect 4558 2505 4559 2569
rect 4493 2489 4559 2505
rect 4493 2425 4494 2489
rect 4558 2425 4559 2489
rect 4493 2409 4559 2425
rect 4493 2345 4494 2409
rect 4558 2345 4559 2409
rect 4493 2329 4559 2345
rect 4493 2265 4494 2329
rect 4558 2265 4559 2329
rect 4493 2111 4559 2265
rect 4619 2111 4679 3143
rect 4739 2173 4799 3203
rect 4859 2111 4919 3143
rect 4979 2173 5039 3203
rect 5099 3049 5165 3139
rect 5099 2985 5100 3049
rect 5164 2985 5165 3049
rect 5099 2969 5165 2985
rect 5099 2905 5100 2969
rect 5164 2905 5165 2969
rect 5099 2889 5165 2905
rect 5099 2825 5100 2889
rect 5164 2825 5165 2889
rect 5099 2809 5165 2825
rect 5099 2745 5100 2809
rect 5164 2745 5165 2809
rect 5099 2729 5165 2745
rect 5099 2665 5100 2729
rect 5164 2665 5165 2729
rect 5099 2649 5165 2665
rect 5099 2585 5100 2649
rect 5164 2585 5165 2649
rect 5099 2569 5165 2585
rect 5099 2505 5100 2569
rect 5164 2505 5165 2569
rect 5099 2489 5165 2505
rect 5099 2425 5100 2489
rect 5164 2425 5165 2489
rect 5099 2409 5165 2425
rect 5099 2345 5100 2409
rect 5164 2345 5165 2409
rect 5099 2329 5165 2345
rect 5099 2265 5100 2329
rect 5164 2265 5165 2329
rect 5099 2111 5165 2265
rect 5225 2173 5285 3203
rect 5345 2111 5405 3143
rect 5465 2173 5525 3203
rect 5585 2111 5645 3143
rect 5705 3049 5771 3139
rect 5705 2985 5706 3049
rect 5770 2985 5771 3049
rect 5705 2969 5771 2985
rect 5705 2905 5706 2969
rect 5770 2905 5771 2969
rect 5705 2889 5771 2905
rect 5705 2825 5706 2889
rect 5770 2825 5771 2889
rect 5705 2809 5771 2825
rect 5705 2745 5706 2809
rect 5770 2745 5771 2809
rect 5705 2729 5771 2745
rect 5705 2665 5706 2729
rect 5770 2665 5771 2729
rect 5705 2649 5771 2665
rect 5705 2585 5706 2649
rect 5770 2585 5771 2649
rect 5705 2569 5771 2585
rect 5705 2505 5706 2569
rect 5770 2505 5771 2569
rect 5705 2489 5771 2505
rect 5705 2425 5706 2489
rect 5770 2425 5771 2489
rect 5705 2409 5771 2425
rect 5705 2345 5706 2409
rect 5770 2345 5771 2409
rect 5705 2329 5771 2345
rect 5705 2265 5706 2329
rect 5770 2265 5771 2329
rect 5705 2111 5771 2265
rect 5831 2111 5891 3143
rect 5951 2173 6011 3203
rect 6071 2111 6131 3143
rect 6191 2173 6251 3203
rect 6311 3049 6377 3139
rect 6311 2985 6312 3049
rect 6376 2985 6377 3049
rect 6311 2969 6377 2985
rect 6311 2905 6312 2969
rect 6376 2905 6377 2969
rect 6311 2889 6377 2905
rect 6311 2825 6312 2889
rect 6376 2825 6377 2889
rect 6311 2809 6377 2825
rect 6311 2745 6312 2809
rect 6376 2745 6377 2809
rect 6311 2729 6377 2745
rect 6311 2665 6312 2729
rect 6376 2665 6377 2729
rect 6311 2649 6377 2665
rect 6311 2585 6312 2649
rect 6376 2585 6377 2649
rect 6311 2569 6377 2585
rect 6311 2505 6312 2569
rect 6376 2505 6377 2569
rect 6311 2489 6377 2505
rect 6311 2425 6312 2489
rect 6376 2425 6377 2489
rect 6311 2409 6377 2425
rect 6311 2345 6312 2409
rect 6376 2345 6377 2409
rect 6311 2329 6377 2345
rect 6311 2265 6312 2329
rect 6376 2265 6377 2329
rect 6437 2671 7212 3203
rect 6437 2607 6810 2671
rect 6874 2670 7085 2671
rect 6874 2607 6941 2670
rect 6437 2606 6941 2607
rect 7005 2607 7085 2670
rect 7149 2607 7212 2671
rect 7005 2606 7212 2607
rect 6437 2588 7212 2606
rect 7420 3049 7486 3139
rect 7420 2985 7421 3049
rect 7485 2985 7486 3049
rect 7420 2969 7486 2985
rect 7420 2905 7421 2969
rect 7485 2905 7486 2969
rect 7420 2889 7486 2905
rect 7420 2825 7421 2889
rect 7485 2825 7486 2889
rect 7420 2809 7486 2825
rect 7420 2745 7421 2809
rect 7485 2745 7486 2809
rect 7420 2729 7486 2745
rect 7420 2665 7421 2729
rect 7485 2665 7486 2729
rect 7420 2649 7486 2665
rect 6437 2349 6866 2588
rect 6437 2285 6470 2349
rect 6534 2285 6866 2349
rect 6437 2273 6866 2285
rect 6311 2111 6377 2265
rect 1463 2109 6377 2111
rect 1463 2045 1567 2109
rect 1631 2045 1647 2109
rect 1711 2045 1727 2109
rect 1791 2045 1807 2109
rect 1871 2045 1887 2109
rect 1951 2045 1967 2109
rect 2031 2045 2173 2109
rect 2237 2045 2253 2109
rect 2317 2045 2333 2109
rect 2397 2045 2413 2109
rect 2477 2045 2493 2109
rect 2557 2045 2573 2109
rect 2637 2045 2779 2109
rect 2843 2045 2859 2109
rect 2923 2045 2939 2109
rect 3003 2045 3019 2109
rect 3083 2045 3099 2109
rect 3163 2045 3179 2109
rect 3243 2045 3385 2109
rect 3449 2045 3465 2109
rect 3529 2045 3545 2109
rect 3609 2045 3625 2109
rect 3689 2045 3705 2109
rect 3769 2045 3785 2109
rect 3849 2045 3991 2109
rect 4055 2045 4071 2109
rect 4135 2045 4151 2109
rect 4215 2045 4231 2109
rect 4295 2045 4311 2109
rect 4375 2045 4391 2109
rect 4455 2045 4597 2109
rect 4661 2045 4677 2109
rect 4741 2045 4757 2109
rect 4821 2045 4837 2109
rect 4901 2045 4917 2109
rect 4981 2045 4997 2109
rect 5061 2045 5203 2109
rect 5267 2045 5283 2109
rect 5347 2045 5363 2109
rect 5427 2045 5443 2109
rect 5507 2045 5523 2109
rect 5587 2045 5603 2109
rect 5667 2045 5809 2109
rect 5873 2045 5889 2109
rect 5953 2045 5969 2109
rect 6033 2045 6049 2109
rect 6113 2045 6129 2109
rect 6193 2045 6209 2109
rect 6273 2045 6377 2109
rect 6638 2140 6866 2273
rect 7420 2585 7421 2649
rect 7485 2585 7486 2649
rect 7420 2569 7486 2585
rect 7420 2505 7421 2569
rect 7485 2505 7486 2569
rect 7420 2489 7486 2505
rect 7420 2425 7421 2489
rect 7485 2425 7486 2489
rect 7420 2409 7486 2425
rect 7420 2345 7421 2409
rect 7485 2345 7486 2409
rect 7420 2329 7486 2345
rect 7420 2265 7421 2329
rect 7485 2265 7486 2329
rect 6638 2125 7198 2140
rect 1463 2043 6377 2045
rect 6437 2088 6635 2098
rect 6437 2024 6558 2088
rect 6622 2024 6635 2088
rect 6437 2014 6635 2024
rect 6638 2061 6828 2125
rect 6892 2061 6948 2125
rect 7012 2061 7091 2125
rect 7155 2061 7198 2125
rect 1085 1860 1757 1862
rect 1085 1796 1189 1860
rect 1253 1796 1269 1860
rect 1333 1796 1349 1860
rect 1413 1796 1429 1860
rect 1493 1796 1509 1860
rect 1573 1796 1589 1860
rect 1653 1796 1757 1860
rect 1085 1794 1757 1796
rect 1085 1640 1151 1794
rect 1085 1576 1086 1640
rect 1150 1576 1151 1640
rect 1085 1560 1151 1576
rect 1085 1496 1086 1560
rect 1150 1496 1151 1560
rect 1085 1480 1151 1496
rect 1085 1416 1086 1480
rect 1150 1416 1151 1480
rect 1085 1400 1151 1416
rect 1085 1336 1086 1400
rect 1150 1336 1151 1400
rect 1085 1320 1151 1336
rect 1085 1256 1086 1320
rect 1150 1256 1151 1320
rect 1085 1240 1151 1256
rect 1085 1176 1086 1240
rect 1150 1176 1151 1240
rect 1085 1160 1151 1176
rect 1085 1096 1086 1160
rect 1150 1096 1151 1160
rect 1085 1080 1151 1096
rect 1085 1016 1086 1080
rect 1150 1016 1151 1080
rect 1085 1000 1151 1016
rect 1085 936 1086 1000
rect 1150 936 1151 1000
rect 1085 920 1151 936
rect 1085 856 1086 920
rect 1150 856 1151 920
rect 1085 766 1151 856
rect 694 702 819 708
rect 1211 702 1271 1732
rect 1331 762 1391 1794
rect 1451 702 1511 1732
rect 1571 762 1631 1794
rect 1691 1640 1757 1794
rect 1691 1576 1692 1640
rect 1756 1576 1757 1640
rect 1691 1560 1757 1576
rect 1691 1496 1692 1560
rect 1756 1496 1757 1560
rect 1691 1480 1757 1496
rect 1691 1416 1692 1480
rect 1756 1416 1757 1480
rect 1691 1400 1757 1416
rect 1691 1336 1692 1400
rect 1756 1336 1757 1400
rect 1691 1320 1757 1336
rect 1691 1256 1692 1320
rect 1756 1256 1757 1320
rect 1691 1240 1757 1256
rect 1691 1176 1692 1240
rect 1756 1176 1757 1240
rect 1691 1160 1757 1176
rect 1691 1096 1692 1160
rect 1756 1096 1757 1160
rect 1691 1080 1757 1096
rect 1691 1016 1692 1080
rect 1756 1016 1757 1080
rect 1691 1000 1757 1016
rect 1691 936 1692 1000
rect 1756 936 1757 1000
rect 1691 920 1757 936
rect 1691 856 1692 920
rect 1756 856 1757 920
rect 1691 766 1757 856
rect 1817 1860 4307 1862
rect 1817 1796 1921 1860
rect 1985 1796 2001 1860
rect 2065 1796 2081 1860
rect 2145 1796 2161 1860
rect 2225 1796 2241 1860
rect 2305 1796 2321 1860
rect 2385 1796 2527 1860
rect 2591 1796 2607 1860
rect 2671 1796 2687 1860
rect 2751 1796 2767 1860
rect 2831 1796 2847 1860
rect 2911 1796 2927 1860
rect 2991 1796 3133 1860
rect 3197 1796 3213 1860
rect 3277 1796 3293 1860
rect 3357 1796 3373 1860
rect 3437 1796 3453 1860
rect 3517 1796 3533 1860
rect 3597 1796 3739 1860
rect 3803 1796 3819 1860
rect 3883 1796 3899 1860
rect 3963 1796 3979 1860
rect 4043 1796 4059 1860
rect 4123 1796 4139 1860
rect 4203 1796 4307 1860
rect 1817 1794 4307 1796
rect 1817 1640 1883 1794
rect 1817 1576 1818 1640
rect 1882 1576 1883 1640
rect 1817 1560 1883 1576
rect 1817 1496 1818 1560
rect 1882 1496 1883 1560
rect 1817 1480 1883 1496
rect 1817 1416 1818 1480
rect 1882 1416 1883 1480
rect 1817 1400 1883 1416
rect 1817 1336 1818 1400
rect 1882 1336 1883 1400
rect 1817 1320 1883 1336
rect 1817 1256 1818 1320
rect 1882 1256 1883 1320
rect 1817 1240 1883 1256
rect 1817 1176 1818 1240
rect 1882 1176 1883 1240
rect 1817 1160 1883 1176
rect 1817 1096 1818 1160
rect 1882 1096 1883 1160
rect 1817 1080 1883 1096
rect 1817 1016 1818 1080
rect 1882 1016 1883 1080
rect 1817 1000 1883 1016
rect 1817 936 1818 1000
rect 1882 936 1883 1000
rect 1817 920 1883 936
rect 1817 856 1818 920
rect 1882 856 1883 920
rect 1817 766 1883 856
rect 1943 702 2003 1732
rect 2063 762 2123 1794
rect 2183 702 2243 1732
rect 2303 762 2363 1794
rect 2423 1640 2489 1794
rect 2423 1576 2424 1640
rect 2488 1576 2489 1640
rect 2423 1560 2489 1576
rect 2423 1496 2424 1560
rect 2488 1496 2489 1560
rect 2423 1480 2489 1496
rect 2423 1416 2424 1480
rect 2488 1416 2489 1480
rect 2423 1400 2489 1416
rect 2423 1336 2424 1400
rect 2488 1336 2489 1400
rect 2423 1320 2489 1336
rect 2423 1256 2424 1320
rect 2488 1256 2489 1320
rect 2423 1240 2489 1256
rect 2423 1176 2424 1240
rect 2488 1176 2489 1240
rect 2423 1160 2489 1176
rect 2423 1096 2424 1160
rect 2488 1096 2489 1160
rect 2423 1080 2489 1096
rect 2423 1016 2424 1080
rect 2488 1016 2489 1080
rect 2423 1000 2489 1016
rect 2423 936 2424 1000
rect 2488 936 2489 1000
rect 2423 920 2489 936
rect 2423 856 2424 920
rect 2488 856 2489 920
rect 2423 766 2489 856
rect 2549 762 2609 1794
rect 2669 702 2729 1732
rect 2789 762 2849 1794
rect 2909 702 2969 1732
rect 3029 1640 3095 1794
rect 3029 1576 3030 1640
rect 3094 1576 3095 1640
rect 3029 1560 3095 1576
rect 3029 1496 3030 1560
rect 3094 1496 3095 1560
rect 3029 1480 3095 1496
rect 3029 1416 3030 1480
rect 3094 1416 3095 1480
rect 3029 1400 3095 1416
rect 3029 1336 3030 1400
rect 3094 1336 3095 1400
rect 3029 1320 3095 1336
rect 3029 1256 3030 1320
rect 3094 1256 3095 1320
rect 3029 1240 3095 1256
rect 3029 1176 3030 1240
rect 3094 1176 3095 1240
rect 3029 1160 3095 1176
rect 3029 1096 3030 1160
rect 3094 1096 3095 1160
rect 3029 1080 3095 1096
rect 3029 1016 3030 1080
rect 3094 1016 3095 1080
rect 3029 1000 3095 1016
rect 3029 936 3030 1000
rect 3094 936 3095 1000
rect 3029 920 3095 936
rect 3029 856 3030 920
rect 3094 856 3095 920
rect 3029 766 3095 856
rect 3155 702 3215 1732
rect 3275 762 3335 1794
rect 3395 702 3455 1732
rect 3515 762 3575 1794
rect 3635 1640 3701 1794
rect 3635 1576 3636 1640
rect 3700 1576 3701 1640
rect 3635 1560 3701 1576
rect 3635 1496 3636 1560
rect 3700 1496 3701 1560
rect 3635 1480 3701 1496
rect 3635 1416 3636 1480
rect 3700 1416 3701 1480
rect 3635 1400 3701 1416
rect 3635 1336 3636 1400
rect 3700 1336 3701 1400
rect 3635 1320 3701 1336
rect 3635 1256 3636 1320
rect 3700 1256 3701 1320
rect 3635 1240 3701 1256
rect 3635 1176 3636 1240
rect 3700 1176 3701 1240
rect 3635 1160 3701 1176
rect 3635 1096 3636 1160
rect 3700 1096 3701 1160
rect 3635 1080 3701 1096
rect 3635 1016 3636 1080
rect 3700 1016 3701 1080
rect 3635 1000 3701 1016
rect 3635 936 3636 1000
rect 3700 936 3701 1000
rect 3635 920 3701 936
rect 3635 856 3636 920
rect 3700 856 3701 920
rect 3635 766 3701 856
rect 3761 762 3821 1794
rect 3881 702 3941 1732
rect 4001 762 4061 1794
rect 4121 702 4181 1732
rect 4241 1640 4307 1794
rect 4241 1576 4242 1640
rect 4306 1576 4307 1640
rect 4241 1560 4307 1576
rect 4241 1496 4242 1560
rect 4306 1496 4307 1560
rect 4241 1480 4307 1496
rect 4241 1416 4242 1480
rect 4306 1416 4307 1480
rect 4241 1400 4307 1416
rect 4241 1336 4242 1400
rect 4306 1336 4307 1400
rect 4241 1320 4307 1336
rect 4241 1256 4242 1320
rect 4306 1256 4307 1320
rect 4241 1240 4307 1256
rect 4241 1176 4242 1240
rect 4306 1176 4307 1240
rect 4241 1160 4307 1176
rect 4241 1096 4242 1160
rect 4306 1096 4307 1160
rect 4241 1080 4307 1096
rect 4241 1016 4242 1080
rect 4306 1016 4307 1080
rect 4241 1000 4307 1016
rect 4241 936 4242 1000
rect 4306 936 4307 1000
rect 4241 920 4307 936
rect 4241 856 4242 920
rect 4306 856 4307 920
rect 4241 766 4307 856
rect 4367 1860 5645 1862
rect 4367 1796 4471 1860
rect 4535 1796 4551 1860
rect 4615 1796 4631 1860
rect 4695 1796 4711 1860
rect 4775 1796 4791 1860
rect 4855 1796 4871 1860
rect 4935 1796 5077 1860
rect 5141 1796 5157 1860
rect 5221 1796 5237 1860
rect 5301 1796 5317 1860
rect 5381 1796 5397 1860
rect 5461 1796 5477 1860
rect 5541 1796 5645 1860
rect 4367 1794 5645 1796
rect 4367 1640 4433 1794
rect 4367 1576 4368 1640
rect 4432 1576 4433 1640
rect 4367 1560 4433 1576
rect 4367 1496 4368 1560
rect 4432 1496 4433 1560
rect 4367 1480 4433 1496
rect 4367 1416 4368 1480
rect 4432 1416 4433 1480
rect 4367 1400 4433 1416
rect 4367 1336 4368 1400
rect 4432 1336 4433 1400
rect 4367 1320 4433 1336
rect 4367 1256 4368 1320
rect 4432 1256 4433 1320
rect 4367 1240 4433 1256
rect 4367 1176 4368 1240
rect 4432 1176 4433 1240
rect 4367 1160 4433 1176
rect 4367 1096 4368 1160
rect 4432 1096 4433 1160
rect 4367 1080 4433 1096
rect 4367 1016 4368 1080
rect 4432 1016 4433 1080
rect 4367 1000 4433 1016
rect 4367 936 4368 1000
rect 4432 936 4433 1000
rect 4367 920 4433 936
rect 4367 856 4368 920
rect 4432 856 4433 920
rect 4367 766 4433 856
rect 4493 702 4553 1732
rect 4613 762 4673 1794
rect 4733 702 4793 1732
rect 4853 762 4913 1794
rect 4973 1640 5039 1794
rect 4973 1576 4974 1640
rect 5038 1576 5039 1640
rect 4973 1560 5039 1576
rect 4973 1496 4974 1560
rect 5038 1496 5039 1560
rect 4973 1480 5039 1496
rect 4973 1416 4974 1480
rect 5038 1416 5039 1480
rect 4973 1400 5039 1416
rect 4973 1336 4974 1400
rect 5038 1336 5039 1400
rect 4973 1320 5039 1336
rect 4973 1256 4974 1320
rect 5038 1256 5039 1320
rect 4973 1240 5039 1256
rect 4973 1176 4974 1240
rect 5038 1176 5039 1240
rect 4973 1160 5039 1176
rect 4973 1096 4974 1160
rect 5038 1096 5039 1160
rect 4973 1080 5039 1096
rect 4973 1016 4974 1080
rect 5038 1016 5039 1080
rect 4973 1000 5039 1016
rect 4973 936 4974 1000
rect 5038 936 5039 1000
rect 4973 920 5039 936
rect 4973 856 4974 920
rect 5038 856 5039 920
rect 4973 766 5039 856
rect 5099 762 5159 1794
rect 5219 702 5279 1732
rect 5339 762 5399 1794
rect 5459 702 5519 1732
rect 5579 1640 5645 1794
rect 5579 1576 5580 1640
rect 5644 1576 5645 1640
rect 5579 1560 5645 1576
rect 5579 1496 5580 1560
rect 5644 1496 5645 1560
rect 5579 1480 5645 1496
rect 5579 1416 5580 1480
rect 5644 1416 5645 1480
rect 5579 1400 5645 1416
rect 5579 1336 5580 1400
rect 5644 1336 5645 1400
rect 5579 1320 5645 1336
rect 5579 1256 5580 1320
rect 5644 1256 5645 1320
rect 5579 1240 5645 1256
rect 5579 1176 5580 1240
rect 5644 1176 5645 1240
rect 5579 1160 5645 1176
rect 5579 1096 5580 1160
rect 5644 1096 5645 1160
rect 5579 1080 5645 1096
rect 5579 1016 5580 1080
rect 5644 1016 5645 1080
rect 5579 1000 5645 1016
rect 5579 936 5580 1000
rect 5644 936 5645 1000
rect 5579 920 5645 936
rect 5579 856 5580 920
rect 5644 856 5645 920
rect 5579 766 5645 856
rect 5705 1860 6377 1862
rect 5705 1796 5809 1860
rect 5873 1796 5889 1860
rect 5953 1796 5969 1860
rect 6033 1796 6049 1860
rect 6113 1796 6129 1860
rect 6193 1796 6209 1860
rect 6273 1796 6377 1860
rect 5705 1794 6377 1796
rect 5705 1640 5771 1794
rect 5705 1576 5706 1640
rect 5770 1576 5771 1640
rect 5705 1560 5771 1576
rect 5705 1496 5706 1560
rect 5770 1496 5771 1560
rect 5705 1480 5771 1496
rect 5705 1416 5706 1480
rect 5770 1416 5771 1480
rect 5705 1400 5771 1416
rect 5705 1336 5706 1400
rect 5770 1336 5771 1400
rect 5705 1320 5771 1336
rect 5705 1256 5706 1320
rect 5770 1256 5771 1320
rect 5705 1240 5771 1256
rect 5705 1176 5706 1240
rect 5770 1176 5771 1240
rect 5705 1160 5771 1176
rect 5705 1096 5706 1160
rect 5770 1096 5771 1160
rect 5705 1080 5771 1096
rect 5705 1016 5706 1080
rect 5770 1016 5771 1080
rect 5705 1000 5771 1016
rect 5705 936 5706 1000
rect 5770 936 5771 1000
rect 5705 920 5771 936
rect 5705 856 5706 920
rect 5770 856 5771 920
rect 5705 766 5771 856
rect 5831 762 5891 1794
rect 5951 702 6011 1732
rect 6071 762 6131 1794
rect 6191 702 6251 1732
rect 6311 1640 6377 1794
rect 6311 1576 6312 1640
rect 6376 1576 6377 1640
rect 6311 1560 6377 1576
rect 6311 1496 6312 1560
rect 6376 1496 6377 1560
rect 6311 1480 6377 1496
rect 6311 1416 6312 1480
rect 6376 1416 6377 1480
rect 6311 1400 6377 1416
rect 6311 1336 6312 1400
rect 6376 1336 6377 1400
rect 6311 1320 6377 1336
rect 6311 1256 6312 1320
rect 6376 1256 6377 1320
rect 6311 1240 6377 1256
rect 6311 1176 6312 1240
rect 6376 1176 6377 1240
rect 6311 1160 6377 1176
rect 6311 1096 6312 1160
rect 6376 1096 6377 1160
rect 6311 1080 6377 1096
rect 6311 1016 6312 1080
rect 6376 1016 6377 1080
rect 6311 1000 6377 1016
rect 6311 936 6312 1000
rect 6376 936 6377 1000
rect 6311 920 6377 936
rect 6311 856 6312 920
rect 6376 856 6377 920
rect 6311 766 6377 856
rect 6437 1633 6497 2014
rect 6638 1895 7198 2061
rect 7420 2111 7486 2265
rect 7546 2173 7606 3203
rect 7666 2111 7726 3143
rect 7786 2173 7846 3203
rect 7906 2111 7966 3143
rect 8026 3049 8092 3139
rect 8026 2985 8027 3049
rect 8091 2985 8092 3049
rect 8026 2969 8092 2985
rect 8026 2905 8027 2969
rect 8091 2905 8092 2969
rect 8026 2889 8092 2905
rect 8026 2825 8027 2889
rect 8091 2825 8092 2889
rect 8026 2809 8092 2825
rect 8026 2745 8027 2809
rect 8091 2745 8092 2809
rect 8026 2729 8092 2745
rect 8026 2665 8027 2729
rect 8091 2665 8092 2729
rect 8026 2649 8092 2665
rect 8026 2585 8027 2649
rect 8091 2585 8092 2649
rect 8026 2569 8092 2585
rect 8026 2505 8027 2569
rect 8091 2505 8092 2569
rect 8026 2489 8092 2505
rect 8026 2425 8027 2489
rect 8091 2425 8092 2489
rect 8026 2409 8092 2425
rect 8026 2345 8027 2409
rect 8091 2345 8092 2409
rect 8026 2329 8092 2345
rect 8026 2265 8027 2329
rect 8091 2265 8092 2329
rect 8026 2111 8092 2265
rect 7420 2109 8092 2111
rect 7420 2045 7524 2109
rect 7588 2045 7604 2109
rect 7668 2045 7684 2109
rect 7748 2045 7764 2109
rect 7828 2045 7844 2109
rect 7908 2045 7924 2109
rect 7988 2045 8092 2109
rect 7420 2043 8092 2045
rect 8152 3049 8218 3139
rect 8152 2985 8153 3049
rect 8217 2985 8218 3049
rect 8152 2969 8218 2985
rect 8152 2905 8153 2969
rect 8217 2905 8218 2969
rect 8152 2889 8218 2905
rect 8152 2825 8153 2889
rect 8217 2825 8218 2889
rect 8152 2809 8218 2825
rect 8152 2745 8153 2809
rect 8217 2745 8218 2809
rect 8152 2729 8218 2745
rect 8152 2665 8153 2729
rect 8217 2665 8218 2729
rect 8152 2649 8218 2665
rect 8152 2585 8153 2649
rect 8217 2585 8218 2649
rect 8152 2569 8218 2585
rect 8152 2505 8153 2569
rect 8217 2505 8218 2569
rect 8152 2489 8218 2505
rect 8152 2425 8153 2489
rect 8217 2425 8218 2489
rect 8152 2409 8218 2425
rect 8152 2345 8153 2409
rect 8217 2345 8218 2409
rect 8152 2329 8218 2345
rect 8152 2265 8153 2329
rect 8217 2265 8218 2329
rect 8152 2111 8218 2265
rect 8278 2173 8338 3203
rect 8398 2111 8458 3143
rect 8518 2173 8578 3203
rect 8638 2111 8698 3143
rect 8758 3049 8824 3139
rect 8758 2985 8759 3049
rect 8823 2985 8824 3049
rect 8758 2969 8824 2985
rect 8758 2905 8759 2969
rect 8823 2905 8824 2969
rect 8758 2889 8824 2905
rect 8758 2825 8759 2889
rect 8823 2825 8824 2889
rect 8758 2809 8824 2825
rect 8758 2745 8759 2809
rect 8823 2745 8824 2809
rect 8758 2729 8824 2745
rect 8758 2665 8759 2729
rect 8823 2665 8824 2729
rect 8758 2649 8824 2665
rect 8758 2585 8759 2649
rect 8823 2585 8824 2649
rect 8758 2569 8824 2585
rect 8758 2505 8759 2569
rect 8823 2505 8824 2569
rect 8758 2489 8824 2505
rect 8758 2425 8759 2489
rect 8823 2425 8824 2489
rect 8758 2409 8824 2425
rect 8758 2345 8759 2409
rect 8823 2345 8824 2409
rect 8758 2329 8824 2345
rect 8758 2265 8759 2329
rect 8823 2265 8824 2329
rect 8758 2111 8824 2265
rect 8884 2111 8944 3143
rect 9004 2173 9064 3203
rect 9124 2111 9184 3143
rect 9244 2173 9304 3203
rect 9364 3049 9430 3139
rect 9364 2985 9365 3049
rect 9429 2985 9430 3049
rect 9364 2969 9430 2985
rect 9364 2905 9365 2969
rect 9429 2905 9430 2969
rect 9364 2889 9430 2905
rect 9364 2825 9365 2889
rect 9429 2825 9430 2889
rect 9364 2809 9430 2825
rect 9364 2745 9365 2809
rect 9429 2745 9430 2809
rect 9364 2729 9430 2745
rect 9364 2665 9365 2729
rect 9429 2665 9430 2729
rect 9364 2649 9430 2665
rect 9364 2585 9365 2649
rect 9429 2585 9430 2649
rect 9364 2569 9430 2585
rect 9364 2505 9365 2569
rect 9429 2505 9430 2569
rect 9364 2489 9430 2505
rect 9364 2425 9365 2489
rect 9429 2425 9430 2489
rect 9364 2409 9430 2425
rect 9364 2345 9365 2409
rect 9429 2345 9430 2409
rect 9364 2329 9430 2345
rect 9364 2265 9365 2329
rect 9429 2265 9430 2329
rect 9364 2111 9430 2265
rect 9490 2173 9550 3203
rect 9610 2111 9670 3143
rect 9730 2173 9790 3203
rect 9850 2111 9910 3143
rect 9970 3049 10036 3139
rect 9970 2985 9971 3049
rect 10035 2985 10036 3049
rect 9970 2969 10036 2985
rect 9970 2905 9971 2969
rect 10035 2905 10036 2969
rect 9970 2889 10036 2905
rect 9970 2825 9971 2889
rect 10035 2825 10036 2889
rect 9970 2809 10036 2825
rect 9970 2745 9971 2809
rect 10035 2745 10036 2809
rect 9970 2729 10036 2745
rect 9970 2665 9971 2729
rect 10035 2665 10036 2729
rect 9970 2649 10036 2665
rect 9970 2585 9971 2649
rect 10035 2585 10036 2649
rect 9970 2569 10036 2585
rect 9970 2505 9971 2569
rect 10035 2505 10036 2569
rect 9970 2489 10036 2505
rect 9970 2425 9971 2489
rect 10035 2425 10036 2489
rect 9970 2409 10036 2425
rect 9970 2345 9971 2409
rect 10035 2345 10036 2409
rect 9970 2329 10036 2345
rect 9970 2265 9971 2329
rect 10035 2265 10036 2329
rect 9970 2111 10036 2265
rect 10096 2111 10156 3143
rect 10216 2173 10276 3203
rect 10336 2111 10396 3143
rect 10456 2173 10516 3203
rect 10576 3049 10642 3139
rect 10576 2985 10577 3049
rect 10641 2985 10642 3049
rect 10576 2969 10642 2985
rect 10576 2905 10577 2969
rect 10641 2905 10642 2969
rect 10576 2889 10642 2905
rect 10576 2825 10577 2889
rect 10641 2825 10642 2889
rect 10576 2809 10642 2825
rect 10576 2745 10577 2809
rect 10641 2745 10642 2809
rect 10576 2729 10642 2745
rect 10576 2665 10577 2729
rect 10641 2665 10642 2729
rect 10576 2649 10642 2665
rect 10576 2585 10577 2649
rect 10641 2585 10642 2649
rect 10576 2569 10642 2585
rect 10576 2505 10577 2569
rect 10641 2505 10642 2569
rect 10576 2489 10642 2505
rect 10576 2425 10577 2489
rect 10641 2425 10642 2489
rect 10576 2409 10642 2425
rect 10576 2345 10577 2409
rect 10641 2345 10642 2409
rect 10576 2329 10642 2345
rect 10576 2265 10577 2329
rect 10641 2265 10642 2329
rect 10576 2111 10642 2265
rect 10702 2173 10762 3203
rect 10822 2111 10882 3143
rect 10942 2173 11002 3203
rect 11062 2111 11122 3143
rect 11182 3049 11248 3139
rect 11182 2985 11183 3049
rect 11247 2985 11248 3049
rect 11182 2969 11248 2985
rect 11182 2905 11183 2969
rect 11247 2905 11248 2969
rect 11182 2889 11248 2905
rect 11182 2825 11183 2889
rect 11247 2825 11248 2889
rect 11182 2809 11248 2825
rect 11182 2745 11183 2809
rect 11247 2745 11248 2809
rect 11182 2729 11248 2745
rect 11182 2665 11183 2729
rect 11247 2665 11248 2729
rect 11182 2649 11248 2665
rect 11182 2585 11183 2649
rect 11247 2585 11248 2649
rect 11182 2569 11248 2585
rect 11182 2505 11183 2569
rect 11247 2505 11248 2569
rect 11182 2489 11248 2505
rect 11182 2425 11183 2489
rect 11247 2425 11248 2489
rect 11182 2409 11248 2425
rect 11182 2345 11183 2409
rect 11247 2345 11248 2409
rect 11182 2329 11248 2345
rect 11182 2265 11183 2329
rect 11247 2265 11248 2329
rect 11182 2111 11248 2265
rect 11308 2111 11368 3143
rect 11428 2173 11488 3203
rect 11548 2111 11608 3143
rect 11668 2173 11728 3203
rect 11788 3049 11854 3139
rect 11788 2985 11789 3049
rect 11853 2985 11854 3049
rect 11788 2969 11854 2985
rect 11788 2905 11789 2969
rect 11853 2905 11854 2969
rect 11788 2889 11854 2905
rect 11788 2825 11789 2889
rect 11853 2825 11854 2889
rect 11788 2809 11854 2825
rect 11788 2745 11789 2809
rect 11853 2745 11854 2809
rect 11788 2729 11854 2745
rect 11788 2665 11789 2729
rect 11853 2665 11854 2729
rect 11788 2649 11854 2665
rect 11788 2585 11789 2649
rect 11853 2585 11854 2649
rect 11788 2569 11854 2585
rect 11788 2505 11789 2569
rect 11853 2505 11854 2569
rect 11788 2489 11854 2505
rect 11788 2425 11789 2489
rect 11853 2425 11854 2489
rect 11788 2409 11854 2425
rect 11788 2345 11789 2409
rect 11853 2345 11854 2409
rect 11788 2329 11854 2345
rect 11788 2265 11789 2329
rect 11853 2265 11854 2329
rect 11788 2111 11854 2265
rect 11914 2173 11974 3203
rect 12034 2111 12094 3143
rect 12154 2173 12214 3203
rect 12274 2111 12334 3143
rect 12394 3049 12460 3139
rect 12394 2985 12395 3049
rect 12459 2985 12460 3049
rect 12394 2969 12460 2985
rect 12394 2905 12395 2969
rect 12459 2905 12460 2969
rect 12394 2889 12460 2905
rect 12394 2825 12395 2889
rect 12459 2825 12460 2889
rect 12394 2809 12460 2825
rect 12394 2745 12395 2809
rect 12459 2745 12460 2809
rect 12394 2729 12460 2745
rect 12394 2665 12395 2729
rect 12459 2665 12460 2729
rect 12394 2649 12460 2665
rect 12394 2585 12395 2649
rect 12459 2585 12460 2649
rect 12394 2569 12460 2585
rect 12394 2505 12395 2569
rect 12459 2505 12460 2569
rect 12394 2489 12460 2505
rect 12394 2425 12395 2489
rect 12459 2425 12460 2489
rect 12394 2409 12460 2425
rect 12394 2345 12395 2409
rect 12459 2345 12460 2409
rect 12394 2329 12460 2345
rect 12394 2265 12395 2329
rect 12459 2265 12460 2329
rect 12394 2111 12460 2265
rect 12520 2111 12580 3143
rect 12640 2173 12700 3203
rect 12760 2111 12820 3143
rect 12880 2173 12940 3203
rect 13000 3049 13066 3139
rect 13000 2985 13001 3049
rect 13065 2985 13066 3049
rect 13000 2969 13066 2985
rect 13000 2905 13001 2969
rect 13065 2905 13066 2969
rect 13000 2889 13066 2905
rect 13000 2825 13001 2889
rect 13065 2825 13066 2889
rect 13000 2809 13066 2825
rect 13000 2745 13001 2809
rect 13065 2745 13066 2809
rect 13000 2729 13066 2745
rect 13000 2665 13001 2729
rect 13065 2665 13066 2729
rect 13000 2649 13066 2665
rect 13000 2585 13001 2649
rect 13065 2585 13066 2649
rect 13000 2569 13066 2585
rect 13000 2505 13001 2569
rect 13065 2505 13066 2569
rect 13000 2489 13066 2505
rect 13000 2425 13001 2489
rect 13065 2425 13066 2489
rect 13000 2409 13066 2425
rect 13000 2345 13001 2409
rect 13065 2345 13066 2409
rect 13000 2329 13066 2345
rect 13000 2265 13001 2329
rect 13065 2265 13066 2329
rect 13126 2349 13444 3203
rect 13126 2285 13159 2349
rect 13223 2285 13444 2349
rect 13126 2273 13444 2285
rect 13000 2111 13066 2265
rect 8152 2109 13066 2111
rect 8152 2045 8256 2109
rect 8320 2045 8336 2109
rect 8400 2045 8416 2109
rect 8480 2045 8496 2109
rect 8560 2045 8576 2109
rect 8640 2045 8656 2109
rect 8720 2045 8862 2109
rect 8926 2045 8942 2109
rect 9006 2045 9022 2109
rect 9086 2045 9102 2109
rect 9166 2045 9182 2109
rect 9246 2045 9262 2109
rect 9326 2045 9468 2109
rect 9532 2045 9548 2109
rect 9612 2045 9628 2109
rect 9692 2045 9708 2109
rect 9772 2045 9788 2109
rect 9852 2045 9868 2109
rect 9932 2045 10074 2109
rect 10138 2045 10154 2109
rect 10218 2045 10234 2109
rect 10298 2045 10314 2109
rect 10378 2045 10394 2109
rect 10458 2045 10474 2109
rect 10538 2045 10680 2109
rect 10744 2045 10760 2109
rect 10824 2045 10840 2109
rect 10904 2045 10920 2109
rect 10984 2045 11000 2109
rect 11064 2045 11080 2109
rect 11144 2045 11286 2109
rect 11350 2045 11366 2109
rect 11430 2045 11446 2109
rect 11510 2045 11526 2109
rect 11590 2045 11606 2109
rect 11670 2045 11686 2109
rect 11750 2045 11892 2109
rect 11956 2045 11972 2109
rect 12036 2045 12052 2109
rect 12116 2045 12132 2109
rect 12196 2045 12212 2109
rect 12276 2045 12292 2109
rect 12356 2045 12498 2109
rect 12562 2045 12578 2109
rect 12642 2045 12658 2109
rect 12722 2045 12738 2109
rect 12802 2045 12818 2109
rect 12882 2045 12898 2109
rect 12962 2045 13066 2109
rect 8152 2043 13066 2045
rect 13126 2088 13324 2098
rect 6557 1885 7198 1895
rect 6557 1821 6558 1885
rect 6622 1821 7198 1885
rect 13126 2024 13247 2088
rect 13311 2024 13324 2088
rect 13126 2014 13324 2024
rect 6557 1811 7198 1821
rect 6638 1633 7198 1811
rect 6437 1623 7198 1633
rect 6437 1559 6467 1623
rect 6531 1559 7198 1623
rect 6437 702 7198 1559
rect 7774 1860 8446 1862
rect 7774 1796 7878 1860
rect 7942 1796 7958 1860
rect 8022 1796 8038 1860
rect 8102 1796 8118 1860
rect 8182 1796 8198 1860
rect 8262 1796 8278 1860
rect 8342 1796 8446 1860
rect 7774 1794 8446 1796
rect 7774 1640 7840 1794
rect 7774 1576 7775 1640
rect 7839 1576 7840 1640
rect 7774 1560 7840 1576
rect 7774 1496 7775 1560
rect 7839 1496 7840 1560
rect 7774 1480 7840 1496
rect 7774 1416 7775 1480
rect 7839 1416 7840 1480
rect 7774 1400 7840 1416
rect 7774 1336 7775 1400
rect 7839 1336 7840 1400
rect 7774 1320 7840 1336
rect 7774 1256 7775 1320
rect 7839 1256 7840 1320
rect 7774 1240 7840 1256
rect 7774 1176 7775 1240
rect 7839 1176 7840 1240
rect 7774 1160 7840 1176
rect 7774 1096 7775 1160
rect 7839 1096 7840 1160
rect 7774 1080 7840 1096
rect 7774 1016 7775 1080
rect 7839 1016 7840 1080
rect 7774 1000 7840 1016
rect 7774 936 7775 1000
rect 7839 936 7840 1000
rect 7774 920 7840 936
rect 7774 856 7775 920
rect 7839 856 7840 920
rect 7774 766 7840 856
rect 7383 702 7508 708
rect 7900 702 7960 1732
rect 8020 762 8080 1794
rect 8140 702 8200 1732
rect 8260 762 8320 1794
rect 8380 1640 8446 1794
rect 8380 1576 8381 1640
rect 8445 1576 8446 1640
rect 8380 1560 8446 1576
rect 8380 1496 8381 1560
rect 8445 1496 8446 1560
rect 8380 1480 8446 1496
rect 8380 1416 8381 1480
rect 8445 1416 8446 1480
rect 8380 1400 8446 1416
rect 8380 1336 8381 1400
rect 8445 1336 8446 1400
rect 8380 1320 8446 1336
rect 8380 1256 8381 1320
rect 8445 1256 8446 1320
rect 8380 1240 8446 1256
rect 8380 1176 8381 1240
rect 8445 1176 8446 1240
rect 8380 1160 8446 1176
rect 8380 1096 8381 1160
rect 8445 1096 8446 1160
rect 8380 1080 8446 1096
rect 8380 1016 8381 1080
rect 8445 1016 8446 1080
rect 8380 1000 8446 1016
rect 8380 936 8381 1000
rect 8445 936 8446 1000
rect 8380 920 8446 936
rect 8380 856 8381 920
rect 8445 856 8446 920
rect 8380 766 8446 856
rect 8506 1860 10996 1862
rect 8506 1796 8610 1860
rect 8674 1796 8690 1860
rect 8754 1796 8770 1860
rect 8834 1796 8850 1860
rect 8914 1796 8930 1860
rect 8994 1796 9010 1860
rect 9074 1796 9216 1860
rect 9280 1796 9296 1860
rect 9360 1796 9376 1860
rect 9440 1796 9456 1860
rect 9520 1796 9536 1860
rect 9600 1796 9616 1860
rect 9680 1796 9822 1860
rect 9886 1796 9902 1860
rect 9966 1796 9982 1860
rect 10046 1796 10062 1860
rect 10126 1796 10142 1860
rect 10206 1796 10222 1860
rect 10286 1796 10428 1860
rect 10492 1796 10508 1860
rect 10572 1796 10588 1860
rect 10652 1796 10668 1860
rect 10732 1796 10748 1860
rect 10812 1796 10828 1860
rect 10892 1796 10996 1860
rect 8506 1794 10996 1796
rect 8506 1640 8572 1794
rect 8506 1576 8507 1640
rect 8571 1576 8572 1640
rect 8506 1560 8572 1576
rect 8506 1496 8507 1560
rect 8571 1496 8572 1560
rect 8506 1480 8572 1496
rect 8506 1416 8507 1480
rect 8571 1416 8572 1480
rect 8506 1400 8572 1416
rect 8506 1336 8507 1400
rect 8571 1336 8572 1400
rect 8506 1320 8572 1336
rect 8506 1256 8507 1320
rect 8571 1256 8572 1320
rect 8506 1240 8572 1256
rect 8506 1176 8507 1240
rect 8571 1176 8572 1240
rect 8506 1160 8572 1176
rect 8506 1096 8507 1160
rect 8571 1096 8572 1160
rect 8506 1080 8572 1096
rect 8506 1016 8507 1080
rect 8571 1016 8572 1080
rect 8506 1000 8572 1016
rect 8506 936 8507 1000
rect 8571 936 8572 1000
rect 8506 920 8572 936
rect 8506 856 8507 920
rect 8571 856 8572 920
rect 8506 766 8572 856
rect 8632 702 8692 1732
rect 8752 762 8812 1794
rect 8872 702 8932 1732
rect 8992 762 9052 1794
rect 9112 1640 9178 1794
rect 9112 1576 9113 1640
rect 9177 1576 9178 1640
rect 9112 1560 9178 1576
rect 9112 1496 9113 1560
rect 9177 1496 9178 1560
rect 9112 1480 9178 1496
rect 9112 1416 9113 1480
rect 9177 1416 9178 1480
rect 9112 1400 9178 1416
rect 9112 1336 9113 1400
rect 9177 1336 9178 1400
rect 9112 1320 9178 1336
rect 9112 1256 9113 1320
rect 9177 1256 9178 1320
rect 9112 1240 9178 1256
rect 9112 1176 9113 1240
rect 9177 1176 9178 1240
rect 9112 1160 9178 1176
rect 9112 1096 9113 1160
rect 9177 1096 9178 1160
rect 9112 1080 9178 1096
rect 9112 1016 9113 1080
rect 9177 1016 9178 1080
rect 9112 1000 9178 1016
rect 9112 936 9113 1000
rect 9177 936 9178 1000
rect 9112 920 9178 936
rect 9112 856 9113 920
rect 9177 856 9178 920
rect 9112 766 9178 856
rect 9238 762 9298 1794
rect 9358 702 9418 1732
rect 9478 762 9538 1794
rect 9598 702 9658 1732
rect 9718 1640 9784 1794
rect 9718 1576 9719 1640
rect 9783 1576 9784 1640
rect 9718 1560 9784 1576
rect 9718 1496 9719 1560
rect 9783 1496 9784 1560
rect 9718 1480 9784 1496
rect 9718 1416 9719 1480
rect 9783 1416 9784 1480
rect 9718 1400 9784 1416
rect 9718 1336 9719 1400
rect 9783 1336 9784 1400
rect 9718 1320 9784 1336
rect 9718 1256 9719 1320
rect 9783 1256 9784 1320
rect 9718 1240 9784 1256
rect 9718 1176 9719 1240
rect 9783 1176 9784 1240
rect 9718 1160 9784 1176
rect 9718 1096 9719 1160
rect 9783 1096 9784 1160
rect 9718 1080 9784 1096
rect 9718 1016 9719 1080
rect 9783 1016 9784 1080
rect 9718 1000 9784 1016
rect 9718 936 9719 1000
rect 9783 936 9784 1000
rect 9718 920 9784 936
rect 9718 856 9719 920
rect 9783 856 9784 920
rect 9718 766 9784 856
rect 9844 702 9904 1732
rect 9964 762 10024 1794
rect 10084 702 10144 1732
rect 10204 762 10264 1794
rect 10324 1640 10390 1794
rect 10324 1576 10325 1640
rect 10389 1576 10390 1640
rect 10324 1560 10390 1576
rect 10324 1496 10325 1560
rect 10389 1496 10390 1560
rect 10324 1480 10390 1496
rect 10324 1416 10325 1480
rect 10389 1416 10390 1480
rect 10324 1400 10390 1416
rect 10324 1336 10325 1400
rect 10389 1336 10390 1400
rect 10324 1320 10390 1336
rect 10324 1256 10325 1320
rect 10389 1256 10390 1320
rect 10324 1240 10390 1256
rect 10324 1176 10325 1240
rect 10389 1176 10390 1240
rect 10324 1160 10390 1176
rect 10324 1096 10325 1160
rect 10389 1096 10390 1160
rect 10324 1080 10390 1096
rect 10324 1016 10325 1080
rect 10389 1016 10390 1080
rect 10324 1000 10390 1016
rect 10324 936 10325 1000
rect 10389 936 10390 1000
rect 10324 920 10390 936
rect 10324 856 10325 920
rect 10389 856 10390 920
rect 10324 766 10390 856
rect 10450 762 10510 1794
rect 10570 702 10630 1732
rect 10690 762 10750 1794
rect 10810 702 10870 1732
rect 10930 1640 10996 1794
rect 10930 1576 10931 1640
rect 10995 1576 10996 1640
rect 10930 1560 10996 1576
rect 10930 1496 10931 1560
rect 10995 1496 10996 1560
rect 10930 1480 10996 1496
rect 10930 1416 10931 1480
rect 10995 1416 10996 1480
rect 10930 1400 10996 1416
rect 10930 1336 10931 1400
rect 10995 1336 10996 1400
rect 10930 1320 10996 1336
rect 10930 1256 10931 1320
rect 10995 1256 10996 1320
rect 10930 1240 10996 1256
rect 10930 1176 10931 1240
rect 10995 1176 10996 1240
rect 10930 1160 10996 1176
rect 10930 1096 10931 1160
rect 10995 1096 10996 1160
rect 10930 1080 10996 1096
rect 10930 1016 10931 1080
rect 10995 1016 10996 1080
rect 10930 1000 10996 1016
rect 10930 936 10931 1000
rect 10995 936 10996 1000
rect 10930 920 10996 936
rect 10930 856 10931 920
rect 10995 856 10996 920
rect 10930 766 10996 856
rect 11056 1860 12334 1862
rect 11056 1796 11160 1860
rect 11224 1796 11240 1860
rect 11304 1796 11320 1860
rect 11384 1796 11400 1860
rect 11464 1796 11480 1860
rect 11544 1796 11560 1860
rect 11624 1796 11766 1860
rect 11830 1796 11846 1860
rect 11910 1796 11926 1860
rect 11990 1796 12006 1860
rect 12070 1796 12086 1860
rect 12150 1796 12166 1860
rect 12230 1796 12334 1860
rect 11056 1794 12334 1796
rect 11056 1640 11122 1794
rect 11056 1576 11057 1640
rect 11121 1576 11122 1640
rect 11056 1560 11122 1576
rect 11056 1496 11057 1560
rect 11121 1496 11122 1560
rect 11056 1480 11122 1496
rect 11056 1416 11057 1480
rect 11121 1416 11122 1480
rect 11056 1400 11122 1416
rect 11056 1336 11057 1400
rect 11121 1336 11122 1400
rect 11056 1320 11122 1336
rect 11056 1256 11057 1320
rect 11121 1256 11122 1320
rect 11056 1240 11122 1256
rect 11056 1176 11057 1240
rect 11121 1176 11122 1240
rect 11056 1160 11122 1176
rect 11056 1096 11057 1160
rect 11121 1096 11122 1160
rect 11056 1080 11122 1096
rect 11056 1016 11057 1080
rect 11121 1016 11122 1080
rect 11056 1000 11122 1016
rect 11056 936 11057 1000
rect 11121 936 11122 1000
rect 11056 920 11122 936
rect 11056 856 11057 920
rect 11121 856 11122 920
rect 11056 766 11122 856
rect 11182 702 11242 1732
rect 11302 762 11362 1794
rect 11422 702 11482 1732
rect 11542 762 11602 1794
rect 11662 1640 11728 1794
rect 11662 1576 11663 1640
rect 11727 1576 11728 1640
rect 11662 1560 11728 1576
rect 11662 1496 11663 1560
rect 11727 1496 11728 1560
rect 11662 1480 11728 1496
rect 11662 1416 11663 1480
rect 11727 1416 11728 1480
rect 11662 1400 11728 1416
rect 11662 1336 11663 1400
rect 11727 1336 11728 1400
rect 11662 1320 11728 1336
rect 11662 1256 11663 1320
rect 11727 1256 11728 1320
rect 11662 1240 11728 1256
rect 11662 1176 11663 1240
rect 11727 1176 11728 1240
rect 11662 1160 11728 1176
rect 11662 1096 11663 1160
rect 11727 1096 11728 1160
rect 11662 1080 11728 1096
rect 11662 1016 11663 1080
rect 11727 1016 11728 1080
rect 11662 1000 11728 1016
rect 11662 936 11663 1000
rect 11727 936 11728 1000
rect 11662 920 11728 936
rect 11662 856 11663 920
rect 11727 856 11728 920
rect 11662 766 11728 856
rect 11788 762 11848 1794
rect 11908 702 11968 1732
rect 12028 762 12088 1794
rect 12148 702 12208 1732
rect 12268 1640 12334 1794
rect 12268 1576 12269 1640
rect 12333 1576 12334 1640
rect 12268 1560 12334 1576
rect 12268 1496 12269 1560
rect 12333 1496 12334 1560
rect 12268 1480 12334 1496
rect 12268 1416 12269 1480
rect 12333 1416 12334 1480
rect 12268 1400 12334 1416
rect 12268 1336 12269 1400
rect 12333 1336 12334 1400
rect 12268 1320 12334 1336
rect 12268 1256 12269 1320
rect 12333 1256 12334 1320
rect 12268 1240 12334 1256
rect 12268 1176 12269 1240
rect 12333 1176 12334 1240
rect 12268 1160 12334 1176
rect 12268 1096 12269 1160
rect 12333 1096 12334 1160
rect 12268 1080 12334 1096
rect 12268 1016 12269 1080
rect 12333 1016 12334 1080
rect 12268 1000 12334 1016
rect 12268 936 12269 1000
rect 12333 936 12334 1000
rect 12268 920 12334 936
rect 12268 856 12269 920
rect 12333 856 12334 920
rect 12268 766 12334 856
rect 12394 1860 13066 1862
rect 12394 1796 12498 1860
rect 12562 1796 12578 1860
rect 12642 1796 12658 1860
rect 12722 1796 12738 1860
rect 12802 1796 12818 1860
rect 12882 1796 12898 1860
rect 12962 1796 13066 1860
rect 12394 1794 13066 1796
rect 12394 1640 12460 1794
rect 12394 1576 12395 1640
rect 12459 1576 12460 1640
rect 12394 1560 12460 1576
rect 12394 1496 12395 1560
rect 12459 1496 12460 1560
rect 12394 1480 12460 1496
rect 12394 1416 12395 1480
rect 12459 1416 12460 1480
rect 12394 1400 12460 1416
rect 12394 1336 12395 1400
rect 12459 1336 12460 1400
rect 12394 1320 12460 1336
rect 12394 1256 12395 1320
rect 12459 1256 12460 1320
rect 12394 1240 12460 1256
rect 12394 1176 12395 1240
rect 12459 1176 12460 1240
rect 12394 1160 12460 1176
rect 12394 1096 12395 1160
rect 12459 1096 12460 1160
rect 12394 1080 12460 1096
rect 12394 1016 12395 1080
rect 12459 1016 12460 1080
rect 12394 1000 12460 1016
rect 12394 936 12395 1000
rect 12459 936 12460 1000
rect 12394 920 12460 936
rect 12394 856 12395 920
rect 12459 856 12460 920
rect 12394 766 12460 856
rect 12520 762 12580 1794
rect 12640 702 12700 1732
rect 12760 762 12820 1794
rect 12880 702 12940 1732
rect 13000 1640 13066 1794
rect 13000 1576 13001 1640
rect 13065 1576 13066 1640
rect 13000 1560 13066 1576
rect 13000 1496 13001 1560
rect 13065 1496 13066 1560
rect 13000 1480 13066 1496
rect 13000 1416 13001 1480
rect 13065 1416 13066 1480
rect 13000 1400 13066 1416
rect 13000 1336 13001 1400
rect 13065 1336 13066 1400
rect 13000 1320 13066 1336
rect 13000 1256 13001 1320
rect 13065 1256 13066 1320
rect 13000 1240 13066 1256
rect 13000 1176 13001 1240
rect 13065 1176 13066 1240
rect 13000 1160 13066 1176
rect 13000 1096 13001 1160
rect 13065 1096 13066 1160
rect 13000 1080 13066 1096
rect 13000 1016 13001 1080
rect 13065 1016 13066 1080
rect 13000 1000 13066 1016
rect 13000 936 13001 1000
rect 13065 936 13066 1000
rect 13000 920 13066 936
rect 13000 856 13001 920
rect 13065 856 13066 920
rect 13000 766 13066 856
rect 13126 1633 13186 2014
rect 13384 1895 13444 2273
rect 13246 1885 13444 1895
rect 13246 1821 13247 1885
rect 13311 1821 13444 1885
rect 13246 1811 13444 1821
rect 13126 1623 13444 1633
rect 13126 1559 13156 1623
rect 13220 1559 13444 1623
rect 13126 702 13444 1559
rect 78 700 13444 702
rect 78 698 1189 700
rect 78 634 724 698
rect 788 636 1189 698
rect 1253 636 1269 700
rect 1333 636 1349 700
rect 1413 636 1429 700
rect 1493 636 1509 700
rect 1573 636 1589 700
rect 1653 636 1921 700
rect 1985 636 2001 700
rect 2065 636 2081 700
rect 2145 636 2161 700
rect 2225 636 2241 700
rect 2305 636 2321 700
rect 2385 636 2527 700
rect 2591 636 2607 700
rect 2671 636 2687 700
rect 2751 636 2767 700
rect 2831 636 2847 700
rect 2911 636 2927 700
rect 2991 636 3133 700
rect 3197 636 3213 700
rect 3277 636 3293 700
rect 3357 636 3373 700
rect 3437 636 3453 700
rect 3517 636 3533 700
rect 3597 636 3739 700
rect 3803 636 3819 700
rect 3883 636 3899 700
rect 3963 636 3979 700
rect 4043 636 4059 700
rect 4123 636 4139 700
rect 4203 636 4471 700
rect 4535 636 4551 700
rect 4615 636 4631 700
rect 4695 636 4711 700
rect 4775 636 4791 700
rect 4855 636 4871 700
rect 4935 636 5077 700
rect 5141 636 5157 700
rect 5221 636 5237 700
rect 5301 636 5317 700
rect 5381 636 5397 700
rect 5461 636 5477 700
rect 5541 636 5809 700
rect 5873 636 5889 700
rect 5953 636 5969 700
rect 6033 636 6049 700
rect 6113 636 6129 700
rect 6193 636 6209 700
rect 6273 698 7878 700
rect 6273 636 7413 698
rect 788 634 7413 636
rect 7477 636 7878 698
rect 7942 636 7958 700
rect 8022 636 8038 700
rect 8102 636 8118 700
rect 8182 636 8198 700
rect 8262 636 8278 700
rect 8342 636 8610 700
rect 8674 636 8690 700
rect 8754 636 8770 700
rect 8834 636 8850 700
rect 8914 636 8930 700
rect 8994 636 9010 700
rect 9074 636 9216 700
rect 9280 636 9296 700
rect 9360 636 9376 700
rect 9440 636 9456 700
rect 9520 636 9536 700
rect 9600 636 9616 700
rect 9680 636 9822 700
rect 9886 636 9902 700
rect 9966 636 9982 700
rect 10046 636 10062 700
rect 10126 636 10142 700
rect 10206 636 10222 700
rect 10286 636 10428 700
rect 10492 636 10508 700
rect 10572 636 10588 700
rect 10652 636 10668 700
rect 10732 636 10748 700
rect 10812 636 10828 700
rect 10892 636 11160 700
rect 11224 636 11240 700
rect 11304 636 11320 700
rect 11384 636 11400 700
rect 11464 636 11480 700
rect 11544 636 11560 700
rect 11624 636 11766 700
rect 11830 636 11846 700
rect 11910 636 11926 700
rect 11990 636 12006 700
rect 12070 636 12086 700
rect 12150 636 12166 700
rect 12230 636 12498 700
rect 12562 636 12578 700
rect 12642 636 12658 700
rect 12722 636 12738 700
rect 12802 636 12818 700
rect 12882 636 12898 700
rect 12962 636 13444 700
rect 7477 634 13444 636
rect 78 624 13444 634
rect 78 622 574 624
rect 6638 622 7263 624
rect 6638 614 6866 622
rect 6275 324 6771 326
rect 13030 324 13526 326
rect 94 314 6771 324
rect 94 312 6061 314
rect 94 248 576 312
rect 640 248 656 312
rect 720 248 736 312
rect 800 248 816 312
rect 880 248 896 312
rect 960 248 976 312
rect 1040 248 1308 312
rect 1372 248 1388 312
rect 1452 248 1468 312
rect 1532 248 1548 312
rect 1612 248 1628 312
rect 1692 248 1708 312
rect 1772 248 1914 312
rect 1978 248 1994 312
rect 2058 248 2074 312
rect 2138 248 2154 312
rect 2218 248 2234 312
rect 2298 248 2314 312
rect 2378 248 2646 312
rect 2710 248 2726 312
rect 2790 248 2806 312
rect 2870 248 2886 312
rect 2950 248 2966 312
rect 3030 248 3046 312
rect 3110 248 3252 312
rect 3316 248 3332 312
rect 3396 248 3412 312
rect 3476 248 3492 312
rect 3556 248 3572 312
rect 3636 248 3652 312
rect 3716 248 3858 312
rect 3922 248 3938 312
rect 4002 248 4018 312
rect 4082 248 4098 312
rect 4162 248 4178 312
rect 4242 248 4258 312
rect 4322 248 4464 312
rect 4528 248 4544 312
rect 4608 248 4624 312
rect 4688 248 4704 312
rect 4768 248 4784 312
rect 4848 248 4864 312
rect 4928 248 5196 312
rect 5260 248 5276 312
rect 5340 248 5356 312
rect 5420 248 5436 312
rect 5500 248 5516 312
rect 5580 248 5596 312
rect 5660 250 6061 312
rect 6125 250 6771 314
rect 5660 248 6771 250
rect 94 246 6771 248
rect 6849 314 13526 324
rect 6849 312 12816 314
rect 6849 248 7331 312
rect 7395 248 7411 312
rect 7475 248 7491 312
rect 7555 248 7571 312
rect 7635 248 7651 312
rect 7715 248 7731 312
rect 7795 248 8063 312
rect 8127 248 8143 312
rect 8207 248 8223 312
rect 8287 248 8303 312
rect 8367 248 8383 312
rect 8447 248 8463 312
rect 8527 248 8669 312
rect 8733 248 8749 312
rect 8813 248 8829 312
rect 8893 248 8909 312
rect 8973 248 8989 312
rect 9053 248 9069 312
rect 9133 248 9401 312
rect 9465 248 9481 312
rect 9545 248 9561 312
rect 9625 248 9641 312
rect 9705 248 9721 312
rect 9785 248 9801 312
rect 9865 248 10007 312
rect 10071 248 10087 312
rect 10151 248 10167 312
rect 10231 248 10247 312
rect 10311 248 10327 312
rect 10391 248 10407 312
rect 10471 248 10613 312
rect 10677 248 10693 312
rect 10757 248 10773 312
rect 10837 248 10853 312
rect 10917 248 10933 312
rect 10997 248 11013 312
rect 11077 248 11219 312
rect 11283 248 11299 312
rect 11363 248 11379 312
rect 11443 248 11459 312
rect 11523 248 11539 312
rect 11603 248 11619 312
rect 11683 248 11951 312
rect 12015 248 12031 312
rect 12095 248 12111 312
rect 12175 248 12191 312
rect 12255 248 12271 312
rect 12335 248 12351 312
rect 12415 250 12816 312
rect 12880 250 13526 314
rect 12415 248 13526 250
rect 6849 246 13526 248
rect 94 -611 412 246
rect 94 -675 318 -611
rect 382 -675 412 -611
rect 94 -685 412 -675
rect 94 -873 292 -863
rect 94 -937 227 -873
rect 291 -937 292 -873
rect 94 -947 292 -937
rect 94 -1325 154 -947
rect 352 -1066 412 -685
rect 472 92 538 182
rect 472 28 473 92
rect 537 28 538 92
rect 472 12 538 28
rect 472 -52 473 12
rect 537 -52 538 12
rect 472 -68 538 -52
rect 472 -132 473 -68
rect 537 -132 538 -68
rect 472 -148 538 -132
rect 472 -212 473 -148
rect 537 -212 538 -148
rect 472 -228 538 -212
rect 472 -292 473 -228
rect 537 -292 538 -228
rect 472 -308 538 -292
rect 472 -372 473 -308
rect 537 -372 538 -308
rect 472 -388 538 -372
rect 472 -452 473 -388
rect 537 -452 538 -388
rect 472 -468 538 -452
rect 472 -532 473 -468
rect 537 -532 538 -468
rect 472 -548 538 -532
rect 472 -612 473 -548
rect 537 -612 538 -548
rect 472 -628 538 -612
rect 472 -692 473 -628
rect 537 -692 538 -628
rect 472 -846 538 -692
rect 598 -784 658 246
rect 718 -846 778 186
rect 838 -784 898 246
rect 958 -846 1018 186
rect 1078 92 1144 182
rect 1078 28 1079 92
rect 1143 28 1144 92
rect 1078 12 1144 28
rect 1078 -52 1079 12
rect 1143 -52 1144 12
rect 1078 -68 1144 -52
rect 1078 -132 1079 -68
rect 1143 -132 1144 -68
rect 1078 -148 1144 -132
rect 1078 -212 1079 -148
rect 1143 -212 1144 -148
rect 1078 -228 1144 -212
rect 1078 -292 1079 -228
rect 1143 -292 1144 -228
rect 1078 -308 1144 -292
rect 1078 -372 1079 -308
rect 1143 -372 1144 -308
rect 1078 -388 1144 -372
rect 1078 -452 1079 -388
rect 1143 -452 1144 -388
rect 1078 -468 1144 -452
rect 1078 -532 1079 -468
rect 1143 -532 1144 -468
rect 1078 -548 1144 -532
rect 1078 -612 1079 -548
rect 1143 -612 1144 -548
rect 1078 -628 1144 -612
rect 1078 -692 1079 -628
rect 1143 -692 1144 -628
rect 1078 -846 1144 -692
rect 472 -848 1144 -846
rect 472 -912 576 -848
rect 640 -912 656 -848
rect 720 -912 736 -848
rect 800 -912 816 -848
rect 880 -912 896 -848
rect 960 -912 976 -848
rect 1040 -912 1144 -848
rect 472 -914 1144 -912
rect 1204 92 1270 182
rect 1204 28 1205 92
rect 1269 28 1270 92
rect 1204 12 1270 28
rect 1204 -52 1205 12
rect 1269 -52 1270 12
rect 1204 -68 1270 -52
rect 1204 -132 1205 -68
rect 1269 -132 1270 -68
rect 1204 -148 1270 -132
rect 1204 -212 1205 -148
rect 1269 -212 1270 -148
rect 1204 -228 1270 -212
rect 1204 -292 1205 -228
rect 1269 -292 1270 -228
rect 1204 -308 1270 -292
rect 1204 -372 1205 -308
rect 1269 -372 1270 -308
rect 1204 -388 1270 -372
rect 1204 -452 1205 -388
rect 1269 -452 1270 -388
rect 1204 -468 1270 -452
rect 1204 -532 1205 -468
rect 1269 -532 1270 -468
rect 1204 -548 1270 -532
rect 1204 -612 1205 -548
rect 1269 -612 1270 -548
rect 1204 -628 1270 -612
rect 1204 -692 1205 -628
rect 1269 -692 1270 -628
rect 1204 -846 1270 -692
rect 1330 -784 1390 246
rect 1450 -846 1510 186
rect 1570 -784 1630 246
rect 1690 -846 1750 186
rect 1810 92 1876 182
rect 1810 28 1811 92
rect 1875 28 1876 92
rect 1810 12 1876 28
rect 1810 -52 1811 12
rect 1875 -52 1876 12
rect 1810 -68 1876 -52
rect 1810 -132 1811 -68
rect 1875 -132 1876 -68
rect 1810 -148 1876 -132
rect 1810 -212 1811 -148
rect 1875 -212 1876 -148
rect 1810 -228 1876 -212
rect 1810 -292 1811 -228
rect 1875 -292 1876 -228
rect 1810 -308 1876 -292
rect 1810 -372 1811 -308
rect 1875 -372 1876 -308
rect 1810 -388 1876 -372
rect 1810 -452 1811 -388
rect 1875 -452 1876 -388
rect 1810 -468 1876 -452
rect 1810 -532 1811 -468
rect 1875 -532 1876 -468
rect 1810 -548 1876 -532
rect 1810 -612 1811 -548
rect 1875 -612 1876 -548
rect 1810 -628 1876 -612
rect 1810 -692 1811 -628
rect 1875 -692 1876 -628
rect 1810 -846 1876 -692
rect 1936 -846 1996 186
rect 2056 -784 2116 246
rect 2176 -846 2236 186
rect 2296 -784 2356 246
rect 2416 92 2482 182
rect 2416 28 2417 92
rect 2481 28 2482 92
rect 2416 12 2482 28
rect 2416 -52 2417 12
rect 2481 -52 2482 12
rect 2416 -68 2482 -52
rect 2416 -132 2417 -68
rect 2481 -132 2482 -68
rect 2416 -148 2482 -132
rect 2416 -212 2417 -148
rect 2481 -212 2482 -148
rect 2416 -228 2482 -212
rect 2416 -292 2417 -228
rect 2481 -292 2482 -228
rect 2416 -308 2482 -292
rect 2416 -372 2417 -308
rect 2481 -372 2482 -308
rect 2416 -388 2482 -372
rect 2416 -452 2417 -388
rect 2481 -452 2482 -388
rect 2416 -468 2482 -452
rect 2416 -532 2417 -468
rect 2481 -532 2482 -468
rect 2416 -548 2482 -532
rect 2416 -612 2417 -548
rect 2481 -612 2482 -548
rect 2416 -628 2482 -612
rect 2416 -692 2417 -628
rect 2481 -692 2482 -628
rect 2416 -846 2482 -692
rect 1204 -848 2482 -846
rect 1204 -912 1308 -848
rect 1372 -912 1388 -848
rect 1452 -912 1468 -848
rect 1532 -912 1548 -848
rect 1612 -912 1628 -848
rect 1692 -912 1708 -848
rect 1772 -912 1914 -848
rect 1978 -912 1994 -848
rect 2058 -912 2074 -848
rect 2138 -912 2154 -848
rect 2218 -912 2234 -848
rect 2298 -912 2314 -848
rect 2378 -912 2482 -848
rect 1204 -914 2482 -912
rect 2542 92 2608 182
rect 2542 28 2543 92
rect 2607 28 2608 92
rect 2542 12 2608 28
rect 2542 -52 2543 12
rect 2607 -52 2608 12
rect 2542 -68 2608 -52
rect 2542 -132 2543 -68
rect 2607 -132 2608 -68
rect 2542 -148 2608 -132
rect 2542 -212 2543 -148
rect 2607 -212 2608 -148
rect 2542 -228 2608 -212
rect 2542 -292 2543 -228
rect 2607 -292 2608 -228
rect 2542 -308 2608 -292
rect 2542 -372 2543 -308
rect 2607 -372 2608 -308
rect 2542 -388 2608 -372
rect 2542 -452 2543 -388
rect 2607 -452 2608 -388
rect 2542 -468 2608 -452
rect 2542 -532 2543 -468
rect 2607 -532 2608 -468
rect 2542 -548 2608 -532
rect 2542 -612 2543 -548
rect 2607 -612 2608 -548
rect 2542 -628 2608 -612
rect 2542 -692 2543 -628
rect 2607 -692 2608 -628
rect 2542 -846 2608 -692
rect 2668 -784 2728 246
rect 2788 -846 2848 186
rect 2908 -784 2968 246
rect 3028 -846 3088 186
rect 3148 92 3214 182
rect 3148 28 3149 92
rect 3213 28 3214 92
rect 3148 12 3214 28
rect 3148 -52 3149 12
rect 3213 -52 3214 12
rect 3148 -68 3214 -52
rect 3148 -132 3149 -68
rect 3213 -132 3214 -68
rect 3148 -148 3214 -132
rect 3148 -212 3149 -148
rect 3213 -212 3214 -148
rect 3148 -228 3214 -212
rect 3148 -292 3149 -228
rect 3213 -292 3214 -228
rect 3148 -308 3214 -292
rect 3148 -372 3149 -308
rect 3213 -372 3214 -308
rect 3148 -388 3214 -372
rect 3148 -452 3149 -388
rect 3213 -452 3214 -388
rect 3148 -468 3214 -452
rect 3148 -532 3149 -468
rect 3213 -532 3214 -468
rect 3148 -548 3214 -532
rect 3148 -612 3149 -548
rect 3213 -612 3214 -548
rect 3148 -628 3214 -612
rect 3148 -692 3149 -628
rect 3213 -692 3214 -628
rect 3148 -846 3214 -692
rect 3274 -846 3334 186
rect 3394 -784 3454 246
rect 3514 -846 3574 186
rect 3634 -784 3694 246
rect 3754 92 3820 182
rect 3754 28 3755 92
rect 3819 28 3820 92
rect 3754 12 3820 28
rect 3754 -52 3755 12
rect 3819 -52 3820 12
rect 3754 -68 3820 -52
rect 3754 -132 3755 -68
rect 3819 -132 3820 -68
rect 3754 -148 3820 -132
rect 3754 -212 3755 -148
rect 3819 -212 3820 -148
rect 3754 -228 3820 -212
rect 3754 -292 3755 -228
rect 3819 -292 3820 -228
rect 3754 -308 3820 -292
rect 3754 -372 3755 -308
rect 3819 -372 3820 -308
rect 3754 -388 3820 -372
rect 3754 -452 3755 -388
rect 3819 -452 3820 -388
rect 3754 -468 3820 -452
rect 3754 -532 3755 -468
rect 3819 -532 3820 -468
rect 3754 -548 3820 -532
rect 3754 -612 3755 -548
rect 3819 -612 3820 -548
rect 3754 -628 3820 -612
rect 3754 -692 3755 -628
rect 3819 -692 3820 -628
rect 3754 -846 3820 -692
rect 3880 -784 3940 246
rect 4000 -846 4060 186
rect 4120 -784 4180 246
rect 4240 -846 4300 186
rect 4360 92 4426 182
rect 4360 28 4361 92
rect 4425 28 4426 92
rect 4360 12 4426 28
rect 4360 -52 4361 12
rect 4425 -52 4426 12
rect 4360 -68 4426 -52
rect 4360 -132 4361 -68
rect 4425 -132 4426 -68
rect 4360 -148 4426 -132
rect 4360 -212 4361 -148
rect 4425 -212 4426 -148
rect 4360 -228 4426 -212
rect 4360 -292 4361 -228
rect 4425 -292 4426 -228
rect 4360 -308 4426 -292
rect 4360 -372 4361 -308
rect 4425 -372 4426 -308
rect 4360 -388 4426 -372
rect 4360 -452 4361 -388
rect 4425 -452 4426 -388
rect 4360 -468 4426 -452
rect 4360 -532 4361 -468
rect 4425 -532 4426 -468
rect 4360 -548 4426 -532
rect 4360 -612 4361 -548
rect 4425 -612 4426 -548
rect 4360 -628 4426 -612
rect 4360 -692 4361 -628
rect 4425 -692 4426 -628
rect 4360 -846 4426 -692
rect 4486 -846 4546 186
rect 4606 -784 4666 246
rect 4726 -846 4786 186
rect 4846 -784 4906 246
rect 4966 92 5032 182
rect 4966 28 4967 92
rect 5031 28 5032 92
rect 4966 12 5032 28
rect 4966 -52 4967 12
rect 5031 -52 5032 12
rect 4966 -68 5032 -52
rect 4966 -132 4967 -68
rect 5031 -132 5032 -68
rect 4966 -148 5032 -132
rect 4966 -212 4967 -148
rect 5031 -212 5032 -148
rect 4966 -228 5032 -212
rect 4966 -292 4967 -228
rect 5031 -292 5032 -228
rect 4966 -308 5032 -292
rect 4966 -372 4967 -308
rect 5031 -372 5032 -308
rect 4966 -388 5032 -372
rect 4966 -452 4967 -388
rect 5031 -452 5032 -388
rect 4966 -468 5032 -452
rect 4966 -532 4967 -468
rect 5031 -532 5032 -468
rect 4966 -548 5032 -532
rect 4966 -612 4967 -548
rect 5031 -612 5032 -548
rect 4966 -628 5032 -612
rect 4966 -692 4967 -628
rect 5031 -692 5032 -628
rect 4966 -846 5032 -692
rect 2542 -848 5032 -846
rect 2542 -912 2646 -848
rect 2710 -912 2726 -848
rect 2790 -912 2806 -848
rect 2870 -912 2886 -848
rect 2950 -912 2966 -848
rect 3030 -912 3046 -848
rect 3110 -912 3252 -848
rect 3316 -912 3332 -848
rect 3396 -912 3412 -848
rect 3476 -912 3492 -848
rect 3556 -912 3572 -848
rect 3636 -912 3652 -848
rect 3716 -912 3858 -848
rect 3922 -912 3938 -848
rect 4002 -912 4018 -848
rect 4082 -912 4098 -848
rect 4162 -912 4178 -848
rect 4242 -912 4258 -848
rect 4322 -912 4464 -848
rect 4528 -912 4544 -848
rect 4608 -912 4624 -848
rect 4688 -912 4704 -848
rect 4768 -912 4784 -848
rect 4848 -912 4864 -848
rect 4928 -912 5032 -848
rect 2542 -914 5032 -912
rect 5092 92 5158 182
rect 5092 28 5093 92
rect 5157 28 5158 92
rect 5092 12 5158 28
rect 5092 -52 5093 12
rect 5157 -52 5158 12
rect 5092 -68 5158 -52
rect 5092 -132 5093 -68
rect 5157 -132 5158 -68
rect 5092 -148 5158 -132
rect 5092 -212 5093 -148
rect 5157 -212 5158 -148
rect 5092 -228 5158 -212
rect 5092 -292 5093 -228
rect 5157 -292 5158 -228
rect 5092 -308 5158 -292
rect 5092 -372 5093 -308
rect 5157 -372 5158 -308
rect 5092 -388 5158 -372
rect 5092 -452 5093 -388
rect 5157 -452 5158 -388
rect 5092 -468 5158 -452
rect 5092 -532 5093 -468
rect 5157 -532 5158 -468
rect 5092 -548 5158 -532
rect 5092 -612 5093 -548
rect 5157 -612 5158 -548
rect 5092 -628 5158 -612
rect 5092 -692 5093 -628
rect 5157 -692 5158 -628
rect 5092 -846 5158 -692
rect 5218 -846 5278 186
rect 5338 -784 5398 246
rect 5458 -846 5518 186
rect 5578 -784 5638 246
rect 6030 240 6155 246
rect 5698 92 5764 182
rect 5698 28 5699 92
rect 5763 28 5764 92
rect 5698 12 5764 28
rect 5698 -52 5699 12
rect 5763 -52 5764 12
rect 5698 -68 5764 -52
rect 5698 -132 5699 -68
rect 5763 -132 5764 -68
rect 5698 -148 5764 -132
rect 5698 -212 5699 -148
rect 5763 -212 5764 -148
rect 5698 -228 5764 -212
rect 5698 -292 5699 -228
rect 5763 -292 5764 -228
rect 5698 -308 5764 -292
rect 5698 -372 5699 -308
rect 5763 -372 5764 -308
rect 5698 -388 5764 -372
rect 5698 -452 5699 -388
rect 5763 -452 5764 -388
rect 5698 -468 5764 -452
rect 5698 -532 5699 -468
rect 5763 -532 5764 -468
rect 5698 -548 5764 -532
rect 5698 -612 5699 -548
rect 5763 -612 5764 -548
rect 5698 -628 5764 -612
rect 5698 -692 5699 -628
rect 5763 -692 5764 -628
rect 5698 -846 5764 -692
rect 5092 -848 5764 -846
rect 5092 -912 5196 -848
rect 5260 -912 5276 -848
rect 5340 -912 5356 -848
rect 5420 -912 5436 -848
rect 5500 -912 5516 -848
rect 5580 -912 5596 -848
rect 5660 -912 5764 -848
rect 5092 -914 5764 -912
rect 214 -1076 412 -1066
rect 214 -1140 227 -1076
rect 291 -1140 412 -1076
rect 214 -1150 412 -1140
rect 472 -1097 5386 -1095
rect 472 -1161 576 -1097
rect 640 -1161 656 -1097
rect 720 -1161 736 -1097
rect 800 -1161 816 -1097
rect 880 -1161 896 -1097
rect 960 -1161 976 -1097
rect 1040 -1161 1182 -1097
rect 1246 -1161 1262 -1097
rect 1326 -1161 1342 -1097
rect 1406 -1161 1422 -1097
rect 1486 -1161 1502 -1097
rect 1566 -1161 1582 -1097
rect 1646 -1161 1788 -1097
rect 1852 -1161 1868 -1097
rect 1932 -1161 1948 -1097
rect 2012 -1161 2028 -1097
rect 2092 -1161 2108 -1097
rect 2172 -1161 2188 -1097
rect 2252 -1161 2394 -1097
rect 2458 -1161 2474 -1097
rect 2538 -1161 2554 -1097
rect 2618 -1161 2634 -1097
rect 2698 -1161 2714 -1097
rect 2778 -1161 2794 -1097
rect 2858 -1161 3000 -1097
rect 3064 -1161 3080 -1097
rect 3144 -1161 3160 -1097
rect 3224 -1161 3240 -1097
rect 3304 -1161 3320 -1097
rect 3384 -1161 3400 -1097
rect 3464 -1161 3606 -1097
rect 3670 -1161 3686 -1097
rect 3750 -1161 3766 -1097
rect 3830 -1161 3846 -1097
rect 3910 -1161 3926 -1097
rect 3990 -1161 4006 -1097
rect 4070 -1161 4212 -1097
rect 4276 -1161 4292 -1097
rect 4356 -1161 4372 -1097
rect 4436 -1161 4452 -1097
rect 4516 -1161 4532 -1097
rect 4596 -1161 4612 -1097
rect 4676 -1161 4818 -1097
rect 4882 -1161 4898 -1097
rect 4962 -1161 4978 -1097
rect 5042 -1161 5058 -1097
rect 5122 -1161 5138 -1097
rect 5202 -1161 5218 -1097
rect 5282 -1161 5386 -1097
rect 472 -1163 5386 -1161
rect 472 -1317 538 -1163
rect 94 -1337 412 -1325
rect 94 -1401 315 -1337
rect 379 -1401 412 -1337
rect 94 -2255 412 -1401
rect 472 -1381 473 -1317
rect 537 -1381 538 -1317
rect 472 -1397 538 -1381
rect 472 -1461 473 -1397
rect 537 -1461 538 -1397
rect 472 -1477 538 -1461
rect 472 -1541 473 -1477
rect 537 -1541 538 -1477
rect 472 -1557 538 -1541
rect 472 -1621 473 -1557
rect 537 -1621 538 -1557
rect 472 -1637 538 -1621
rect 472 -1701 473 -1637
rect 537 -1701 538 -1637
rect 472 -1717 538 -1701
rect 472 -1781 473 -1717
rect 537 -1781 538 -1717
rect 472 -1797 538 -1781
rect 472 -1861 473 -1797
rect 537 -1861 538 -1797
rect 472 -1877 538 -1861
rect 472 -1941 473 -1877
rect 537 -1941 538 -1877
rect 472 -1957 538 -1941
rect 472 -2021 473 -1957
rect 537 -2021 538 -1957
rect 472 -2037 538 -2021
rect 472 -2101 473 -2037
rect 537 -2101 538 -2037
rect 472 -2191 538 -2101
rect 598 -2255 658 -1225
rect 718 -2195 778 -1163
rect 838 -2255 898 -1225
rect 958 -2195 1018 -1163
rect 1078 -1317 1144 -1163
rect 1078 -1381 1079 -1317
rect 1143 -1381 1144 -1317
rect 1078 -1397 1144 -1381
rect 1078 -1461 1079 -1397
rect 1143 -1461 1144 -1397
rect 1078 -1477 1144 -1461
rect 1078 -1541 1079 -1477
rect 1143 -1541 1144 -1477
rect 1078 -1557 1144 -1541
rect 1078 -1621 1079 -1557
rect 1143 -1621 1144 -1557
rect 1078 -1637 1144 -1621
rect 1078 -1701 1079 -1637
rect 1143 -1701 1144 -1637
rect 1078 -1717 1144 -1701
rect 1078 -1781 1079 -1717
rect 1143 -1781 1144 -1717
rect 1078 -1797 1144 -1781
rect 1078 -1861 1079 -1797
rect 1143 -1861 1144 -1797
rect 1078 -1877 1144 -1861
rect 1078 -1941 1079 -1877
rect 1143 -1941 1144 -1877
rect 1078 -1957 1144 -1941
rect 1078 -2021 1079 -1957
rect 1143 -2021 1144 -1957
rect 1078 -2037 1144 -2021
rect 1078 -2101 1079 -2037
rect 1143 -2101 1144 -2037
rect 1078 -2191 1144 -2101
rect 1204 -2195 1264 -1163
rect 1324 -2255 1384 -1225
rect 1444 -2195 1504 -1163
rect 1564 -2255 1624 -1225
rect 1684 -1317 1750 -1163
rect 1684 -1381 1685 -1317
rect 1749 -1381 1750 -1317
rect 1684 -1397 1750 -1381
rect 1684 -1461 1685 -1397
rect 1749 -1461 1750 -1397
rect 1684 -1477 1750 -1461
rect 1684 -1541 1685 -1477
rect 1749 -1541 1750 -1477
rect 1684 -1557 1750 -1541
rect 1684 -1621 1685 -1557
rect 1749 -1621 1750 -1557
rect 1684 -1637 1750 -1621
rect 1684 -1701 1685 -1637
rect 1749 -1701 1750 -1637
rect 1684 -1717 1750 -1701
rect 1684 -1781 1685 -1717
rect 1749 -1781 1750 -1717
rect 1684 -1797 1750 -1781
rect 1684 -1861 1685 -1797
rect 1749 -1861 1750 -1797
rect 1684 -1877 1750 -1861
rect 1684 -1941 1685 -1877
rect 1749 -1941 1750 -1877
rect 1684 -1957 1750 -1941
rect 1684 -2021 1685 -1957
rect 1749 -2021 1750 -1957
rect 1684 -2037 1750 -2021
rect 1684 -2101 1685 -2037
rect 1749 -2101 1750 -2037
rect 1684 -2191 1750 -2101
rect 1810 -2255 1870 -1225
rect 1930 -2195 1990 -1163
rect 2050 -2255 2110 -1225
rect 2170 -2195 2230 -1163
rect 2290 -1317 2356 -1163
rect 2290 -1381 2291 -1317
rect 2355 -1381 2356 -1317
rect 2290 -1397 2356 -1381
rect 2290 -1461 2291 -1397
rect 2355 -1461 2356 -1397
rect 2290 -1477 2356 -1461
rect 2290 -1541 2291 -1477
rect 2355 -1541 2356 -1477
rect 2290 -1557 2356 -1541
rect 2290 -1621 2291 -1557
rect 2355 -1621 2356 -1557
rect 2290 -1637 2356 -1621
rect 2290 -1701 2291 -1637
rect 2355 -1701 2356 -1637
rect 2290 -1717 2356 -1701
rect 2290 -1781 2291 -1717
rect 2355 -1781 2356 -1717
rect 2290 -1797 2356 -1781
rect 2290 -1861 2291 -1797
rect 2355 -1861 2356 -1797
rect 2290 -1877 2356 -1861
rect 2290 -1941 2291 -1877
rect 2355 -1941 2356 -1877
rect 2290 -1957 2356 -1941
rect 2290 -2021 2291 -1957
rect 2355 -2021 2356 -1957
rect 2290 -2037 2356 -2021
rect 2290 -2101 2291 -2037
rect 2355 -2101 2356 -2037
rect 2290 -2191 2356 -2101
rect 2416 -2195 2476 -1163
rect 2536 -2255 2596 -1225
rect 2656 -2195 2716 -1163
rect 2776 -2255 2836 -1225
rect 2896 -1317 2962 -1163
rect 2896 -1381 2897 -1317
rect 2961 -1381 2962 -1317
rect 2896 -1397 2962 -1381
rect 2896 -1461 2897 -1397
rect 2961 -1461 2962 -1397
rect 2896 -1477 2962 -1461
rect 2896 -1541 2897 -1477
rect 2961 -1541 2962 -1477
rect 2896 -1557 2962 -1541
rect 2896 -1621 2897 -1557
rect 2961 -1621 2962 -1557
rect 2896 -1637 2962 -1621
rect 2896 -1701 2897 -1637
rect 2961 -1701 2962 -1637
rect 2896 -1717 2962 -1701
rect 2896 -1781 2897 -1717
rect 2961 -1781 2962 -1717
rect 2896 -1797 2962 -1781
rect 2896 -1861 2897 -1797
rect 2961 -1861 2962 -1797
rect 2896 -1877 2962 -1861
rect 2896 -1941 2897 -1877
rect 2961 -1941 2962 -1877
rect 2896 -1957 2962 -1941
rect 2896 -2021 2897 -1957
rect 2961 -2021 2962 -1957
rect 2896 -2037 2962 -2021
rect 2896 -2101 2897 -2037
rect 2961 -2101 2962 -2037
rect 2896 -2191 2962 -2101
rect 3022 -2255 3082 -1225
rect 3142 -2195 3202 -1163
rect 3262 -2255 3322 -1225
rect 3382 -2195 3442 -1163
rect 3502 -1317 3568 -1163
rect 3502 -1381 3503 -1317
rect 3567 -1381 3568 -1317
rect 3502 -1397 3568 -1381
rect 3502 -1461 3503 -1397
rect 3567 -1461 3568 -1397
rect 3502 -1477 3568 -1461
rect 3502 -1541 3503 -1477
rect 3567 -1541 3568 -1477
rect 3502 -1557 3568 -1541
rect 3502 -1621 3503 -1557
rect 3567 -1621 3568 -1557
rect 3502 -1637 3568 -1621
rect 3502 -1701 3503 -1637
rect 3567 -1701 3568 -1637
rect 3502 -1717 3568 -1701
rect 3502 -1781 3503 -1717
rect 3567 -1781 3568 -1717
rect 3502 -1797 3568 -1781
rect 3502 -1861 3503 -1797
rect 3567 -1861 3568 -1797
rect 3502 -1877 3568 -1861
rect 3502 -1941 3503 -1877
rect 3567 -1941 3568 -1877
rect 3502 -1957 3568 -1941
rect 3502 -2021 3503 -1957
rect 3567 -2021 3568 -1957
rect 3502 -2037 3568 -2021
rect 3502 -2101 3503 -2037
rect 3567 -2101 3568 -2037
rect 3502 -2191 3568 -2101
rect 3628 -2195 3688 -1163
rect 3748 -2255 3808 -1225
rect 3868 -2195 3928 -1163
rect 3988 -2255 4048 -1225
rect 4108 -1317 4174 -1163
rect 4108 -1381 4109 -1317
rect 4173 -1381 4174 -1317
rect 4108 -1397 4174 -1381
rect 4108 -1461 4109 -1397
rect 4173 -1461 4174 -1397
rect 4108 -1477 4174 -1461
rect 4108 -1541 4109 -1477
rect 4173 -1541 4174 -1477
rect 4108 -1557 4174 -1541
rect 4108 -1621 4109 -1557
rect 4173 -1621 4174 -1557
rect 4108 -1637 4174 -1621
rect 4108 -1701 4109 -1637
rect 4173 -1701 4174 -1637
rect 4108 -1717 4174 -1701
rect 4108 -1781 4109 -1717
rect 4173 -1781 4174 -1717
rect 4108 -1797 4174 -1781
rect 4108 -1861 4109 -1797
rect 4173 -1861 4174 -1797
rect 4108 -1877 4174 -1861
rect 4108 -1941 4109 -1877
rect 4173 -1941 4174 -1877
rect 4108 -1957 4174 -1941
rect 4108 -2021 4109 -1957
rect 4173 -2021 4174 -1957
rect 4108 -2037 4174 -2021
rect 4108 -2101 4109 -2037
rect 4173 -2101 4174 -2037
rect 4108 -2191 4174 -2101
rect 4234 -2255 4294 -1225
rect 4354 -2195 4414 -1163
rect 4474 -2255 4534 -1225
rect 4594 -2195 4654 -1163
rect 4714 -1317 4780 -1163
rect 4714 -1381 4715 -1317
rect 4779 -1381 4780 -1317
rect 4714 -1397 4780 -1381
rect 4714 -1461 4715 -1397
rect 4779 -1461 4780 -1397
rect 4714 -1477 4780 -1461
rect 4714 -1541 4715 -1477
rect 4779 -1541 4780 -1477
rect 4714 -1557 4780 -1541
rect 4714 -1621 4715 -1557
rect 4779 -1621 4780 -1557
rect 4714 -1637 4780 -1621
rect 4714 -1701 4715 -1637
rect 4779 -1701 4780 -1637
rect 4714 -1717 4780 -1701
rect 4714 -1781 4715 -1717
rect 4779 -1781 4780 -1717
rect 4714 -1797 4780 -1781
rect 4714 -1861 4715 -1797
rect 4779 -1861 4780 -1797
rect 4714 -1877 4780 -1861
rect 4714 -1941 4715 -1877
rect 4779 -1941 4780 -1877
rect 4714 -1957 4780 -1941
rect 4714 -2021 4715 -1957
rect 4779 -2021 4780 -1957
rect 4714 -2037 4780 -2021
rect 4714 -2101 4715 -2037
rect 4779 -2101 4780 -2037
rect 4714 -2191 4780 -2101
rect 4840 -2195 4900 -1163
rect 4960 -2255 5020 -1225
rect 5080 -2195 5140 -1163
rect 5200 -2255 5260 -1225
rect 5320 -1317 5386 -1163
rect 5320 -1381 5321 -1317
rect 5385 -1381 5386 -1317
rect 5320 -1397 5386 -1381
rect 5320 -1461 5321 -1397
rect 5385 -1461 5386 -1397
rect 5320 -1477 5386 -1461
rect 5320 -1541 5321 -1477
rect 5385 -1541 5386 -1477
rect 5320 -1557 5386 -1541
rect 5320 -1621 5321 -1557
rect 5385 -1621 5386 -1557
rect 5320 -1637 5386 -1621
rect 5320 -1701 5321 -1637
rect 5385 -1701 5386 -1637
rect 5320 -1717 5386 -1701
rect 5320 -1781 5321 -1717
rect 5385 -1781 5386 -1717
rect 5320 -1797 5386 -1781
rect 5320 -1861 5321 -1797
rect 5385 -1861 5386 -1797
rect 5320 -1877 5386 -1861
rect 5320 -1941 5321 -1877
rect 5385 -1941 5386 -1877
rect 5320 -1957 5386 -1941
rect 5320 -2021 5321 -1957
rect 5385 -2021 5386 -1957
rect 5320 -2037 5386 -2021
rect 5320 -2101 5321 -2037
rect 5385 -2101 5386 -2037
rect 5320 -2191 5386 -2101
rect 5446 -1097 6118 -1095
rect 5446 -1161 5550 -1097
rect 5614 -1161 5630 -1097
rect 5694 -1161 5710 -1097
rect 5774 -1161 5790 -1097
rect 5854 -1161 5870 -1097
rect 5934 -1161 5950 -1097
rect 6014 -1161 6118 -1097
rect 5446 -1163 6118 -1161
rect 5446 -1317 5512 -1163
rect 5446 -1381 5447 -1317
rect 5511 -1381 5512 -1317
rect 5446 -1397 5512 -1381
rect 5446 -1461 5447 -1397
rect 5511 -1461 5512 -1397
rect 5446 -1477 5512 -1461
rect 5446 -1541 5447 -1477
rect 5511 -1541 5512 -1477
rect 5446 -1557 5512 -1541
rect 5446 -1621 5447 -1557
rect 5511 -1621 5512 -1557
rect 5446 -1637 5512 -1621
rect 5446 -1701 5447 -1637
rect 5511 -1701 5512 -1637
rect 5446 -1717 5512 -1701
rect 5446 -1781 5447 -1717
rect 5511 -1781 5512 -1717
rect 5446 -1797 5512 -1781
rect 5446 -1861 5447 -1797
rect 5511 -1861 5512 -1797
rect 5446 -1877 5512 -1861
rect 5446 -1941 5447 -1877
rect 5511 -1941 5512 -1877
rect 5446 -1957 5512 -1941
rect 5446 -2021 5447 -1957
rect 5511 -2021 5512 -1957
rect 5446 -2037 5512 -2021
rect 5446 -2101 5447 -2037
rect 5511 -2101 5512 -2037
rect 5446 -2191 5512 -2101
rect 5572 -2195 5632 -1163
rect 5692 -2255 5752 -1225
rect 5812 -2195 5872 -1163
rect 5932 -2255 5992 -1225
rect 6052 -1317 6118 -1163
rect 6340 -1098 6770 246
rect 6849 -611 7167 246
rect 6849 -675 7073 -611
rect 7137 -675 7167 -611
rect 6849 -685 7167 -675
rect 6849 -873 7047 -863
rect 6849 -937 6982 -873
rect 7046 -937 7047 -873
rect 6849 -947 7047 -937
rect 6340 -1113 6771 -1098
rect 6340 -1177 6383 -1113
rect 6447 -1177 6526 -1113
rect 6590 -1177 6646 -1113
rect 6710 -1177 6771 -1113
rect 6340 -1192 6771 -1177
rect 6052 -1381 6053 -1317
rect 6117 -1381 6118 -1317
rect 6052 -1397 6118 -1381
rect 6052 -1461 6053 -1397
rect 6117 -1461 6118 -1397
rect 6052 -1477 6118 -1461
rect 6052 -1541 6053 -1477
rect 6117 -1541 6118 -1477
rect 6052 -1557 6118 -1541
rect 6052 -1621 6053 -1557
rect 6117 -1621 6118 -1557
rect 6052 -1637 6118 -1621
rect 6052 -1701 6053 -1637
rect 6117 -1701 6118 -1637
rect 6849 -1325 6909 -947
rect 7107 -1066 7167 -685
rect 7227 92 7293 182
rect 7227 28 7228 92
rect 7292 28 7293 92
rect 7227 12 7293 28
rect 7227 -52 7228 12
rect 7292 -52 7293 12
rect 7227 -68 7293 -52
rect 7227 -132 7228 -68
rect 7292 -132 7293 -68
rect 7227 -148 7293 -132
rect 7227 -212 7228 -148
rect 7292 -212 7293 -148
rect 7227 -228 7293 -212
rect 7227 -292 7228 -228
rect 7292 -292 7293 -228
rect 7227 -308 7293 -292
rect 7227 -372 7228 -308
rect 7292 -372 7293 -308
rect 7227 -388 7293 -372
rect 7227 -452 7228 -388
rect 7292 -452 7293 -388
rect 7227 -468 7293 -452
rect 7227 -532 7228 -468
rect 7292 -532 7293 -468
rect 7227 -548 7293 -532
rect 7227 -612 7228 -548
rect 7292 -612 7293 -548
rect 7227 -628 7293 -612
rect 7227 -692 7228 -628
rect 7292 -692 7293 -628
rect 7227 -846 7293 -692
rect 7353 -784 7413 246
rect 7473 -846 7533 186
rect 7593 -784 7653 246
rect 7713 -846 7773 186
rect 7833 92 7899 182
rect 7833 28 7834 92
rect 7898 28 7899 92
rect 7833 12 7899 28
rect 7833 -52 7834 12
rect 7898 -52 7899 12
rect 7833 -68 7899 -52
rect 7833 -132 7834 -68
rect 7898 -132 7899 -68
rect 7833 -148 7899 -132
rect 7833 -212 7834 -148
rect 7898 -212 7899 -148
rect 7833 -228 7899 -212
rect 7833 -292 7834 -228
rect 7898 -292 7899 -228
rect 7833 -308 7899 -292
rect 7833 -372 7834 -308
rect 7898 -372 7899 -308
rect 7833 -388 7899 -372
rect 7833 -452 7834 -388
rect 7898 -452 7899 -388
rect 7833 -468 7899 -452
rect 7833 -532 7834 -468
rect 7898 -532 7899 -468
rect 7833 -548 7899 -532
rect 7833 -612 7834 -548
rect 7898 -612 7899 -548
rect 7833 -628 7899 -612
rect 7833 -692 7834 -628
rect 7898 -692 7899 -628
rect 7833 -846 7899 -692
rect 7227 -848 7899 -846
rect 7227 -912 7331 -848
rect 7395 -912 7411 -848
rect 7475 -912 7491 -848
rect 7555 -912 7571 -848
rect 7635 -912 7651 -848
rect 7715 -912 7731 -848
rect 7795 -912 7899 -848
rect 7227 -914 7899 -912
rect 7959 92 8025 182
rect 7959 28 7960 92
rect 8024 28 8025 92
rect 7959 12 8025 28
rect 7959 -52 7960 12
rect 8024 -52 8025 12
rect 7959 -68 8025 -52
rect 7959 -132 7960 -68
rect 8024 -132 8025 -68
rect 7959 -148 8025 -132
rect 7959 -212 7960 -148
rect 8024 -212 8025 -148
rect 7959 -228 8025 -212
rect 7959 -292 7960 -228
rect 8024 -292 8025 -228
rect 7959 -308 8025 -292
rect 7959 -372 7960 -308
rect 8024 -372 8025 -308
rect 7959 -388 8025 -372
rect 7959 -452 7960 -388
rect 8024 -452 8025 -388
rect 7959 -468 8025 -452
rect 7959 -532 7960 -468
rect 8024 -532 8025 -468
rect 7959 -548 8025 -532
rect 7959 -612 7960 -548
rect 8024 -612 8025 -548
rect 7959 -628 8025 -612
rect 7959 -692 7960 -628
rect 8024 -692 8025 -628
rect 7959 -846 8025 -692
rect 8085 -784 8145 246
rect 8205 -846 8265 186
rect 8325 -784 8385 246
rect 8445 -846 8505 186
rect 8565 92 8631 182
rect 8565 28 8566 92
rect 8630 28 8631 92
rect 8565 12 8631 28
rect 8565 -52 8566 12
rect 8630 -52 8631 12
rect 8565 -68 8631 -52
rect 8565 -132 8566 -68
rect 8630 -132 8631 -68
rect 8565 -148 8631 -132
rect 8565 -212 8566 -148
rect 8630 -212 8631 -148
rect 8565 -228 8631 -212
rect 8565 -292 8566 -228
rect 8630 -292 8631 -228
rect 8565 -308 8631 -292
rect 8565 -372 8566 -308
rect 8630 -372 8631 -308
rect 8565 -388 8631 -372
rect 8565 -452 8566 -388
rect 8630 -452 8631 -388
rect 8565 -468 8631 -452
rect 8565 -532 8566 -468
rect 8630 -532 8631 -468
rect 8565 -548 8631 -532
rect 8565 -612 8566 -548
rect 8630 -612 8631 -548
rect 8565 -628 8631 -612
rect 8565 -692 8566 -628
rect 8630 -692 8631 -628
rect 8565 -846 8631 -692
rect 8691 -846 8751 186
rect 8811 -784 8871 246
rect 8931 -846 8991 186
rect 9051 -784 9111 246
rect 9171 92 9237 182
rect 9171 28 9172 92
rect 9236 28 9237 92
rect 9171 12 9237 28
rect 9171 -52 9172 12
rect 9236 -52 9237 12
rect 9171 -68 9237 -52
rect 9171 -132 9172 -68
rect 9236 -132 9237 -68
rect 9171 -148 9237 -132
rect 9171 -212 9172 -148
rect 9236 -212 9237 -148
rect 9171 -228 9237 -212
rect 9171 -292 9172 -228
rect 9236 -292 9237 -228
rect 9171 -308 9237 -292
rect 9171 -372 9172 -308
rect 9236 -372 9237 -308
rect 9171 -388 9237 -372
rect 9171 -452 9172 -388
rect 9236 -452 9237 -388
rect 9171 -468 9237 -452
rect 9171 -532 9172 -468
rect 9236 -532 9237 -468
rect 9171 -548 9237 -532
rect 9171 -612 9172 -548
rect 9236 -612 9237 -548
rect 9171 -628 9237 -612
rect 9171 -692 9172 -628
rect 9236 -692 9237 -628
rect 9171 -846 9237 -692
rect 7959 -848 9237 -846
rect 7959 -912 8063 -848
rect 8127 -912 8143 -848
rect 8207 -912 8223 -848
rect 8287 -912 8303 -848
rect 8367 -912 8383 -848
rect 8447 -912 8463 -848
rect 8527 -912 8669 -848
rect 8733 -912 8749 -848
rect 8813 -912 8829 -848
rect 8893 -912 8909 -848
rect 8973 -912 8989 -848
rect 9053 -912 9069 -848
rect 9133 -912 9237 -848
rect 7959 -914 9237 -912
rect 9297 92 9363 182
rect 9297 28 9298 92
rect 9362 28 9363 92
rect 9297 12 9363 28
rect 9297 -52 9298 12
rect 9362 -52 9363 12
rect 9297 -68 9363 -52
rect 9297 -132 9298 -68
rect 9362 -132 9363 -68
rect 9297 -148 9363 -132
rect 9297 -212 9298 -148
rect 9362 -212 9363 -148
rect 9297 -228 9363 -212
rect 9297 -292 9298 -228
rect 9362 -292 9363 -228
rect 9297 -308 9363 -292
rect 9297 -372 9298 -308
rect 9362 -372 9363 -308
rect 9297 -388 9363 -372
rect 9297 -452 9298 -388
rect 9362 -452 9363 -388
rect 9297 -468 9363 -452
rect 9297 -532 9298 -468
rect 9362 -532 9363 -468
rect 9297 -548 9363 -532
rect 9297 -612 9298 -548
rect 9362 -612 9363 -548
rect 9297 -628 9363 -612
rect 9297 -692 9298 -628
rect 9362 -692 9363 -628
rect 9297 -846 9363 -692
rect 9423 -784 9483 246
rect 9543 -846 9603 186
rect 9663 -784 9723 246
rect 9783 -846 9843 186
rect 9903 92 9969 182
rect 9903 28 9904 92
rect 9968 28 9969 92
rect 9903 12 9969 28
rect 9903 -52 9904 12
rect 9968 -52 9969 12
rect 9903 -68 9969 -52
rect 9903 -132 9904 -68
rect 9968 -132 9969 -68
rect 9903 -148 9969 -132
rect 9903 -212 9904 -148
rect 9968 -212 9969 -148
rect 9903 -228 9969 -212
rect 9903 -292 9904 -228
rect 9968 -292 9969 -228
rect 9903 -308 9969 -292
rect 9903 -372 9904 -308
rect 9968 -372 9969 -308
rect 9903 -388 9969 -372
rect 9903 -452 9904 -388
rect 9968 -452 9969 -388
rect 9903 -468 9969 -452
rect 9903 -532 9904 -468
rect 9968 -532 9969 -468
rect 9903 -548 9969 -532
rect 9903 -612 9904 -548
rect 9968 -612 9969 -548
rect 9903 -628 9969 -612
rect 9903 -692 9904 -628
rect 9968 -692 9969 -628
rect 9903 -846 9969 -692
rect 10029 -846 10089 186
rect 10149 -784 10209 246
rect 10269 -846 10329 186
rect 10389 -784 10449 246
rect 10509 92 10575 182
rect 10509 28 10510 92
rect 10574 28 10575 92
rect 10509 12 10575 28
rect 10509 -52 10510 12
rect 10574 -52 10575 12
rect 10509 -68 10575 -52
rect 10509 -132 10510 -68
rect 10574 -132 10575 -68
rect 10509 -148 10575 -132
rect 10509 -212 10510 -148
rect 10574 -212 10575 -148
rect 10509 -228 10575 -212
rect 10509 -292 10510 -228
rect 10574 -292 10575 -228
rect 10509 -308 10575 -292
rect 10509 -372 10510 -308
rect 10574 -372 10575 -308
rect 10509 -388 10575 -372
rect 10509 -452 10510 -388
rect 10574 -452 10575 -388
rect 10509 -468 10575 -452
rect 10509 -532 10510 -468
rect 10574 -532 10575 -468
rect 10509 -548 10575 -532
rect 10509 -612 10510 -548
rect 10574 -612 10575 -548
rect 10509 -628 10575 -612
rect 10509 -692 10510 -628
rect 10574 -692 10575 -628
rect 10509 -846 10575 -692
rect 10635 -784 10695 246
rect 10755 -846 10815 186
rect 10875 -784 10935 246
rect 10995 -846 11055 186
rect 11115 92 11181 182
rect 11115 28 11116 92
rect 11180 28 11181 92
rect 11115 12 11181 28
rect 11115 -52 11116 12
rect 11180 -52 11181 12
rect 11115 -68 11181 -52
rect 11115 -132 11116 -68
rect 11180 -132 11181 -68
rect 11115 -148 11181 -132
rect 11115 -212 11116 -148
rect 11180 -212 11181 -148
rect 11115 -228 11181 -212
rect 11115 -292 11116 -228
rect 11180 -292 11181 -228
rect 11115 -308 11181 -292
rect 11115 -372 11116 -308
rect 11180 -372 11181 -308
rect 11115 -388 11181 -372
rect 11115 -452 11116 -388
rect 11180 -452 11181 -388
rect 11115 -468 11181 -452
rect 11115 -532 11116 -468
rect 11180 -532 11181 -468
rect 11115 -548 11181 -532
rect 11115 -612 11116 -548
rect 11180 -612 11181 -548
rect 11115 -628 11181 -612
rect 11115 -692 11116 -628
rect 11180 -692 11181 -628
rect 11115 -846 11181 -692
rect 11241 -846 11301 186
rect 11361 -784 11421 246
rect 11481 -846 11541 186
rect 11601 -784 11661 246
rect 11721 92 11787 182
rect 11721 28 11722 92
rect 11786 28 11787 92
rect 11721 12 11787 28
rect 11721 -52 11722 12
rect 11786 -52 11787 12
rect 11721 -68 11787 -52
rect 11721 -132 11722 -68
rect 11786 -132 11787 -68
rect 11721 -148 11787 -132
rect 11721 -212 11722 -148
rect 11786 -212 11787 -148
rect 11721 -228 11787 -212
rect 11721 -292 11722 -228
rect 11786 -292 11787 -228
rect 11721 -308 11787 -292
rect 11721 -372 11722 -308
rect 11786 -372 11787 -308
rect 11721 -388 11787 -372
rect 11721 -452 11722 -388
rect 11786 -452 11787 -388
rect 11721 -468 11787 -452
rect 11721 -532 11722 -468
rect 11786 -532 11787 -468
rect 11721 -548 11787 -532
rect 11721 -612 11722 -548
rect 11786 -612 11787 -548
rect 11721 -628 11787 -612
rect 11721 -692 11722 -628
rect 11786 -692 11787 -628
rect 11721 -846 11787 -692
rect 9297 -848 11787 -846
rect 9297 -912 9401 -848
rect 9465 -912 9481 -848
rect 9545 -912 9561 -848
rect 9625 -912 9641 -848
rect 9705 -912 9721 -848
rect 9785 -912 9801 -848
rect 9865 -912 10007 -848
rect 10071 -912 10087 -848
rect 10151 -912 10167 -848
rect 10231 -912 10247 -848
rect 10311 -912 10327 -848
rect 10391 -912 10407 -848
rect 10471 -912 10613 -848
rect 10677 -912 10693 -848
rect 10757 -912 10773 -848
rect 10837 -912 10853 -848
rect 10917 -912 10933 -848
rect 10997 -912 11013 -848
rect 11077 -912 11219 -848
rect 11283 -912 11299 -848
rect 11363 -912 11379 -848
rect 11443 -912 11459 -848
rect 11523 -912 11539 -848
rect 11603 -912 11619 -848
rect 11683 -912 11787 -848
rect 9297 -914 11787 -912
rect 11847 92 11913 182
rect 11847 28 11848 92
rect 11912 28 11913 92
rect 11847 12 11913 28
rect 11847 -52 11848 12
rect 11912 -52 11913 12
rect 11847 -68 11913 -52
rect 11847 -132 11848 -68
rect 11912 -132 11913 -68
rect 11847 -148 11913 -132
rect 11847 -212 11848 -148
rect 11912 -212 11913 -148
rect 11847 -228 11913 -212
rect 11847 -292 11848 -228
rect 11912 -292 11913 -228
rect 11847 -308 11913 -292
rect 11847 -372 11848 -308
rect 11912 -372 11913 -308
rect 11847 -388 11913 -372
rect 11847 -452 11848 -388
rect 11912 -452 11913 -388
rect 11847 -468 11913 -452
rect 11847 -532 11848 -468
rect 11912 -532 11913 -468
rect 11847 -548 11913 -532
rect 11847 -612 11848 -548
rect 11912 -612 11913 -548
rect 11847 -628 11913 -612
rect 11847 -692 11848 -628
rect 11912 -692 11913 -628
rect 11847 -846 11913 -692
rect 11973 -846 12033 186
rect 12093 -784 12153 246
rect 12213 -846 12273 186
rect 12333 -784 12393 246
rect 12785 240 12910 246
rect 12453 92 12519 182
rect 12453 28 12454 92
rect 12518 28 12519 92
rect 12453 12 12519 28
rect 12453 -52 12454 12
rect 12518 -52 12519 12
rect 12453 -68 12519 -52
rect 12453 -132 12454 -68
rect 12518 -132 12519 -68
rect 12453 -148 12519 -132
rect 12453 -212 12454 -148
rect 12518 -212 12519 -148
rect 12453 -228 12519 -212
rect 12453 -292 12454 -228
rect 12518 -292 12519 -228
rect 12453 -308 12519 -292
rect 12453 -372 12454 -308
rect 12518 -372 12519 -308
rect 12453 -388 12519 -372
rect 12453 -452 12454 -388
rect 12518 -452 12519 -388
rect 12453 -468 12519 -452
rect 12453 -532 12454 -468
rect 12518 -532 12519 -468
rect 12453 -548 12519 -532
rect 12453 -612 12454 -548
rect 12518 -612 12519 -548
rect 12453 -628 12519 -612
rect 12453 -692 12454 -628
rect 12518 -692 12519 -628
rect 12453 -846 12519 -692
rect 11847 -848 12519 -846
rect 11847 -912 11951 -848
rect 12015 -912 12031 -848
rect 12095 -912 12111 -848
rect 12175 -912 12191 -848
rect 12255 -912 12271 -848
rect 12335 -912 12351 -848
rect 12415 -912 12519 -848
rect 11847 -914 12519 -912
rect 6969 -1076 7167 -1066
rect 6969 -1140 6982 -1076
rect 7046 -1140 7167 -1076
rect 6969 -1150 7167 -1140
rect 7227 -1097 12141 -1095
rect 7227 -1161 7331 -1097
rect 7395 -1161 7411 -1097
rect 7475 -1161 7491 -1097
rect 7555 -1161 7571 -1097
rect 7635 -1161 7651 -1097
rect 7715 -1161 7731 -1097
rect 7795 -1161 7937 -1097
rect 8001 -1161 8017 -1097
rect 8081 -1161 8097 -1097
rect 8161 -1161 8177 -1097
rect 8241 -1161 8257 -1097
rect 8321 -1161 8337 -1097
rect 8401 -1161 8543 -1097
rect 8607 -1161 8623 -1097
rect 8687 -1161 8703 -1097
rect 8767 -1161 8783 -1097
rect 8847 -1161 8863 -1097
rect 8927 -1161 8943 -1097
rect 9007 -1161 9149 -1097
rect 9213 -1161 9229 -1097
rect 9293 -1161 9309 -1097
rect 9373 -1161 9389 -1097
rect 9453 -1161 9469 -1097
rect 9533 -1161 9549 -1097
rect 9613 -1161 9755 -1097
rect 9819 -1161 9835 -1097
rect 9899 -1161 9915 -1097
rect 9979 -1161 9995 -1097
rect 10059 -1161 10075 -1097
rect 10139 -1161 10155 -1097
rect 10219 -1161 10361 -1097
rect 10425 -1161 10441 -1097
rect 10505 -1161 10521 -1097
rect 10585 -1161 10601 -1097
rect 10665 -1161 10681 -1097
rect 10745 -1161 10761 -1097
rect 10825 -1161 10967 -1097
rect 11031 -1161 11047 -1097
rect 11111 -1161 11127 -1097
rect 11191 -1161 11207 -1097
rect 11271 -1161 11287 -1097
rect 11351 -1161 11367 -1097
rect 11431 -1161 11573 -1097
rect 11637 -1161 11653 -1097
rect 11717 -1161 11733 -1097
rect 11797 -1161 11813 -1097
rect 11877 -1161 11893 -1097
rect 11957 -1161 11973 -1097
rect 12037 -1161 12141 -1097
rect 7227 -1163 12141 -1161
rect 7227 -1317 7293 -1163
rect 6849 -1337 7167 -1325
rect 6849 -1401 7070 -1337
rect 7134 -1401 7167 -1337
rect 6052 -1717 6118 -1701
rect 6052 -1781 6053 -1717
rect 6117 -1781 6118 -1717
rect 6052 -1797 6118 -1781
rect 6052 -1861 6053 -1797
rect 6117 -1861 6118 -1797
rect 6052 -1877 6118 -1861
rect 6052 -1941 6053 -1877
rect 6117 -1941 6118 -1877
rect 6052 -1957 6118 -1941
rect 6052 -2021 6053 -1957
rect 6117 -2021 6118 -1957
rect 6052 -2037 6118 -2021
rect 6052 -2101 6053 -2037
rect 6117 -2101 6118 -2037
rect 6052 -2191 6118 -2101
rect 6326 -1658 6788 -1640
rect 6326 -1659 6533 -1658
rect 6326 -1723 6389 -1659
rect 6453 -1722 6533 -1659
rect 6597 -1659 6788 -1658
rect 6597 -1722 6664 -1659
rect 6453 -1723 6664 -1722
rect 6728 -1723 6788 -1659
rect 6326 -2255 6788 -1723
rect 94 -2257 6788 -2255
rect 94 -2321 576 -2257
rect 640 -2321 656 -2257
rect 720 -2321 736 -2257
rect 800 -2321 816 -2257
rect 880 -2321 896 -2257
rect 960 -2321 976 -2257
rect 1040 -2321 1182 -2257
rect 1246 -2321 1262 -2257
rect 1326 -2321 1342 -2257
rect 1406 -2321 1422 -2257
rect 1486 -2321 1502 -2257
rect 1566 -2321 1582 -2257
rect 1646 -2321 1788 -2257
rect 1852 -2321 1868 -2257
rect 1932 -2321 1948 -2257
rect 2012 -2321 2028 -2257
rect 2092 -2321 2108 -2257
rect 2172 -2321 2188 -2257
rect 2252 -2321 2394 -2257
rect 2458 -2321 2474 -2257
rect 2538 -2321 2554 -2257
rect 2618 -2321 2634 -2257
rect 2698 -2321 2714 -2257
rect 2778 -2321 2794 -2257
rect 2858 -2321 3000 -2257
rect 3064 -2321 3080 -2257
rect 3144 -2321 3160 -2257
rect 3224 -2321 3240 -2257
rect 3304 -2321 3320 -2257
rect 3384 -2321 3400 -2257
rect 3464 -2321 3606 -2257
rect 3670 -2321 3686 -2257
rect 3750 -2321 3766 -2257
rect 3830 -2321 3846 -2257
rect 3910 -2321 3926 -2257
rect 3990 -2321 4006 -2257
rect 4070 -2321 4212 -2257
rect 4276 -2321 4292 -2257
rect 4356 -2321 4372 -2257
rect 4436 -2321 4452 -2257
rect 4516 -2321 4532 -2257
rect 4596 -2321 4612 -2257
rect 4676 -2321 4818 -2257
rect 4882 -2321 4898 -2257
rect 4962 -2321 4978 -2257
rect 5042 -2321 5058 -2257
rect 5122 -2321 5138 -2257
rect 5202 -2321 5218 -2257
rect 5282 -2321 5550 -2257
rect 5614 -2321 5630 -2257
rect 5694 -2321 5710 -2257
rect 5774 -2321 5790 -2257
rect 5854 -2321 5870 -2257
rect 5934 -2321 5950 -2257
rect 6014 -2264 6788 -2257
rect 6014 -2321 6047 -2264
rect 94 -2328 6047 -2321
rect 6111 -2328 6788 -2264
rect 94 -2333 6788 -2328
rect 6849 -2255 7167 -1401
rect 7227 -1381 7228 -1317
rect 7292 -1381 7293 -1317
rect 7227 -1397 7293 -1381
rect 7227 -1461 7228 -1397
rect 7292 -1461 7293 -1397
rect 7227 -1477 7293 -1461
rect 7227 -1541 7228 -1477
rect 7292 -1541 7293 -1477
rect 7227 -1557 7293 -1541
rect 7227 -1621 7228 -1557
rect 7292 -1621 7293 -1557
rect 7227 -1637 7293 -1621
rect 7227 -1701 7228 -1637
rect 7292 -1701 7293 -1637
rect 7227 -1717 7293 -1701
rect 7227 -1781 7228 -1717
rect 7292 -1781 7293 -1717
rect 7227 -1797 7293 -1781
rect 7227 -1861 7228 -1797
rect 7292 -1861 7293 -1797
rect 7227 -1877 7293 -1861
rect 7227 -1941 7228 -1877
rect 7292 -1941 7293 -1877
rect 7227 -1957 7293 -1941
rect 7227 -2021 7228 -1957
rect 7292 -2021 7293 -1957
rect 7227 -2037 7293 -2021
rect 7227 -2101 7228 -2037
rect 7292 -2101 7293 -2037
rect 7227 -2191 7293 -2101
rect 7353 -2255 7413 -1225
rect 7473 -2195 7533 -1163
rect 7593 -2255 7653 -1225
rect 7713 -2195 7773 -1163
rect 7833 -1317 7899 -1163
rect 7833 -1381 7834 -1317
rect 7898 -1381 7899 -1317
rect 7833 -1397 7899 -1381
rect 7833 -1461 7834 -1397
rect 7898 -1461 7899 -1397
rect 7833 -1477 7899 -1461
rect 7833 -1541 7834 -1477
rect 7898 -1541 7899 -1477
rect 7833 -1557 7899 -1541
rect 7833 -1621 7834 -1557
rect 7898 -1621 7899 -1557
rect 7833 -1637 7899 -1621
rect 7833 -1701 7834 -1637
rect 7898 -1701 7899 -1637
rect 7833 -1717 7899 -1701
rect 7833 -1781 7834 -1717
rect 7898 -1781 7899 -1717
rect 7833 -1797 7899 -1781
rect 7833 -1861 7834 -1797
rect 7898 -1861 7899 -1797
rect 7833 -1877 7899 -1861
rect 7833 -1941 7834 -1877
rect 7898 -1941 7899 -1877
rect 7833 -1957 7899 -1941
rect 7833 -2021 7834 -1957
rect 7898 -2021 7899 -1957
rect 7833 -2037 7899 -2021
rect 7833 -2101 7834 -2037
rect 7898 -2101 7899 -2037
rect 7833 -2191 7899 -2101
rect 7959 -2195 8019 -1163
rect 8079 -2255 8139 -1225
rect 8199 -2195 8259 -1163
rect 8319 -2255 8379 -1225
rect 8439 -1317 8505 -1163
rect 8439 -1381 8440 -1317
rect 8504 -1381 8505 -1317
rect 8439 -1397 8505 -1381
rect 8439 -1461 8440 -1397
rect 8504 -1461 8505 -1397
rect 8439 -1477 8505 -1461
rect 8439 -1541 8440 -1477
rect 8504 -1541 8505 -1477
rect 8439 -1557 8505 -1541
rect 8439 -1621 8440 -1557
rect 8504 -1621 8505 -1557
rect 8439 -1637 8505 -1621
rect 8439 -1701 8440 -1637
rect 8504 -1701 8505 -1637
rect 8439 -1717 8505 -1701
rect 8439 -1781 8440 -1717
rect 8504 -1781 8505 -1717
rect 8439 -1797 8505 -1781
rect 8439 -1861 8440 -1797
rect 8504 -1861 8505 -1797
rect 8439 -1877 8505 -1861
rect 8439 -1941 8440 -1877
rect 8504 -1941 8505 -1877
rect 8439 -1957 8505 -1941
rect 8439 -2021 8440 -1957
rect 8504 -2021 8505 -1957
rect 8439 -2037 8505 -2021
rect 8439 -2101 8440 -2037
rect 8504 -2101 8505 -2037
rect 8439 -2191 8505 -2101
rect 8565 -2255 8625 -1225
rect 8685 -2195 8745 -1163
rect 8805 -2255 8865 -1225
rect 8925 -2195 8985 -1163
rect 9045 -1317 9111 -1163
rect 9045 -1381 9046 -1317
rect 9110 -1381 9111 -1317
rect 9045 -1397 9111 -1381
rect 9045 -1461 9046 -1397
rect 9110 -1461 9111 -1397
rect 9045 -1477 9111 -1461
rect 9045 -1541 9046 -1477
rect 9110 -1541 9111 -1477
rect 9045 -1557 9111 -1541
rect 9045 -1621 9046 -1557
rect 9110 -1621 9111 -1557
rect 9045 -1637 9111 -1621
rect 9045 -1701 9046 -1637
rect 9110 -1701 9111 -1637
rect 9045 -1717 9111 -1701
rect 9045 -1781 9046 -1717
rect 9110 -1781 9111 -1717
rect 9045 -1797 9111 -1781
rect 9045 -1861 9046 -1797
rect 9110 -1861 9111 -1797
rect 9045 -1877 9111 -1861
rect 9045 -1941 9046 -1877
rect 9110 -1941 9111 -1877
rect 9045 -1957 9111 -1941
rect 9045 -2021 9046 -1957
rect 9110 -2021 9111 -1957
rect 9045 -2037 9111 -2021
rect 9045 -2101 9046 -2037
rect 9110 -2101 9111 -2037
rect 9045 -2191 9111 -2101
rect 9171 -2195 9231 -1163
rect 9291 -2255 9351 -1225
rect 9411 -2195 9471 -1163
rect 9531 -2255 9591 -1225
rect 9651 -1317 9717 -1163
rect 9651 -1381 9652 -1317
rect 9716 -1381 9717 -1317
rect 9651 -1397 9717 -1381
rect 9651 -1461 9652 -1397
rect 9716 -1461 9717 -1397
rect 9651 -1477 9717 -1461
rect 9651 -1541 9652 -1477
rect 9716 -1541 9717 -1477
rect 9651 -1557 9717 -1541
rect 9651 -1621 9652 -1557
rect 9716 -1621 9717 -1557
rect 9651 -1637 9717 -1621
rect 9651 -1701 9652 -1637
rect 9716 -1701 9717 -1637
rect 9651 -1717 9717 -1701
rect 9651 -1781 9652 -1717
rect 9716 -1781 9717 -1717
rect 9651 -1797 9717 -1781
rect 9651 -1861 9652 -1797
rect 9716 -1861 9717 -1797
rect 9651 -1877 9717 -1861
rect 9651 -1941 9652 -1877
rect 9716 -1941 9717 -1877
rect 9651 -1957 9717 -1941
rect 9651 -2021 9652 -1957
rect 9716 -2021 9717 -1957
rect 9651 -2037 9717 -2021
rect 9651 -2101 9652 -2037
rect 9716 -2101 9717 -2037
rect 9651 -2191 9717 -2101
rect 9777 -2255 9837 -1225
rect 9897 -2195 9957 -1163
rect 10017 -2255 10077 -1225
rect 10137 -2195 10197 -1163
rect 10257 -1317 10323 -1163
rect 10257 -1381 10258 -1317
rect 10322 -1381 10323 -1317
rect 10257 -1397 10323 -1381
rect 10257 -1461 10258 -1397
rect 10322 -1461 10323 -1397
rect 10257 -1477 10323 -1461
rect 10257 -1541 10258 -1477
rect 10322 -1541 10323 -1477
rect 10257 -1557 10323 -1541
rect 10257 -1621 10258 -1557
rect 10322 -1621 10323 -1557
rect 10257 -1637 10323 -1621
rect 10257 -1701 10258 -1637
rect 10322 -1701 10323 -1637
rect 10257 -1717 10323 -1701
rect 10257 -1781 10258 -1717
rect 10322 -1781 10323 -1717
rect 10257 -1797 10323 -1781
rect 10257 -1861 10258 -1797
rect 10322 -1861 10323 -1797
rect 10257 -1877 10323 -1861
rect 10257 -1941 10258 -1877
rect 10322 -1941 10323 -1877
rect 10257 -1957 10323 -1941
rect 10257 -2021 10258 -1957
rect 10322 -2021 10323 -1957
rect 10257 -2037 10323 -2021
rect 10257 -2101 10258 -2037
rect 10322 -2101 10323 -2037
rect 10257 -2191 10323 -2101
rect 10383 -2195 10443 -1163
rect 10503 -2255 10563 -1225
rect 10623 -2195 10683 -1163
rect 10743 -2255 10803 -1225
rect 10863 -1317 10929 -1163
rect 10863 -1381 10864 -1317
rect 10928 -1381 10929 -1317
rect 10863 -1397 10929 -1381
rect 10863 -1461 10864 -1397
rect 10928 -1461 10929 -1397
rect 10863 -1477 10929 -1461
rect 10863 -1541 10864 -1477
rect 10928 -1541 10929 -1477
rect 10863 -1557 10929 -1541
rect 10863 -1621 10864 -1557
rect 10928 -1621 10929 -1557
rect 10863 -1637 10929 -1621
rect 10863 -1701 10864 -1637
rect 10928 -1701 10929 -1637
rect 10863 -1717 10929 -1701
rect 10863 -1781 10864 -1717
rect 10928 -1781 10929 -1717
rect 10863 -1797 10929 -1781
rect 10863 -1861 10864 -1797
rect 10928 -1861 10929 -1797
rect 10863 -1877 10929 -1861
rect 10863 -1941 10864 -1877
rect 10928 -1941 10929 -1877
rect 10863 -1957 10929 -1941
rect 10863 -2021 10864 -1957
rect 10928 -2021 10929 -1957
rect 10863 -2037 10929 -2021
rect 10863 -2101 10864 -2037
rect 10928 -2101 10929 -2037
rect 10863 -2191 10929 -2101
rect 10989 -2255 11049 -1225
rect 11109 -2195 11169 -1163
rect 11229 -2255 11289 -1225
rect 11349 -2195 11409 -1163
rect 11469 -1317 11535 -1163
rect 11469 -1381 11470 -1317
rect 11534 -1381 11535 -1317
rect 11469 -1397 11535 -1381
rect 11469 -1461 11470 -1397
rect 11534 -1461 11535 -1397
rect 11469 -1477 11535 -1461
rect 11469 -1541 11470 -1477
rect 11534 -1541 11535 -1477
rect 11469 -1557 11535 -1541
rect 11469 -1621 11470 -1557
rect 11534 -1621 11535 -1557
rect 11469 -1637 11535 -1621
rect 11469 -1701 11470 -1637
rect 11534 -1701 11535 -1637
rect 11469 -1717 11535 -1701
rect 11469 -1781 11470 -1717
rect 11534 -1781 11535 -1717
rect 11469 -1797 11535 -1781
rect 11469 -1861 11470 -1797
rect 11534 -1861 11535 -1797
rect 11469 -1877 11535 -1861
rect 11469 -1941 11470 -1877
rect 11534 -1941 11535 -1877
rect 11469 -1957 11535 -1941
rect 11469 -2021 11470 -1957
rect 11534 -2021 11535 -1957
rect 11469 -2037 11535 -2021
rect 11469 -2101 11470 -2037
rect 11534 -2101 11535 -2037
rect 11469 -2191 11535 -2101
rect 11595 -2195 11655 -1163
rect 11715 -2255 11775 -1225
rect 11835 -2195 11895 -1163
rect 11955 -2255 12015 -1225
rect 12075 -1317 12141 -1163
rect 12075 -1381 12076 -1317
rect 12140 -1381 12141 -1317
rect 12075 -1397 12141 -1381
rect 12075 -1461 12076 -1397
rect 12140 -1461 12141 -1397
rect 12075 -1477 12141 -1461
rect 12075 -1541 12076 -1477
rect 12140 -1541 12141 -1477
rect 12075 -1557 12141 -1541
rect 12075 -1621 12076 -1557
rect 12140 -1621 12141 -1557
rect 12075 -1637 12141 -1621
rect 12075 -1701 12076 -1637
rect 12140 -1701 12141 -1637
rect 12075 -1717 12141 -1701
rect 12075 -1781 12076 -1717
rect 12140 -1781 12141 -1717
rect 12075 -1797 12141 -1781
rect 12075 -1861 12076 -1797
rect 12140 -1861 12141 -1797
rect 12075 -1877 12141 -1861
rect 12075 -1941 12076 -1877
rect 12140 -1941 12141 -1877
rect 12075 -1957 12141 -1941
rect 12075 -2021 12076 -1957
rect 12140 -2021 12141 -1957
rect 12075 -2037 12141 -2021
rect 12075 -2101 12076 -2037
rect 12140 -2101 12141 -2037
rect 12075 -2191 12141 -2101
rect 12201 -1097 12873 -1095
rect 12201 -1161 12305 -1097
rect 12369 -1161 12385 -1097
rect 12449 -1161 12465 -1097
rect 12529 -1161 12545 -1097
rect 12609 -1161 12625 -1097
rect 12689 -1161 12705 -1097
rect 12769 -1161 12873 -1097
rect 12201 -1163 12873 -1161
rect 12201 -1317 12267 -1163
rect 12201 -1381 12202 -1317
rect 12266 -1381 12267 -1317
rect 12201 -1397 12267 -1381
rect 12201 -1461 12202 -1397
rect 12266 -1461 12267 -1397
rect 12201 -1477 12267 -1461
rect 12201 -1541 12202 -1477
rect 12266 -1541 12267 -1477
rect 12201 -1557 12267 -1541
rect 12201 -1621 12202 -1557
rect 12266 -1621 12267 -1557
rect 12201 -1637 12267 -1621
rect 12201 -1701 12202 -1637
rect 12266 -1701 12267 -1637
rect 12201 -1717 12267 -1701
rect 12201 -1781 12202 -1717
rect 12266 -1781 12267 -1717
rect 12201 -1797 12267 -1781
rect 12201 -1861 12202 -1797
rect 12266 -1861 12267 -1797
rect 12201 -1877 12267 -1861
rect 12201 -1941 12202 -1877
rect 12266 -1941 12267 -1877
rect 12201 -1957 12267 -1941
rect 12201 -2021 12202 -1957
rect 12266 -2021 12267 -1957
rect 12201 -2037 12267 -2021
rect 12201 -2101 12202 -2037
rect 12266 -2101 12267 -2037
rect 12201 -2191 12267 -2101
rect 12327 -2195 12387 -1163
rect 12447 -2255 12507 -1225
rect 12567 -2195 12627 -1163
rect 12687 -2255 12747 -1225
rect 12807 -1317 12873 -1163
rect 13095 -1098 13525 246
rect 13095 -1113 13526 -1098
rect 13095 -1177 13138 -1113
rect 13202 -1177 13281 -1113
rect 13345 -1177 13401 -1113
rect 13465 -1177 13526 -1113
rect 13095 -1192 13526 -1177
rect 12807 -1381 12808 -1317
rect 12872 -1381 12873 -1317
rect 12807 -1397 12873 -1381
rect 12807 -1461 12808 -1397
rect 12872 -1461 12873 -1397
rect 12807 -1477 12873 -1461
rect 12807 -1541 12808 -1477
rect 12872 -1541 12873 -1477
rect 12807 -1557 12873 -1541
rect 12807 -1621 12808 -1557
rect 12872 -1621 12873 -1557
rect 12807 -1637 12873 -1621
rect 12807 -1701 12808 -1637
rect 12872 -1701 12873 -1637
rect 12807 -1717 12873 -1701
rect 12807 -1781 12808 -1717
rect 12872 -1781 12873 -1717
rect 12807 -1797 12873 -1781
rect 12807 -1861 12808 -1797
rect 12872 -1861 12873 -1797
rect 12807 -1877 12873 -1861
rect 12807 -1941 12808 -1877
rect 12872 -1941 12873 -1877
rect 12807 -1957 12873 -1941
rect 12807 -2021 12808 -1957
rect 12872 -2021 12873 -1957
rect 12807 -2037 12873 -2021
rect 12807 -2101 12808 -2037
rect 12872 -2101 12873 -2037
rect 12807 -2191 12873 -2101
rect 13081 -1658 13543 -1640
rect 13081 -1659 13288 -1658
rect 13081 -1723 13144 -1659
rect 13208 -1722 13288 -1659
rect 13352 -1659 13543 -1658
rect 13352 -1722 13419 -1659
rect 13208 -1723 13419 -1722
rect 13483 -1723 13543 -1659
rect 13081 -2255 13543 -1723
rect 6849 -2257 13543 -2255
rect 6849 -2321 7331 -2257
rect 7395 -2321 7411 -2257
rect 7475 -2321 7491 -2257
rect 7555 -2321 7571 -2257
rect 7635 -2321 7651 -2257
rect 7715 -2321 7731 -2257
rect 7795 -2321 7937 -2257
rect 8001 -2321 8017 -2257
rect 8081 -2321 8097 -2257
rect 8161 -2321 8177 -2257
rect 8241 -2321 8257 -2257
rect 8321 -2321 8337 -2257
rect 8401 -2321 8543 -2257
rect 8607 -2321 8623 -2257
rect 8687 -2321 8703 -2257
rect 8767 -2321 8783 -2257
rect 8847 -2321 8863 -2257
rect 8927 -2321 8943 -2257
rect 9007 -2321 9149 -2257
rect 9213 -2321 9229 -2257
rect 9293 -2321 9309 -2257
rect 9373 -2321 9389 -2257
rect 9453 -2321 9469 -2257
rect 9533 -2321 9549 -2257
rect 9613 -2321 9755 -2257
rect 9819 -2321 9835 -2257
rect 9899 -2321 9915 -2257
rect 9979 -2321 9995 -2257
rect 10059 -2321 10075 -2257
rect 10139 -2321 10155 -2257
rect 10219 -2321 10361 -2257
rect 10425 -2321 10441 -2257
rect 10505 -2321 10521 -2257
rect 10585 -2321 10601 -2257
rect 10665 -2321 10681 -2257
rect 10745 -2321 10761 -2257
rect 10825 -2321 10967 -2257
rect 11031 -2321 11047 -2257
rect 11111 -2321 11127 -2257
rect 11191 -2321 11207 -2257
rect 11271 -2321 11287 -2257
rect 11351 -2321 11367 -2257
rect 11431 -2321 11573 -2257
rect 11637 -2321 11653 -2257
rect 11717 -2321 11733 -2257
rect 11797 -2321 11813 -2257
rect 11877 -2321 11893 -2257
rect 11957 -2321 11973 -2257
rect 12037 -2321 12305 -2257
rect 12369 -2321 12385 -2257
rect 12449 -2321 12465 -2257
rect 12529 -2321 12545 -2257
rect 12609 -2321 12625 -2257
rect 12689 -2321 12705 -2257
rect 12769 -2264 13543 -2257
rect 12769 -2321 12802 -2264
rect 6849 -2328 12802 -2321
rect 12866 -2328 13543 -2264
rect 6849 -2333 13543 -2328
rect 6016 -2338 6142 -2333
rect 12771 -2338 12897 -2333
<< labels >>
flabel metal1 37 1929 705 1976 0 FreeSans 320 0 0 0 x4.IN
flabel metal1 6513 1927 6695 1973 0 FreeSans 320 0 0 0 x4.OUT
flabel metal4 61 2671 523 3281 0 FreeSans 320 0 0 0 x4.VDD
flabel metal4 79 622 509 2061 0 FreeSans 320 0 0 0 x4.VSS
flabel metal1 0 2312 138 2346 0 FreeSans 320 0 0 0 x4.code[3]
flabel metal1 18 1726 412 1773 0 FreeSans 320 0 0 0 x4.code_offset
flabel metal1 5771 600 5829 1756 0 FreeSans 320 0 0 0 x4.code[0]
flabel metal1 4915 601 4973 1778 0 FreeSans 320 0 0 0 x4.code[1]
flabel metal1 2489 601 2547 1778 0 FreeSans 320 0 0 0 x4.code[2]
flabel poly 625 1725 727 1755 0 FreeSans 320 0 0 0 x4.x9.input_stack
flabel space 739 1638 773 1698 0 FreeSans 320 0 0 0 x4.x9.output_stack
flabel space 739 672 773 732 0 FreeSans 320 0 0 0 x4.x9.vss
flabel space 1331 762 1391 1796 0 FreeSans 320 0 0 0 x4.x7.CBOT
flabel space 1451 700 1511 1732 0 FreeSans 320 0 0 0 x4.x7.CTOP
flabel space 1337 1002 1507 1172 0 FreeSans 320 0 0 0 x4.x7.SUB
flabel space 1645 1738 1679 1772 0 FreeSans 320 0 0 0 x4.x7.SW
flabel metal4 1347 1384 1373 1416 0 FreeSans 320 0 0 0 x4.x7.x2.CBOT
flabel metal4 1465 794 1491 826 0 FreeSans 320 0 0 0 x4.x7.x2.CTOP
flabel pwell 1337 1002 1507 1172 0 FreeSans 320 0 0 0 x4.x7.x2.SUB
flabel space 2063 762 2123 1796 0 FreeSans 320 0 0 0 x4.x4[3].CBOT
flabel space 2183 700 2243 1732 0 FreeSans 320 0 0 0 x4.x4[3].CTOP
flabel space 2069 1002 2239 1172 0 FreeSans 320 0 0 0 x4.x4[3].SUB
flabel space 2377 1738 2411 1772 0 FreeSans 320 0 0 0 x4.x4[3].SW
flabel metal4 2079 1384 2105 1416 0 FreeSans 320 0 0 0 x4.x4[3].x2.CBOT
flabel metal4 2197 794 2223 826 0 FreeSans 320 0 0 0 x4.x4[3].x2.CTOP
flabel pwell 2069 1002 2239 1172 0 FreeSans 320 0 0 0 x4.x4[3].x2.SUB
flabel space 2789 762 2849 1796 0 FreeSans 320 0 0 0 x4.x4[2].CBOT
flabel space 2669 700 2729 1732 0 FreeSans 320 0 0 0 x4.x4[2].CTOP
flabel space 2673 1002 2843 1172 0 FreeSans 320 0 0 0 x4.x4[2].SUB
flabel space 2501 1738 2535 1772 0 FreeSans 320 0 0 0 x4.x4[2].SW
flabel metal4 2807 1384 2833 1416 0 FreeSans 320 0 0 0 x4.x4[2].x2.CBOT
flabel metal4 2689 794 2715 826 0 FreeSans 320 0 0 0 x4.x4[2].x2.CTOP
flabel pwell 2673 1002 2843 1172 0 FreeSans 320 0 0 0 x4.x4[2].x2.SUB
flabel space 3275 762 3335 1796 0 FreeSans 320 0 0 0 x4.x4[1].CBOT
flabel space 3395 700 3455 1732 0 FreeSans 320 0 0 0 x4.x4[1].CTOP
flabel space 3281 1002 3451 1172 0 FreeSans 320 0 0 0 x4.x4[1].SUB
flabel space 3589 1738 3623 1772 0 FreeSans 320 0 0 0 x4.x4[1].SW
flabel metal4 3291 1384 3317 1416 0 FreeSans 320 0 0 0 x4.x4[1].x2.CBOT
flabel metal4 3409 794 3435 826 0 FreeSans 320 0 0 0 x4.x4[1].x2.CTOP
flabel pwell 3281 1002 3451 1172 0 FreeSans 320 0 0 0 x4.x4[1].x2.SUB
flabel space 4001 762 4061 1796 0 FreeSans 320 0 0 0 x4.x4[0].CBOT
flabel space 3881 700 3941 1732 0 FreeSans 320 0 0 0 x4.x4[0].CTOP
flabel space 3885 1002 4055 1172 0 FreeSans 320 0 0 0 x4.x4[0].SUB
flabel space 3713 1738 3747 1772 0 FreeSans 320 0 0 0 x4.x4[0].SW
flabel metal4 4019 1384 4045 1416 0 FreeSans 320 0 0 0 x4.x4[0].x2.CBOT
flabel metal4 3901 794 3927 826 0 FreeSans 320 0 0 0 x4.x4[0].x2.CTOP
flabel pwell 3885 1002 4055 1172 0 FreeSans 320 0 0 0 x4.x4[0].x2.SUB
flabel space 4613 762 4673 1796 0 FreeSans 320 0 0 0 x4.x3[1].CBOT
flabel space 4733 700 4793 1732 0 FreeSans 320 0 0 0 x4.x3[1].CTOP
flabel space 4619 1002 4789 1172 0 FreeSans 320 0 0 0 x4.x3[1].SUB
flabel space 4927 1738 4961 1772 0 FreeSans 320 0 0 0 x4.x3[1].SW
flabel metal4 4629 1384 4655 1416 0 FreeSans 320 0 0 0 x4.x3[1].x2.CBOT
flabel metal4 4747 794 4773 826 0 FreeSans 320 0 0 0 x4.x3[1].x2.CTOP
flabel pwell 4619 1002 4789 1172 0 FreeSans 320 0 0 0 x4.x3[1].x2.SUB
flabel space 5339 762 5399 1796 0 FreeSans 320 0 0 0 x4.x3[0].CBOT
flabel space 5219 700 5279 1732 0 FreeSans 320 0 0 0 x4.x3[0].CTOP
flabel space 5223 1002 5393 1172 0 FreeSans 320 0 0 0 x4.x3[0].SUB
flabel space 5051 1738 5085 1772 0 FreeSans 320 0 0 0 x4.x3[0].SW
flabel metal4 5357 1384 5383 1416 0 FreeSans 320 0 0 0 x4.x3[0].x2.CBOT
flabel metal4 5239 794 5265 826 0 FreeSans 320 0 0 0 x4.x3[0].x2.CTOP
flabel pwell 5223 1002 5393 1172 0 FreeSans 320 0 0 0 x4.x3[0].x2.SUB
flabel space 6071 762 6131 1796 0 FreeSans 320 0 0 0 x4.x2.CBOT
flabel space 5951 700 6011 1732 0 FreeSans 320 0 0 0 x4.x2.CTOP
flabel space 5955 1002 6125 1172 0 FreeSans 320 0 0 0 x4.x2.SUB
flabel space 5783 1738 5817 1772 0 FreeSans 320 0 0 0 x4.x2.SW
flabel metal4 6089 1384 6115 1416 0 FreeSans 320 0 0 0 x4.x2.x2.CBOT
flabel metal4 5971 794 5997 826 0 FreeSans 320 0 0 0 x4.x2.x2.CTOP
flabel pwell 5955 1002 6125 1172 0 FreeSans 320 0 0 0 x4.x2.x2.SUB
flabel locali 226 2382 260 2416 0 FreeSans 340 0 0 0 x4.x1.Y
flabel locali 226 2314 260 2348 0 FreeSans 340 0 0 0 x4.x1.Y
flabel locali 134 2314 168 2348 0 FreeSans 340 0 0 0 x4.x1.A
flabel metal1 91 2076 125 2110 0 FreeSans 200 0 0 0 x4.x1.VGND
flabel metal1 91 2620 125 2654 0 FreeSans 200 0 0 0 x4.x1.VPWR
rlabel comment 62 2093 62 2093 4 x4.x1.inv_1
rlabel metal1 62 2045 338 2141 1 x4.x1.VGND
rlabel metal1 62 2589 338 2685 1 x4.x1.VPWR
flabel pwell 91 2076 125 2110 0 FreeSans 200 0 0 0 x4.x1.VNB
flabel nwell 91 2620 125 2654 0 FreeSans 200 0 0 0 x4.x1.VPB
flabel locali 324 2382 358 2416 0 FreeSans 340 0 0 0 x4.x5.Y
flabel locali 324 2314 358 2348 0 FreeSans 340 0 0 0 x4.x5.Y
flabel locali 416 2314 450 2348 0 FreeSans 340 0 0 0 x4.x5.A
flabel metal1 459 2076 493 2110 0 FreeSans 200 0 0 0 x4.x5.VGND
flabel metal1 459 2620 493 2654 0 FreeSans 200 0 0 0 x4.x5.VPWR
rlabel comment 522 2093 522 2093 6 x4.x5.inv_1
rlabel metal1 246 2045 522 2141 1 x4.x5.VGND
rlabel metal1 246 2589 522 2685 1 x4.x5.VPWR
flabel pwell 459 2076 493 2110 0 FreeSans 200 0 0 0 x4.x5.VNB
flabel nwell 459 2620 493 2654 0 FreeSans 200 0 0 0 x4.x5.VPB
flabel metal1 669 2382 703 2416 0 FreeSans 320 0 0 0 x4.x8.input_stack
flabel space 713 3165 747 3225 0 FreeSans 320 0 0 0 x4.x8.vdd
flabel space 713 2475 747 2535 0 FreeSans 320 0 0 0 x4.x8.output_stack
flabel space 983 2733 1153 2903 0 FreeSans 320 0 0 0 x4.x6.SUB
flabel space 977 2109 1037 3143 0 FreeSans 320 0 0 0 x4.x6.CBOT
flabel space 1097 2173 1157 3205 0 FreeSans 320 0 0 0 x4.x6.CTOP
flabel space 1290 2142 1324 2176 0 FreeSans 320 0 0 0 x4.x6.SW
flabel metal4 993 2489 1019 2521 0 FreeSans 320 0 0 0 x4.x6.x1.CBOT
flabel metal4 1111 3079 1137 3111 0 FreeSans 320 0 0 0 x4.x6.x1.CTOP
flabel nwell 983 2733 1153 2903 0 FreeSans 320 0 0 0 x4.x6.x1.SUB
flabel space 1715 2733 1885 2903 0 FreeSans 320 0 0 0 x4.x5[7].SUB
flabel space 1709 2109 1769 3143 0 FreeSans 320 0 0 0 x4.x5[7].CBOT
flabel space 1829 2173 1889 3205 0 FreeSans 320 0 0 0 x4.x5[7].CTOP
flabel space 2022 2142 2056 2176 0 FreeSans 320 0 0 0 x4.x5[7].SW
flabel metal4 1725 2489 1751 2521 0 FreeSans 320 0 0 0 x4.x5[7].x1.CBOT
flabel metal4 1843 3079 1869 3111 0 FreeSans 320 0 0 0 x4.x5[7].x1.CTOP
flabel nwell 1715 2733 1885 2903 0 FreeSans 320 0 0 0 x4.x5[7].x1.SUB
flabel space 2319 2733 2489 2903 0 FreeSans 320 0 0 0 x4.x5[6].SUB
flabel space 2435 2109 2495 3143 0 FreeSans 320 0 0 0 x4.x5[6].CBOT
flabel space 2315 2173 2375 3205 0 FreeSans 320 0 0 0 x4.x5[6].CTOP
flabel space 2148 2142 2182 2176 0 FreeSans 320 0 0 0 x4.x5[6].SW
flabel metal4 2453 2489 2479 2521 0 FreeSans 320 0 0 0 x4.x5[6].x1.CBOT
flabel metal4 2335 3079 2361 3111 0 FreeSans 320 0 0 0 x4.x5[6].x1.CTOP
flabel nwell 2319 2733 2489 2903 0 FreeSans 320 0 0 0 x4.x5[6].x1.SUB
flabel space 2927 2733 3097 2903 0 FreeSans 320 0 0 0 x4.x5[5].SUB
flabel space 2921 2109 2981 3143 0 FreeSans 320 0 0 0 x4.x5[5].CBOT
flabel space 3041 2173 3101 3205 0 FreeSans 320 0 0 0 x4.x5[5].CTOP
flabel space 3234 2142 3268 2176 0 FreeSans 320 0 0 0 x4.x5[5].SW
flabel metal4 2937 2489 2963 2521 0 FreeSans 320 0 0 0 x4.x5[5].x1.CBOT
flabel metal4 3055 3079 3081 3111 0 FreeSans 320 0 0 0 x4.x5[5].x1.CTOP
flabel nwell 2927 2733 3097 2903 0 FreeSans 320 0 0 0 x4.x5[5].x1.SUB
flabel space 3531 2733 3701 2903 0 FreeSans 320 0 0 0 x4.x5[4].SUB
flabel space 3647 2109 3707 3143 0 FreeSans 320 0 0 0 x4.x5[4].CBOT
flabel space 3527 2173 3587 3205 0 FreeSans 320 0 0 0 x4.x5[4].CTOP
flabel space 3360 2142 3394 2176 0 FreeSans 320 0 0 0 x4.x5[4].SW
flabel metal4 3665 2489 3691 2521 0 FreeSans 320 0 0 0 x4.x5[4].x1.CBOT
flabel metal4 3547 3079 3573 3111 0 FreeSans 320 0 0 0 x4.x5[4].x1.CTOP
flabel nwell 3531 2733 3701 2903 0 FreeSans 320 0 0 0 x4.x5[4].x1.SUB
flabel space 4139 2733 4309 2903 0 FreeSans 320 0 0 0 x4.x5[3].SUB
flabel space 4133 2109 4193 3143 0 FreeSans 320 0 0 0 x4.x5[3].CBOT
flabel space 4253 2173 4313 3205 0 FreeSans 320 0 0 0 x4.x5[3].CTOP
flabel space 4446 2142 4480 2176 0 FreeSans 320 0 0 0 x4.x5[3].SW
flabel metal4 4149 2489 4175 2521 0 FreeSans 320 0 0 0 x4.x5[3].x1.CBOT
flabel metal4 4267 3079 4293 3111 0 FreeSans 320 0 0 0 x4.x5[3].x1.CTOP
flabel nwell 4139 2733 4309 2903 0 FreeSans 320 0 0 0 x4.x5[3].x1.SUB
flabel space 4743 2733 4913 2903 0 FreeSans 320 0 0 0 x4.x5[2].SUB
flabel space 4859 2109 4919 3143 0 FreeSans 320 0 0 0 x4.x5[2].CBOT
flabel space 4739 2173 4799 3205 0 FreeSans 320 0 0 0 x4.x5[2].CTOP
flabel space 4572 2142 4606 2176 0 FreeSans 320 0 0 0 x4.x5[2].SW
flabel metal4 4877 2489 4903 2521 0 FreeSans 320 0 0 0 x4.x5[2].x1.CBOT
flabel metal4 4759 3079 4785 3111 0 FreeSans 320 0 0 0 x4.x5[2].x1.CTOP
flabel nwell 4743 2733 4913 2903 0 FreeSans 320 0 0 0 x4.x5[2].x1.SUB
flabel space 5351 2733 5521 2903 0 FreeSans 320 0 0 0 x4.x5[1].SUB
flabel space 5345 2109 5405 3143 0 FreeSans 320 0 0 0 x4.x5[1].CBOT
flabel space 5465 2173 5525 3205 0 FreeSans 320 0 0 0 x4.x5[1].CTOP
flabel space 5658 2142 5692 2176 0 FreeSans 320 0 0 0 x4.x5[1].SW
flabel metal4 5361 2489 5387 2521 0 FreeSans 320 0 0 0 x4.x5[1].x1.CBOT
flabel metal4 5479 3079 5505 3111 0 FreeSans 320 0 0 0 x4.x5[1].x1.CTOP
flabel nwell 5351 2733 5521 2903 0 FreeSans 320 0 0 0 x4.x5[1].x1.SUB
flabel space 5955 2733 6125 2903 0 FreeSans 320 0 0 0 x4.x5[0].SUB
flabel space 6071 2109 6131 3143 0 FreeSans 320 0 0 0 x4.x5[0].CBOT
flabel space 5951 2173 6011 3205 0 FreeSans 320 0 0 0 x4.x5[0].CTOP
flabel space 5784 2142 5818 2176 0 FreeSans 320 0 0 0 x4.x5[0].SW
flabel metal4 6089 2489 6115 2521 0 FreeSans 320 0 0 0 x4.x5[0].x1.CBOT
flabel metal4 5971 3079 5997 3111 0 FreeSans 320 0 0 0 x4.x5[0].x1.CTOP
flabel nwell 5955 2733 6125 2903 0 FreeSans 320 0 0 0 x4.x5[0].x1.SUB
flabel metal1 6144 -1028 6812 -981 0 FreeSans 320 0 0 0 x3.IN
flabel metal1 154 -1025 336 -979 0 FreeSans 320 0 0 0 x3.OUT
flabel metal4 6326 -2333 6788 -1723 0 FreeSans 320 0 0 0 x3.VDD
flabel metal4 6340 -1113 6770 326 0 FreeSans 320 0 0 0 x3.VSS
flabel metal1 6711 -1398 6849 -1364 0 FreeSans 320 0 0 0 x3.code[3]
flabel metal1 6437 -825 6831 -778 0 FreeSans 320 0 0 0 x3.code_offset
flabel metal1 1020 -808 1078 348 0 FreeSans 320 0 0 0 x3.code[0]
flabel metal1 1876 -830 1934 347 0 FreeSans 320 0 0 0 x3.code[1]
flabel metal1 4302 -830 4360 347 0 FreeSans 320 0 0 0 x3.code[2]
flabel poly 6122 -807 6224 -777 0 FreeSans 320 0 0 0 x3.x9.input_stack
flabel space 6076 -750 6110 -690 0 FreeSans 320 0 0 0 x3.x9.output_stack
flabel space 6076 216 6110 276 0 FreeSans 320 0 0 0 x3.x9.vss
flabel space 5458 -848 5518 186 0 FreeSans 320 0 0 0 x3.x7.CBOT
flabel space 5338 -784 5398 248 0 FreeSans 320 0 0 0 x3.x7.CTOP
flabel space 5342 -224 5512 -54 0 FreeSans 320 0 0 0 x3.x7.SUB
flabel space 5170 -824 5204 -790 0 FreeSans 320 0 0 0 x3.x7.SW
flabel metal4 5476 -468 5502 -436 0 FreeSans 320 0 0 0 x3.x7.x2.CBOT
flabel metal4 5358 122 5384 154 0 FreeSans 320 0 0 0 x3.x7.x2.CTOP
flabel pwell 5342 -224 5512 -54 0 FreeSans 320 0 0 0 x3.x7.x2.SUB
flabel space 4726 -848 4786 186 0 FreeSans 320 0 0 0 x3.x4[3].CBOT
flabel space 4606 -784 4666 248 0 FreeSans 320 0 0 0 x3.x4[3].CTOP
flabel space 4610 -224 4780 -54 0 FreeSans 320 0 0 0 x3.x4[3].SUB
flabel space 4438 -824 4472 -790 0 FreeSans 320 0 0 0 x3.x4[3].SW
flabel metal4 4744 -468 4770 -436 0 FreeSans 320 0 0 0 x3.x4[3].x2.CBOT
flabel metal4 4626 122 4652 154 0 FreeSans 320 0 0 0 x3.x4[3].x2.CTOP
flabel pwell 4610 -224 4780 -54 0 FreeSans 320 0 0 0 x3.x4[3].x2.SUB
flabel space 4000 -848 4060 186 0 FreeSans 320 0 0 0 x3.x4[2].CBOT
flabel space 4120 -784 4180 248 0 FreeSans 320 0 0 0 x3.x4[2].CTOP
flabel space 4006 -224 4176 -54 0 FreeSans 320 0 0 0 x3.x4[2].SUB
flabel space 4314 -824 4348 -790 0 FreeSans 320 0 0 0 x3.x4[2].SW
flabel metal4 4016 -468 4042 -436 0 FreeSans 320 0 0 0 x3.x4[2].x2.CBOT
flabel metal4 4134 122 4160 154 0 FreeSans 320 0 0 0 x3.x4[2].x2.CTOP
flabel pwell 4006 -224 4176 -54 0 FreeSans 320 0 0 0 x3.x4[2].x2.SUB
flabel space 3514 -848 3574 186 0 FreeSans 320 0 0 0 x3.x4[1].CBOT
flabel space 3394 -784 3454 248 0 FreeSans 320 0 0 0 x3.x4[1].CTOP
flabel space 3398 -224 3568 -54 0 FreeSans 320 0 0 0 x3.x4[1].SUB
flabel space 3226 -824 3260 -790 0 FreeSans 320 0 0 0 x3.x4[1].SW
flabel metal4 3532 -468 3558 -436 0 FreeSans 320 0 0 0 x3.x4[1].x2.CBOT
flabel metal4 3414 122 3440 154 0 FreeSans 320 0 0 0 x3.x4[1].x2.CTOP
flabel pwell 3398 -224 3568 -54 0 FreeSans 320 0 0 0 x3.x4[1].x2.SUB
flabel space 2788 -848 2848 186 0 FreeSans 320 0 0 0 x3.x4[0].CBOT
flabel space 2908 -784 2968 248 0 FreeSans 320 0 0 0 x3.x4[0].CTOP
flabel space 2794 -224 2964 -54 0 FreeSans 320 0 0 0 x3.x4[0].SUB
flabel space 3102 -824 3136 -790 0 FreeSans 320 0 0 0 x3.x4[0].SW
flabel metal4 2804 -468 2830 -436 0 FreeSans 320 0 0 0 x3.x4[0].x2.CBOT
flabel metal4 2922 122 2948 154 0 FreeSans 320 0 0 0 x3.x4[0].x2.CTOP
flabel pwell 2794 -224 2964 -54 0 FreeSans 320 0 0 0 x3.x4[0].x2.SUB
flabel space 2176 -848 2236 186 0 FreeSans 320 0 0 0 x3.x3[1].CBOT
flabel space 2056 -784 2116 248 0 FreeSans 320 0 0 0 x3.x3[1].CTOP
flabel space 2060 -224 2230 -54 0 FreeSans 320 0 0 0 x3.x3[1].SUB
flabel space 1888 -824 1922 -790 0 FreeSans 320 0 0 0 x3.x3[1].SW
flabel metal4 2194 -468 2220 -436 0 FreeSans 320 0 0 0 x3.x3[1].x2.CBOT
flabel metal4 2076 122 2102 154 0 FreeSans 320 0 0 0 x3.x3[1].x2.CTOP
flabel pwell 2060 -224 2230 -54 0 FreeSans 320 0 0 0 x3.x3[1].x2.SUB
flabel space 1450 -848 1510 186 0 FreeSans 320 0 0 0 x3.x3[0].CBOT
flabel space 1570 -784 1630 248 0 FreeSans 320 0 0 0 x3.x3[0].CTOP
flabel space 1456 -224 1626 -54 0 FreeSans 320 0 0 0 x3.x3[0].SUB
flabel space 1764 -824 1798 -790 0 FreeSans 320 0 0 0 x3.x3[0].SW
flabel metal4 1466 -468 1492 -436 0 FreeSans 320 0 0 0 x3.x3[0].x2.CBOT
flabel metal4 1584 122 1610 154 0 FreeSans 320 0 0 0 x3.x3[0].x2.CTOP
flabel pwell 1456 -224 1626 -54 0 FreeSans 320 0 0 0 x3.x3[0].x2.SUB
flabel space 718 -848 778 186 0 FreeSans 320 0 0 0 x3.x2.CBOT
flabel space 838 -784 898 248 0 FreeSans 320 0 0 0 x3.x2.CTOP
flabel space 724 -224 894 -54 0 FreeSans 320 0 0 0 x3.x2.SUB
flabel space 1032 -824 1066 -790 0 FreeSans 320 0 0 0 x3.x2.SW
flabel metal4 734 -468 760 -436 0 FreeSans 320 0 0 0 x3.x2.x2.CBOT
flabel metal4 852 122 878 154 0 FreeSans 320 0 0 0 x3.x2.x2.CTOP
flabel pwell 724 -224 894 -54 0 FreeSans 320 0 0 0 x3.x2.x2.SUB
flabel locali 6589 -1468 6623 -1434 0 FreeSans 340 0 0 0 x3.x1.Y
flabel locali 6589 -1400 6623 -1366 0 FreeSans 340 0 0 0 x3.x1.Y
flabel locali 6681 -1400 6715 -1366 0 FreeSans 340 0 0 0 x3.x1.A
flabel metal1 6724 -1162 6758 -1128 0 FreeSans 200 0 0 0 x3.x1.VGND
flabel metal1 6724 -1706 6758 -1672 0 FreeSans 200 0 0 0 x3.x1.VPWR
rlabel comment 6787 -1145 6787 -1145 8 x3.x1.inv_1
rlabel metal1 6511 -1193 6787 -1097 5 x3.x1.VGND
rlabel metal1 6511 -1737 6787 -1641 5 x3.x1.VPWR
flabel pwell 6724 -1162 6758 -1128 0 FreeSans 200 0 0 0 x3.x1.VNB
flabel nwell 6724 -1706 6758 -1672 0 FreeSans 200 0 0 0 x3.x1.VPB
flabel locali 6491 -1468 6525 -1434 0 FreeSans 340 0 0 0 x3.x5.Y
flabel locali 6491 -1400 6525 -1366 0 FreeSans 340 0 0 0 x3.x5.Y
flabel locali 6399 -1400 6433 -1366 0 FreeSans 340 0 0 0 x3.x5.A
flabel metal1 6356 -1162 6390 -1128 0 FreeSans 200 0 0 0 x3.x5.VGND
flabel metal1 6356 -1706 6390 -1672 0 FreeSans 200 0 0 0 x3.x5.VPWR
rlabel comment 6327 -1145 6327 -1145 2 x3.x5.inv_1
rlabel metal1 6327 -1193 6603 -1097 5 x3.x5.VGND
rlabel metal1 6327 -1737 6603 -1641 5 x3.x5.VPWR
flabel pwell 6356 -1162 6390 -1128 0 FreeSans 200 0 0 0 x3.x5.VNB
flabel nwell 6356 -1706 6390 -1672 0 FreeSans 200 0 0 0 x3.x5.VPB
flabel metal1 6146 -1468 6180 -1434 0 FreeSans 320 0 0 0 x3.x8.input_stack
flabel space 6102 -2277 6136 -2217 0 FreeSans 320 0 0 0 x3.x8.vdd
flabel space 6102 -1587 6136 -1527 0 FreeSans 320 0 0 0 x3.x8.output_stack
flabel space 5696 -1955 5866 -1785 0 FreeSans 320 0 0 0 x3.x6.SUB
flabel space 5812 -2195 5872 -1161 0 FreeSans 320 0 0 0 x3.x6.CBOT
flabel space 5692 -2257 5752 -1225 0 FreeSans 320 0 0 0 x3.x6.CTOP
flabel space 5525 -1228 5559 -1194 0 FreeSans 320 0 0 0 x3.x6.SW
flabel metal4 5830 -1573 5856 -1541 0 FreeSans 320 0 0 0 x3.x6.x1.CBOT
flabel metal4 5712 -2163 5738 -2131 0 FreeSans 320 0 0 0 x3.x6.x1.CTOP
flabel nwell 5696 -1955 5866 -1785 0 FreeSans 320 0 0 0 x3.x6.x1.SUB
flabel space 4964 -1955 5134 -1785 0 FreeSans 320 0 0 0 x3.x5[7].SUB
flabel space 5080 -2195 5140 -1161 0 FreeSans 320 0 0 0 x3.x5[7].CBOT
flabel space 4960 -2257 5020 -1225 0 FreeSans 320 0 0 0 x3.x5[7].CTOP
flabel space 4793 -1228 4827 -1194 0 FreeSans 320 0 0 0 x3.x5[7].SW
flabel metal4 5098 -1573 5124 -1541 0 FreeSans 320 0 0 0 x3.x5[7].x1.CBOT
flabel metal4 4980 -2163 5006 -2131 0 FreeSans 320 0 0 0 x3.x5[7].x1.CTOP
flabel nwell 4964 -1955 5134 -1785 0 FreeSans 320 0 0 0 x3.x5[7].x1.SUB
flabel space 4360 -1955 4530 -1785 0 FreeSans 320 0 0 0 x3.x5[6].SUB
flabel space 4354 -2195 4414 -1161 0 FreeSans 320 0 0 0 x3.x5[6].CBOT
flabel space 4474 -2257 4534 -1225 0 FreeSans 320 0 0 0 x3.x5[6].CTOP
flabel space 4667 -1228 4701 -1194 0 FreeSans 320 0 0 0 x3.x5[6].SW
flabel metal4 4370 -1573 4396 -1541 0 FreeSans 320 0 0 0 x3.x5[6].x1.CBOT
flabel metal4 4488 -2163 4514 -2131 0 FreeSans 320 0 0 0 x3.x5[6].x1.CTOP
flabel nwell 4360 -1955 4530 -1785 0 FreeSans 320 0 0 0 x3.x5[6].x1.SUB
flabel space 3752 -1955 3922 -1785 0 FreeSans 320 0 0 0 x3.x5[5].SUB
flabel space 3868 -2195 3928 -1161 0 FreeSans 320 0 0 0 x3.x5[5].CBOT
flabel space 3748 -2257 3808 -1225 0 FreeSans 320 0 0 0 x3.x5[5].CTOP
flabel space 3581 -1228 3615 -1194 0 FreeSans 320 0 0 0 x3.x5[5].SW
flabel metal4 3886 -1573 3912 -1541 0 FreeSans 320 0 0 0 x3.x5[5].x1.CBOT
flabel metal4 3768 -2163 3794 -2131 0 FreeSans 320 0 0 0 x3.x5[5].x1.CTOP
flabel nwell 3752 -1955 3922 -1785 0 FreeSans 320 0 0 0 x3.x5[5].x1.SUB
flabel space 3148 -1955 3318 -1785 0 FreeSans 320 0 0 0 x3.x5[4].SUB
flabel space 3142 -2195 3202 -1161 0 FreeSans 320 0 0 0 x3.x5[4].CBOT
flabel space 3262 -2257 3322 -1225 0 FreeSans 320 0 0 0 x3.x5[4].CTOP
flabel space 3455 -1228 3489 -1194 0 FreeSans 320 0 0 0 x3.x5[4].SW
flabel metal4 3158 -1573 3184 -1541 0 FreeSans 320 0 0 0 x3.x5[4].x1.CBOT
flabel metal4 3276 -2163 3302 -2131 0 FreeSans 320 0 0 0 x3.x5[4].x1.CTOP
flabel nwell 3148 -1955 3318 -1785 0 FreeSans 320 0 0 0 x3.x5[4].x1.SUB
flabel space 2540 -1955 2710 -1785 0 FreeSans 320 0 0 0 x3.x5[3].SUB
flabel space 2656 -2195 2716 -1161 0 FreeSans 320 0 0 0 x3.x5[3].CBOT
flabel space 2536 -2257 2596 -1225 0 FreeSans 320 0 0 0 x3.x5[3].CTOP
flabel space 2369 -1228 2403 -1194 0 FreeSans 320 0 0 0 x3.x5[3].SW
flabel metal4 2674 -1573 2700 -1541 0 FreeSans 320 0 0 0 x3.x5[3].x1.CBOT
flabel metal4 2556 -2163 2582 -2131 0 FreeSans 320 0 0 0 x3.x5[3].x1.CTOP
flabel nwell 2540 -1955 2710 -1785 0 FreeSans 320 0 0 0 x3.x5[3].x1.SUB
flabel space 1936 -1955 2106 -1785 0 FreeSans 320 0 0 0 x3.x5[2].SUB
flabel space 1930 -2195 1990 -1161 0 FreeSans 320 0 0 0 x3.x5[2].CBOT
flabel space 2050 -2257 2110 -1225 0 FreeSans 320 0 0 0 x3.x5[2].CTOP
flabel space 2243 -1228 2277 -1194 0 FreeSans 320 0 0 0 x3.x5[2].SW
flabel metal4 1946 -1573 1972 -1541 0 FreeSans 320 0 0 0 x3.x5[2].x1.CBOT
flabel metal4 2064 -2163 2090 -2131 0 FreeSans 320 0 0 0 x3.x5[2].x1.CTOP
flabel nwell 1936 -1955 2106 -1785 0 FreeSans 320 0 0 0 x3.x5[2].x1.SUB
flabel space 1328 -1955 1498 -1785 0 FreeSans 320 0 0 0 x3.x5[1].SUB
flabel space 1444 -2195 1504 -1161 0 FreeSans 320 0 0 0 x3.x5[1].CBOT
flabel space 1324 -2257 1384 -1225 0 FreeSans 320 0 0 0 x3.x5[1].CTOP
flabel space 1157 -1228 1191 -1194 0 FreeSans 320 0 0 0 x3.x5[1].SW
flabel metal4 1462 -1573 1488 -1541 0 FreeSans 320 0 0 0 x3.x5[1].x1.CBOT
flabel metal4 1344 -2163 1370 -2131 0 FreeSans 320 0 0 0 x3.x5[1].x1.CTOP
flabel nwell 1328 -1955 1498 -1785 0 FreeSans 320 0 0 0 x3.x5[1].x1.SUB
flabel space 724 -1955 894 -1785 0 FreeSans 320 0 0 0 x3.x5[0].SUB
flabel space 718 -2195 778 -1161 0 FreeSans 320 0 0 0 x3.x5[0].CBOT
flabel space 838 -2257 898 -1225 0 FreeSans 320 0 0 0 x3.x5[0].CTOP
flabel space 1031 -1228 1065 -1194 0 FreeSans 320 0 0 0 x3.x5[0].SW
flabel metal4 734 -1573 760 -1541 0 FreeSans 320 0 0 0 x3.x5[0].x1.CBOT
flabel metal4 852 -2163 878 -2131 0 FreeSans 320 0 0 0 x3.x5[0].x1.CTOP
flabel nwell 724 -1955 894 -1785 0 FreeSans 320 0 0 0 x3.x5[0].x1.SUB
flabel metal1 12899 -1028 13567 -981 0 FreeSans 320 0 0 0 x2.IN
flabel metal1 6909 -1025 7091 -979 0 FreeSans 320 0 0 0 x2.OUT
flabel metal4 13081 -2333 13543 -1723 0 FreeSans 320 0 0 0 x2.VDD
flabel metal4 13095 -1113 13525 326 0 FreeSans 320 0 0 0 x2.VSS
flabel metal1 13466 -1398 13604 -1364 0 FreeSans 320 0 0 0 x2.code[3]
flabel metal1 13192 -825 13586 -778 0 FreeSans 320 0 0 0 x2.code_offset
flabel metal1 7775 -808 7833 348 0 FreeSans 320 0 0 0 x2.code[0]
flabel metal1 8631 -830 8689 347 0 FreeSans 320 0 0 0 x2.code[1]
flabel metal1 11057 -830 11115 347 0 FreeSans 320 0 0 0 x2.code[2]
flabel poly 12877 -807 12979 -777 0 FreeSans 320 0 0 0 x2.x9.input_stack
flabel space 12831 -750 12865 -690 0 FreeSans 320 0 0 0 x2.x9.output_stack
flabel space 12831 216 12865 276 0 FreeSans 320 0 0 0 x2.x9.vss
flabel space 12213 -848 12273 186 0 FreeSans 320 0 0 0 x2.x7.CBOT
flabel space 12093 -784 12153 248 0 FreeSans 320 0 0 0 x2.x7.CTOP
flabel space 12097 -224 12267 -54 0 FreeSans 320 0 0 0 x2.x7.SUB
flabel space 11925 -824 11959 -790 0 FreeSans 320 0 0 0 x2.x7.SW
flabel metal4 12231 -468 12257 -436 0 FreeSans 320 0 0 0 x2.x7.x2.CBOT
flabel metal4 12113 122 12139 154 0 FreeSans 320 0 0 0 x2.x7.x2.CTOP
flabel pwell 12097 -224 12267 -54 0 FreeSans 320 0 0 0 x2.x7.x2.SUB
flabel space 11481 -848 11541 186 0 FreeSans 320 0 0 0 x2.x4[3].CBOT
flabel space 11361 -784 11421 248 0 FreeSans 320 0 0 0 x2.x4[3].CTOP
flabel space 11365 -224 11535 -54 0 FreeSans 320 0 0 0 x2.x4[3].SUB
flabel space 11193 -824 11227 -790 0 FreeSans 320 0 0 0 x2.x4[3].SW
flabel metal4 11499 -468 11525 -436 0 FreeSans 320 0 0 0 x2.x4[3].x2.CBOT
flabel metal4 11381 122 11407 154 0 FreeSans 320 0 0 0 x2.x4[3].x2.CTOP
flabel pwell 11365 -224 11535 -54 0 FreeSans 320 0 0 0 x2.x4[3].x2.SUB
flabel space 10755 -848 10815 186 0 FreeSans 320 0 0 0 x2.x4[2].CBOT
flabel space 10875 -784 10935 248 0 FreeSans 320 0 0 0 x2.x4[2].CTOP
flabel space 10761 -224 10931 -54 0 FreeSans 320 0 0 0 x2.x4[2].SUB
flabel space 11069 -824 11103 -790 0 FreeSans 320 0 0 0 x2.x4[2].SW
flabel metal4 10771 -468 10797 -436 0 FreeSans 320 0 0 0 x2.x4[2].x2.CBOT
flabel metal4 10889 122 10915 154 0 FreeSans 320 0 0 0 x2.x4[2].x2.CTOP
flabel pwell 10761 -224 10931 -54 0 FreeSans 320 0 0 0 x2.x4[2].x2.SUB
flabel space 10269 -848 10329 186 0 FreeSans 320 0 0 0 x2.x4[1].CBOT
flabel space 10149 -784 10209 248 0 FreeSans 320 0 0 0 x2.x4[1].CTOP
flabel space 10153 -224 10323 -54 0 FreeSans 320 0 0 0 x2.x4[1].SUB
flabel space 9981 -824 10015 -790 0 FreeSans 320 0 0 0 x2.x4[1].SW
flabel metal4 10287 -468 10313 -436 0 FreeSans 320 0 0 0 x2.x4[1].x2.CBOT
flabel metal4 10169 122 10195 154 0 FreeSans 320 0 0 0 x2.x4[1].x2.CTOP
flabel pwell 10153 -224 10323 -54 0 FreeSans 320 0 0 0 x2.x4[1].x2.SUB
flabel space 9543 -848 9603 186 0 FreeSans 320 0 0 0 x2.x4[0].CBOT
flabel space 9663 -784 9723 248 0 FreeSans 320 0 0 0 x2.x4[0].CTOP
flabel space 9549 -224 9719 -54 0 FreeSans 320 0 0 0 x2.x4[0].SUB
flabel space 9857 -824 9891 -790 0 FreeSans 320 0 0 0 x2.x4[0].SW
flabel metal4 9559 -468 9585 -436 0 FreeSans 320 0 0 0 x2.x4[0].x2.CBOT
flabel metal4 9677 122 9703 154 0 FreeSans 320 0 0 0 x2.x4[0].x2.CTOP
flabel pwell 9549 -224 9719 -54 0 FreeSans 320 0 0 0 x2.x4[0].x2.SUB
flabel space 8931 -848 8991 186 0 FreeSans 320 0 0 0 x2.x3[1].CBOT
flabel space 8811 -784 8871 248 0 FreeSans 320 0 0 0 x2.x3[1].CTOP
flabel space 8815 -224 8985 -54 0 FreeSans 320 0 0 0 x2.x3[1].SUB
flabel space 8643 -824 8677 -790 0 FreeSans 320 0 0 0 x2.x3[1].SW
flabel metal4 8949 -468 8975 -436 0 FreeSans 320 0 0 0 x2.x3[1].x2.CBOT
flabel metal4 8831 122 8857 154 0 FreeSans 320 0 0 0 x2.x3[1].x2.CTOP
flabel pwell 8815 -224 8985 -54 0 FreeSans 320 0 0 0 x2.x3[1].x2.SUB
flabel space 8205 -848 8265 186 0 FreeSans 320 0 0 0 x2.x3[0].CBOT
flabel space 8325 -784 8385 248 0 FreeSans 320 0 0 0 x2.x3[0].CTOP
flabel space 8211 -224 8381 -54 0 FreeSans 320 0 0 0 x2.x3[0].SUB
flabel space 8519 -824 8553 -790 0 FreeSans 320 0 0 0 x2.x3[0].SW
flabel metal4 8221 -468 8247 -436 0 FreeSans 320 0 0 0 x2.x3[0].x2.CBOT
flabel metal4 8339 122 8365 154 0 FreeSans 320 0 0 0 x2.x3[0].x2.CTOP
flabel pwell 8211 -224 8381 -54 0 FreeSans 320 0 0 0 x2.x3[0].x2.SUB
flabel space 7473 -848 7533 186 0 FreeSans 320 0 0 0 x2.x2.CBOT
flabel space 7593 -784 7653 248 0 FreeSans 320 0 0 0 x2.x2.CTOP
flabel space 7479 -224 7649 -54 0 FreeSans 320 0 0 0 x2.x2.SUB
flabel space 7787 -824 7821 -790 0 FreeSans 320 0 0 0 x2.x2.SW
flabel metal4 7489 -468 7515 -436 0 FreeSans 320 0 0 0 x2.x2.x2.CBOT
flabel metal4 7607 122 7633 154 0 FreeSans 320 0 0 0 x2.x2.x2.CTOP
flabel pwell 7479 -224 7649 -54 0 FreeSans 320 0 0 0 x2.x2.x2.SUB
flabel locali 13344 -1468 13378 -1434 0 FreeSans 340 0 0 0 x2.x1.Y
flabel locali 13344 -1400 13378 -1366 0 FreeSans 340 0 0 0 x2.x1.Y
flabel locali 13436 -1400 13470 -1366 0 FreeSans 340 0 0 0 x2.x1.A
flabel metal1 13479 -1162 13513 -1128 0 FreeSans 200 0 0 0 x2.x1.VGND
flabel metal1 13479 -1706 13513 -1672 0 FreeSans 200 0 0 0 x2.x1.VPWR
rlabel comment 13542 -1145 13542 -1145 8 x2.x1.inv_1
rlabel metal1 13266 -1193 13542 -1097 5 x2.x1.VGND
rlabel metal1 13266 -1737 13542 -1641 5 x2.x1.VPWR
flabel pwell 13479 -1162 13513 -1128 0 FreeSans 200 0 0 0 x2.x1.VNB
flabel nwell 13479 -1706 13513 -1672 0 FreeSans 200 0 0 0 x2.x1.VPB
flabel locali 13246 -1468 13280 -1434 0 FreeSans 340 0 0 0 x2.x5.Y
flabel locali 13246 -1400 13280 -1366 0 FreeSans 340 0 0 0 x2.x5.Y
flabel locali 13154 -1400 13188 -1366 0 FreeSans 340 0 0 0 x2.x5.A
flabel metal1 13111 -1162 13145 -1128 0 FreeSans 200 0 0 0 x2.x5.VGND
flabel metal1 13111 -1706 13145 -1672 0 FreeSans 200 0 0 0 x2.x5.VPWR
rlabel comment 13082 -1145 13082 -1145 2 x2.x5.inv_1
rlabel metal1 13082 -1193 13358 -1097 5 x2.x5.VGND
rlabel metal1 13082 -1737 13358 -1641 5 x2.x5.VPWR
flabel pwell 13111 -1162 13145 -1128 0 FreeSans 200 0 0 0 x2.x5.VNB
flabel nwell 13111 -1706 13145 -1672 0 FreeSans 200 0 0 0 x2.x5.VPB
flabel metal1 12901 -1468 12935 -1434 0 FreeSans 320 0 0 0 x2.x8.input_stack
flabel space 12857 -2277 12891 -2217 0 FreeSans 320 0 0 0 x2.x8.vdd
flabel space 12857 -1587 12891 -1527 0 FreeSans 320 0 0 0 x2.x8.output_stack
flabel space 12451 -1955 12621 -1785 0 FreeSans 320 0 0 0 x2.x6.SUB
flabel space 12567 -2195 12627 -1161 0 FreeSans 320 0 0 0 x2.x6.CBOT
flabel space 12447 -2257 12507 -1225 0 FreeSans 320 0 0 0 x2.x6.CTOP
flabel space 12280 -1228 12314 -1194 0 FreeSans 320 0 0 0 x2.x6.SW
flabel metal4 12585 -1573 12611 -1541 0 FreeSans 320 0 0 0 x2.x6.x1.CBOT
flabel metal4 12467 -2163 12493 -2131 0 FreeSans 320 0 0 0 x2.x6.x1.CTOP
flabel nwell 12451 -1955 12621 -1785 0 FreeSans 320 0 0 0 x2.x6.x1.SUB
flabel space 11719 -1955 11889 -1785 0 FreeSans 320 0 0 0 x2.x5[7].SUB
flabel space 11835 -2195 11895 -1161 0 FreeSans 320 0 0 0 x2.x5[7].CBOT
flabel space 11715 -2257 11775 -1225 0 FreeSans 320 0 0 0 x2.x5[7].CTOP
flabel space 11548 -1228 11582 -1194 0 FreeSans 320 0 0 0 x2.x5[7].SW
flabel metal4 11853 -1573 11879 -1541 0 FreeSans 320 0 0 0 x2.x5[7].x1.CBOT
flabel metal4 11735 -2163 11761 -2131 0 FreeSans 320 0 0 0 x2.x5[7].x1.CTOP
flabel nwell 11719 -1955 11889 -1785 0 FreeSans 320 0 0 0 x2.x5[7].x1.SUB
flabel space 11115 -1955 11285 -1785 0 FreeSans 320 0 0 0 x2.x5[6].SUB
flabel space 11109 -2195 11169 -1161 0 FreeSans 320 0 0 0 x2.x5[6].CBOT
flabel space 11229 -2257 11289 -1225 0 FreeSans 320 0 0 0 x2.x5[6].CTOP
flabel space 11422 -1228 11456 -1194 0 FreeSans 320 0 0 0 x2.x5[6].SW
flabel metal4 11125 -1573 11151 -1541 0 FreeSans 320 0 0 0 x2.x5[6].x1.CBOT
flabel metal4 11243 -2163 11269 -2131 0 FreeSans 320 0 0 0 x2.x5[6].x1.CTOP
flabel nwell 11115 -1955 11285 -1785 0 FreeSans 320 0 0 0 x2.x5[6].x1.SUB
flabel space 10507 -1955 10677 -1785 0 FreeSans 320 0 0 0 x2.x5[5].SUB
flabel space 10623 -2195 10683 -1161 0 FreeSans 320 0 0 0 x2.x5[5].CBOT
flabel space 10503 -2257 10563 -1225 0 FreeSans 320 0 0 0 x2.x5[5].CTOP
flabel space 10336 -1228 10370 -1194 0 FreeSans 320 0 0 0 x2.x5[5].SW
flabel metal4 10641 -1573 10667 -1541 0 FreeSans 320 0 0 0 x2.x5[5].x1.CBOT
flabel metal4 10523 -2163 10549 -2131 0 FreeSans 320 0 0 0 x2.x5[5].x1.CTOP
flabel nwell 10507 -1955 10677 -1785 0 FreeSans 320 0 0 0 x2.x5[5].x1.SUB
flabel space 9903 -1955 10073 -1785 0 FreeSans 320 0 0 0 x2.x5[4].SUB
flabel space 9897 -2195 9957 -1161 0 FreeSans 320 0 0 0 x2.x5[4].CBOT
flabel space 10017 -2257 10077 -1225 0 FreeSans 320 0 0 0 x2.x5[4].CTOP
flabel space 10210 -1228 10244 -1194 0 FreeSans 320 0 0 0 x2.x5[4].SW
flabel metal4 9913 -1573 9939 -1541 0 FreeSans 320 0 0 0 x2.x5[4].x1.CBOT
flabel metal4 10031 -2163 10057 -2131 0 FreeSans 320 0 0 0 x2.x5[4].x1.CTOP
flabel nwell 9903 -1955 10073 -1785 0 FreeSans 320 0 0 0 x2.x5[4].x1.SUB
flabel space 9295 -1955 9465 -1785 0 FreeSans 320 0 0 0 x2.x5[3].SUB
flabel space 9411 -2195 9471 -1161 0 FreeSans 320 0 0 0 x2.x5[3].CBOT
flabel space 9291 -2257 9351 -1225 0 FreeSans 320 0 0 0 x2.x5[3].CTOP
flabel space 9124 -1228 9158 -1194 0 FreeSans 320 0 0 0 x2.x5[3].SW
flabel metal4 9429 -1573 9455 -1541 0 FreeSans 320 0 0 0 x2.x5[3].x1.CBOT
flabel metal4 9311 -2163 9337 -2131 0 FreeSans 320 0 0 0 x2.x5[3].x1.CTOP
flabel nwell 9295 -1955 9465 -1785 0 FreeSans 320 0 0 0 x2.x5[3].x1.SUB
flabel space 8691 -1955 8861 -1785 0 FreeSans 320 0 0 0 x2.x5[2].SUB
flabel space 8685 -2195 8745 -1161 0 FreeSans 320 0 0 0 x2.x5[2].CBOT
flabel space 8805 -2257 8865 -1225 0 FreeSans 320 0 0 0 x2.x5[2].CTOP
flabel space 8998 -1228 9032 -1194 0 FreeSans 320 0 0 0 x2.x5[2].SW
flabel metal4 8701 -1573 8727 -1541 0 FreeSans 320 0 0 0 x2.x5[2].x1.CBOT
flabel metal4 8819 -2163 8845 -2131 0 FreeSans 320 0 0 0 x2.x5[2].x1.CTOP
flabel nwell 8691 -1955 8861 -1785 0 FreeSans 320 0 0 0 x2.x5[2].x1.SUB
flabel space 8083 -1955 8253 -1785 0 FreeSans 320 0 0 0 x2.x5[1].SUB
flabel space 8199 -2195 8259 -1161 0 FreeSans 320 0 0 0 x2.x5[1].CBOT
flabel space 8079 -2257 8139 -1225 0 FreeSans 320 0 0 0 x2.x5[1].CTOP
flabel space 7912 -1228 7946 -1194 0 FreeSans 320 0 0 0 x2.x5[1].SW
flabel metal4 8217 -1573 8243 -1541 0 FreeSans 320 0 0 0 x2.x5[1].x1.CBOT
flabel metal4 8099 -2163 8125 -2131 0 FreeSans 320 0 0 0 x2.x5[1].x1.CTOP
flabel nwell 8083 -1955 8253 -1785 0 FreeSans 320 0 0 0 x2.x5[1].x1.SUB
flabel space 7479 -1955 7649 -1785 0 FreeSans 320 0 0 0 x2.x5[0].SUB
flabel space 7473 -2195 7533 -1161 0 FreeSans 320 0 0 0 x2.x5[0].CBOT
flabel space 7593 -2257 7653 -1225 0 FreeSans 320 0 0 0 x2.x5[0].CTOP
flabel space 7786 -1228 7820 -1194 0 FreeSans 320 0 0 0 x2.x5[0].SW
flabel metal4 7489 -1573 7515 -1541 0 FreeSans 320 0 0 0 x2.x5[0].x1.CBOT
flabel metal4 7607 -2163 7633 -2131 0 FreeSans 320 0 0 0 x2.x5[0].x1.CTOP
flabel nwell 7479 -1955 7649 -1785 0 FreeSans 320 0 0 0 x2.x5[0].x1.SUB
flabel metal1 6726 1929 7394 1976 0 FreeSans 320 0 0 0 x1.IN
flabel metal1 13202 1927 13384 1973 0 FreeSans 320 0 0 0 x1.OUT
flabel metal4 6750 2671 7212 3281 0 FreeSans 320 0 0 0 x1.VDD
flabel metal4 6768 622 7198 2061 0 FreeSans 320 0 0 0 x1.VSS
flabel metal1 6689 2312 6827 2346 0 FreeSans 320 0 0 0 x1.code[3]
flabel metal1 6707 1726 7101 1773 0 FreeSans 320 0 0 0 x1.code_offset
flabel metal1 12460 600 12518 1756 0 FreeSans 320 0 0 0 x1.code[0]
flabel metal1 11604 601 11662 1778 0 FreeSans 320 0 0 0 x1.code[1]
flabel metal1 9178 601 9236 1778 0 FreeSans 320 0 0 0 x1.code[2]
flabel poly 7314 1725 7416 1755 0 FreeSans 320 0 0 0 x1.x9.input_stack
flabel space 7428 1638 7462 1698 0 FreeSans 320 0 0 0 x1.x9.output_stack
flabel space 7428 672 7462 732 0 FreeSans 320 0 0 0 x1.x9.vss
flabel space 8020 762 8080 1796 0 FreeSans 320 0 0 0 x1.x7.CBOT
flabel space 8140 700 8200 1732 0 FreeSans 320 0 0 0 x1.x7.CTOP
flabel space 8026 1002 8196 1172 0 FreeSans 320 0 0 0 x1.x7.SUB
flabel space 8334 1738 8368 1772 0 FreeSans 320 0 0 0 x1.x7.SW
flabel metal4 8036 1384 8062 1416 0 FreeSans 320 0 0 0 x1.x7.x2.CBOT
flabel metal4 8154 794 8180 826 0 FreeSans 320 0 0 0 x1.x7.x2.CTOP
flabel pwell 8026 1002 8196 1172 0 FreeSans 320 0 0 0 x1.x7.x2.SUB
flabel space 8752 762 8812 1796 0 FreeSans 320 0 0 0 x1.x4[3].CBOT
flabel space 8872 700 8932 1732 0 FreeSans 320 0 0 0 x1.x4[3].CTOP
flabel space 8758 1002 8928 1172 0 FreeSans 320 0 0 0 x1.x4[3].SUB
flabel space 9066 1738 9100 1772 0 FreeSans 320 0 0 0 x1.x4[3].SW
flabel metal4 8768 1384 8794 1416 0 FreeSans 320 0 0 0 x1.x4[3].x2.CBOT
flabel metal4 8886 794 8912 826 0 FreeSans 320 0 0 0 x1.x4[3].x2.CTOP
flabel pwell 8758 1002 8928 1172 0 FreeSans 320 0 0 0 x1.x4[3].x2.SUB
flabel space 9478 762 9538 1796 0 FreeSans 320 0 0 0 x1.x4[2].CBOT
flabel space 9358 700 9418 1732 0 FreeSans 320 0 0 0 x1.x4[2].CTOP
flabel space 9362 1002 9532 1172 0 FreeSans 320 0 0 0 x1.x4[2].SUB
flabel space 9190 1738 9224 1772 0 FreeSans 320 0 0 0 x1.x4[2].SW
flabel metal4 9496 1384 9522 1416 0 FreeSans 320 0 0 0 x1.x4[2].x2.CBOT
flabel metal4 9378 794 9404 826 0 FreeSans 320 0 0 0 x1.x4[2].x2.CTOP
flabel pwell 9362 1002 9532 1172 0 FreeSans 320 0 0 0 x1.x4[2].x2.SUB
flabel space 9964 762 10024 1796 0 FreeSans 320 0 0 0 x1.x4[1].CBOT
flabel space 10084 700 10144 1732 0 FreeSans 320 0 0 0 x1.x4[1].CTOP
flabel space 9970 1002 10140 1172 0 FreeSans 320 0 0 0 x1.x4[1].SUB
flabel space 10278 1738 10312 1772 0 FreeSans 320 0 0 0 x1.x4[1].SW
flabel metal4 9980 1384 10006 1416 0 FreeSans 320 0 0 0 x1.x4[1].x2.CBOT
flabel metal4 10098 794 10124 826 0 FreeSans 320 0 0 0 x1.x4[1].x2.CTOP
flabel pwell 9970 1002 10140 1172 0 FreeSans 320 0 0 0 x1.x4[1].x2.SUB
flabel space 10690 762 10750 1796 0 FreeSans 320 0 0 0 x1.x4[0].CBOT
flabel space 10570 700 10630 1732 0 FreeSans 320 0 0 0 x1.x4[0].CTOP
flabel space 10574 1002 10744 1172 0 FreeSans 320 0 0 0 x1.x4[0].SUB
flabel space 10402 1738 10436 1772 0 FreeSans 320 0 0 0 x1.x4[0].SW
flabel metal4 10708 1384 10734 1416 0 FreeSans 320 0 0 0 x1.x4[0].x2.CBOT
flabel metal4 10590 794 10616 826 0 FreeSans 320 0 0 0 x1.x4[0].x2.CTOP
flabel pwell 10574 1002 10744 1172 0 FreeSans 320 0 0 0 x1.x4[0].x2.SUB
flabel space 11302 762 11362 1796 0 FreeSans 320 0 0 0 x1.x3[1].CBOT
flabel space 11422 700 11482 1732 0 FreeSans 320 0 0 0 x1.x3[1].CTOP
flabel space 11308 1002 11478 1172 0 FreeSans 320 0 0 0 x1.x3[1].SUB
flabel space 11616 1738 11650 1772 0 FreeSans 320 0 0 0 x1.x3[1].SW
flabel metal4 11318 1384 11344 1416 0 FreeSans 320 0 0 0 x1.x3[1].x2.CBOT
flabel metal4 11436 794 11462 826 0 FreeSans 320 0 0 0 x1.x3[1].x2.CTOP
flabel pwell 11308 1002 11478 1172 0 FreeSans 320 0 0 0 x1.x3[1].x2.SUB
flabel space 12028 762 12088 1796 0 FreeSans 320 0 0 0 x1.x3[0].CBOT
flabel space 11908 700 11968 1732 0 FreeSans 320 0 0 0 x1.x3[0].CTOP
flabel space 11912 1002 12082 1172 0 FreeSans 320 0 0 0 x1.x3[0].SUB
flabel space 11740 1738 11774 1772 0 FreeSans 320 0 0 0 x1.x3[0].SW
flabel metal4 12046 1384 12072 1416 0 FreeSans 320 0 0 0 x1.x3[0].x2.CBOT
flabel metal4 11928 794 11954 826 0 FreeSans 320 0 0 0 x1.x3[0].x2.CTOP
flabel pwell 11912 1002 12082 1172 0 FreeSans 320 0 0 0 x1.x3[0].x2.SUB
flabel space 12760 762 12820 1796 0 FreeSans 320 0 0 0 x1.x2.CBOT
flabel space 12640 700 12700 1732 0 FreeSans 320 0 0 0 x1.x2.CTOP
flabel space 12644 1002 12814 1172 0 FreeSans 320 0 0 0 x1.x2.SUB
flabel space 12472 1738 12506 1772 0 FreeSans 320 0 0 0 x1.x2.SW
flabel metal4 12778 1384 12804 1416 0 FreeSans 320 0 0 0 x1.x2.x2.CBOT
flabel metal4 12660 794 12686 826 0 FreeSans 320 0 0 0 x1.x2.x2.CTOP
flabel pwell 12644 1002 12814 1172 0 FreeSans 320 0 0 0 x1.x2.x2.SUB
flabel locali 6915 2382 6949 2416 0 FreeSans 340 0 0 0 x1.x1.Y
flabel locali 6915 2314 6949 2348 0 FreeSans 340 0 0 0 x1.x1.Y
flabel locali 6823 2314 6857 2348 0 FreeSans 340 0 0 0 x1.x1.A
flabel metal1 6780 2076 6814 2110 0 FreeSans 200 0 0 0 x1.x1.VGND
flabel metal1 6780 2620 6814 2654 0 FreeSans 200 0 0 0 x1.x1.VPWR
rlabel comment 6751 2093 6751 2093 4 x1.x1.inv_1
rlabel metal1 6751 2045 7027 2141 1 x1.x1.VGND
rlabel metal1 6751 2589 7027 2685 1 x1.x1.VPWR
flabel pwell 6780 2076 6814 2110 0 FreeSans 200 0 0 0 x1.x1.VNB
flabel nwell 6780 2620 6814 2654 0 FreeSans 200 0 0 0 x1.x1.VPB
flabel locali 7013 2382 7047 2416 0 FreeSans 340 0 0 0 x1.x5.Y
flabel locali 7013 2314 7047 2348 0 FreeSans 340 0 0 0 x1.x5.Y
flabel locali 7105 2314 7139 2348 0 FreeSans 340 0 0 0 x1.x5.A
flabel metal1 7148 2076 7182 2110 0 FreeSans 200 0 0 0 x1.x5.VGND
flabel metal1 7148 2620 7182 2654 0 FreeSans 200 0 0 0 x1.x5.VPWR
rlabel comment 7211 2093 7211 2093 6 x1.x5.inv_1
rlabel metal1 6935 2045 7211 2141 1 x1.x5.VGND
rlabel metal1 6935 2589 7211 2685 1 x1.x5.VPWR
flabel pwell 7148 2076 7182 2110 0 FreeSans 200 0 0 0 x1.x5.VNB
flabel nwell 7148 2620 7182 2654 0 FreeSans 200 0 0 0 x1.x5.VPB
flabel metal1 7358 2382 7392 2416 0 FreeSans 320 0 0 0 x1.x8.input_stack
flabel space 7402 3165 7436 3225 0 FreeSans 320 0 0 0 x1.x8.vdd
flabel space 7402 2475 7436 2535 0 FreeSans 320 0 0 0 x1.x8.output_stack
flabel space 7672 2733 7842 2903 0 FreeSans 320 0 0 0 x1.x6.SUB
flabel space 7666 2109 7726 3143 0 FreeSans 320 0 0 0 x1.x6.CBOT
flabel space 7786 2173 7846 3205 0 FreeSans 320 0 0 0 x1.x6.CTOP
flabel space 7979 2142 8013 2176 0 FreeSans 320 0 0 0 x1.x6.SW
flabel metal4 7682 2489 7708 2521 0 FreeSans 320 0 0 0 x1.x6.x1.CBOT
flabel metal4 7800 3079 7826 3111 0 FreeSans 320 0 0 0 x1.x6.x1.CTOP
flabel nwell 7672 2733 7842 2903 0 FreeSans 320 0 0 0 x1.x6.x1.SUB
flabel space 8404 2733 8574 2903 0 FreeSans 320 0 0 0 x1.x5[7].SUB
flabel space 8398 2109 8458 3143 0 FreeSans 320 0 0 0 x1.x5[7].CBOT
flabel space 8518 2173 8578 3205 0 FreeSans 320 0 0 0 x1.x5[7].CTOP
flabel space 8711 2142 8745 2176 0 FreeSans 320 0 0 0 x1.x5[7].SW
flabel metal4 8414 2489 8440 2521 0 FreeSans 320 0 0 0 x1.x5[7].x1.CBOT
flabel metal4 8532 3079 8558 3111 0 FreeSans 320 0 0 0 x1.x5[7].x1.CTOP
flabel nwell 8404 2733 8574 2903 0 FreeSans 320 0 0 0 x1.x5[7].x1.SUB
flabel space 9008 2733 9178 2903 0 FreeSans 320 0 0 0 x1.x5[6].SUB
flabel space 9124 2109 9184 3143 0 FreeSans 320 0 0 0 x1.x5[6].CBOT
flabel space 9004 2173 9064 3205 0 FreeSans 320 0 0 0 x1.x5[6].CTOP
flabel space 8837 2142 8871 2176 0 FreeSans 320 0 0 0 x1.x5[6].SW
flabel metal4 9142 2489 9168 2521 0 FreeSans 320 0 0 0 x1.x5[6].x1.CBOT
flabel metal4 9024 3079 9050 3111 0 FreeSans 320 0 0 0 x1.x5[6].x1.CTOP
flabel nwell 9008 2733 9178 2903 0 FreeSans 320 0 0 0 x1.x5[6].x1.SUB
flabel space 9616 2733 9786 2903 0 FreeSans 320 0 0 0 x1.x5[5].SUB
flabel space 9610 2109 9670 3143 0 FreeSans 320 0 0 0 x1.x5[5].CBOT
flabel space 9730 2173 9790 3205 0 FreeSans 320 0 0 0 x1.x5[5].CTOP
flabel space 9923 2142 9957 2176 0 FreeSans 320 0 0 0 x1.x5[5].SW
flabel metal4 9626 2489 9652 2521 0 FreeSans 320 0 0 0 x1.x5[5].x1.CBOT
flabel metal4 9744 3079 9770 3111 0 FreeSans 320 0 0 0 x1.x5[5].x1.CTOP
flabel nwell 9616 2733 9786 2903 0 FreeSans 320 0 0 0 x1.x5[5].x1.SUB
flabel space 10220 2733 10390 2903 0 FreeSans 320 0 0 0 x1.x5[4].SUB
flabel space 10336 2109 10396 3143 0 FreeSans 320 0 0 0 x1.x5[4].CBOT
flabel space 10216 2173 10276 3205 0 FreeSans 320 0 0 0 x1.x5[4].CTOP
flabel space 10049 2142 10083 2176 0 FreeSans 320 0 0 0 x1.x5[4].SW
flabel metal4 10354 2489 10380 2521 0 FreeSans 320 0 0 0 x1.x5[4].x1.CBOT
flabel metal4 10236 3079 10262 3111 0 FreeSans 320 0 0 0 x1.x5[4].x1.CTOP
flabel nwell 10220 2733 10390 2903 0 FreeSans 320 0 0 0 x1.x5[4].x1.SUB
flabel space 10828 2733 10998 2903 0 FreeSans 320 0 0 0 x1.x5[3].SUB
flabel space 10822 2109 10882 3143 0 FreeSans 320 0 0 0 x1.x5[3].CBOT
flabel space 10942 2173 11002 3205 0 FreeSans 320 0 0 0 x1.x5[3].CTOP
flabel space 11135 2142 11169 2176 0 FreeSans 320 0 0 0 x1.x5[3].SW
flabel metal4 10838 2489 10864 2521 0 FreeSans 320 0 0 0 x1.x5[3].x1.CBOT
flabel metal4 10956 3079 10982 3111 0 FreeSans 320 0 0 0 x1.x5[3].x1.CTOP
flabel nwell 10828 2733 10998 2903 0 FreeSans 320 0 0 0 x1.x5[3].x1.SUB
flabel space 11432 2733 11602 2903 0 FreeSans 320 0 0 0 x1.x5[2].SUB
flabel space 11548 2109 11608 3143 0 FreeSans 320 0 0 0 x1.x5[2].CBOT
flabel space 11428 2173 11488 3205 0 FreeSans 320 0 0 0 x1.x5[2].CTOP
flabel space 11261 2142 11295 2176 0 FreeSans 320 0 0 0 x1.x5[2].SW
flabel metal4 11566 2489 11592 2521 0 FreeSans 320 0 0 0 x1.x5[2].x1.CBOT
flabel metal4 11448 3079 11474 3111 0 FreeSans 320 0 0 0 x1.x5[2].x1.CTOP
flabel nwell 11432 2733 11602 2903 0 FreeSans 320 0 0 0 x1.x5[2].x1.SUB
flabel space 12040 2733 12210 2903 0 FreeSans 320 0 0 0 x1.x5[1].SUB
flabel space 12034 2109 12094 3143 0 FreeSans 320 0 0 0 x1.x5[1].CBOT
flabel space 12154 2173 12214 3205 0 FreeSans 320 0 0 0 x1.x5[1].CTOP
flabel space 12347 2142 12381 2176 0 FreeSans 320 0 0 0 x1.x5[1].SW
flabel metal4 12050 2489 12076 2521 0 FreeSans 320 0 0 0 x1.x5[1].x1.CBOT
flabel metal4 12168 3079 12194 3111 0 FreeSans 320 0 0 0 x1.x5[1].x1.CTOP
flabel nwell 12040 2733 12210 2903 0 FreeSans 320 0 0 0 x1.x5[1].x1.SUB
flabel space 12644 2733 12814 2903 0 FreeSans 320 0 0 0 x1.x5[0].SUB
flabel space 12760 2109 12820 3143 0 FreeSans 320 0 0 0 x1.x5[0].CBOT
flabel space 12640 2173 12700 3205 0 FreeSans 320 0 0 0 x1.x5[0].CTOP
flabel space 12473 2142 12507 2176 0 FreeSans 320 0 0 0 x1.x5[0].SW
flabel metal4 12778 2489 12804 2521 0 FreeSans 320 0 0 0 x1.x5[0].x1.CBOT
flabel metal4 12660 3079 12686 3111 0 FreeSans 320 0 0 0 x1.x5[0].x1.CTOP
flabel nwell 12644 2733 12814 2903 0 FreeSans 320 0 0 0 x1.x5[0].x1.SUB
<< end >>
