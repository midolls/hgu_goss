* NGSPICE file created from hgu_sarlogic_8bit_logic_flat.ext - technology: sky130A

.subckt hgu_sarlogic_8bit_logic_flat sel_bit[0] sel_bit[1] reset eob comparator_out
+ D[7] D[5] check[0] check[5] check[1] check[4] check[2] check[3] D[2] D[1] D[4] D[0]
+ clk_sar D[6] D[3] check[6] VSS VDD
X0 VDD a_10680_2340# D[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1 VDD a_8289_4086# check[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 VDD D[0] a_8236_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3 VDD a_2389_5648# eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X4 a_12030_3213# a_11856_3239# a_12146_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X5 a_4971_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_2147_5083# a_1682_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X7 a_1822_4801# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X8 a_11330_2340# a_11628_2640# a_11564_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X9 VSS a_12030_3213# a_12737_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_4213_3239# a_4367_3213# a_4073_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 a_8591_4801# check[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_9710_4296# a_9238_4086# a_9954_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X13 VSS x30.Q_N a_7185_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X14 VDD a_11250_4775# a_11160_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X15 VSS a_5992_4086# x45.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 a_3599_2340# a_3912_2366# a_4018_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X17 x72.Q_N a_7246_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X18 VSS x27.Q_N a_4018_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X19 a_4854_3213# x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X20 a_7072_3239# a_5844_3239# a_6930_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X21 a_9442_4086# a_8697_4112# a_9578_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X22 VSS x4.X a_9151_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VDD a_7246_3213# a_7158_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X24 VDD a_5897_4086# check[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X25 a_11089_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X26 a_4793_2366# a_4925_2550# a_4657_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 VDD x75.Q a_5844_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_6978_4801# a_6466_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_4388_2732# a_3599_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X30 a_2788_5674# check[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X31 a_10794_3239# a_10628_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 VSS D[0] a_8236_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VDD x4.X a_4368_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X34 a_9465_4801# a_8403_4801# a_9370_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X35 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 a_12048_4394# a_11089_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X37 a_9101_3521# a_8683_3605# a_8857_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X38 a_7247_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X39 VDD a_6846_4086# a_6845_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X40 VSS x20.Q_N a_1626_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X41 D[2] a_12737_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X42 a_11250_4775# a_11076_5167# a_11390_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X43 a_4680_3239# a_3452_3239# a_4538_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X44 a_2479_2648# a_1520_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X45 VDD a_4854_3213# a_4766_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X46 a_11184_4801# a_10795_4801# a_11076_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X47 VSS a_1338_5674# x5.X VSS sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X48 a_2784_5996# check[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X49 a_4593_4112# a_4453_4386# a_4155_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X50 a_1996_2732# a_1207_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X51 a_7181_3239# a_5844_3239# a_7072_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X52 a_6198_3239# comparator_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X53 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X54 a_2265_2340# a_1520_2366# a_2401_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X55 a_12031_4775# a_11857_4801# a_12147_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X56 VSS x75.Q a_5844_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 VDD VDD a_1976_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VSS a_7050_4086# a_6985_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X59 a_1762_2340# a_2060_2640# a_1996_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X60 VDD check[1] a_2969_6040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X61 a_2883_5674# a_2853_5648# a_2788_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X62 a_7562_4478# a_7050_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X63 a_10775_2340# a_11088_2366# a_11194_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X64 a_6504_2648# a_6304_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X65 a_4214_4801# a_4368_4775# a_4074_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X66 VSS x36.Q_N a_11194_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X67 a_10794_3239# a_10628_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 a_4855_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X70 a_7073_4801# a_5845_4801# a_6931_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 VDD a_4454_4086# a_4453_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X72 VDD a_7247_4775# a_7159_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X73 x4.A a_897_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 x30.Q_N a_7247_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X75 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X76 a_12345_2732# a_11833_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X77 VSS check[0] a_5372_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X78 a_8803_4112# a_8939_4086# a_8384_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X79 VSS x4.X a_9152_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X80 a_3806_3239# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X81 VDD x20.Q_N a_1207_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X82 VSS check[1] a_2993_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X83 VSS VDD a_8803_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X84 VSS a_10776_4086# x39.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X85 a_6291_3605# a_5844_3239# a_6198_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X86 x75.Q_N a_4854_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X87 VSS x5.X a_8237_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X88 VSS a_6465_3213# a_6399_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X89 a_1822_4801# a_1976_4775# a_1682_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X90 VDD a_10775_2340# x63.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X91 a_9102_5083# a_8684_5167# a_8858_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X92 a_11856_3239# a_10628_3239# a_11714_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X93 a_4681_4801# a_3453_4801# a_4539_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X94 VDD a_4855_4775# a_4767_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X95 a_9953_2366# a_9441_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X96 check[3] a_12738_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X97 a_1112_2340# a_1207_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X98 a_11769_4112# a_11629_4386# a_11331_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X99 a_2579_4801# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X100 a_4155_4086# a_4453_4386# a_4389_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X101 a_7480_3521# a_7072_3239# a_7246_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X102 VSS VDD a_9578_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X103 a_5992_4086# a_6305_4112# a_6411_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X104 VDD comparator_out a_12547_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X105 a_6199_4801# check[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X106 a_7182_4801# a_5845_4801# a_7073_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X107 VSS VDD a_6411_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X108 VDD x4.X a_6759_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X109 x33.Q_N a_9639_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X110 VSS x27.Q_N a_4793_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X111 a_3899_3605# a_3452_3239# a_3806_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X112 VSS x5.X a_5845_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X113 D[1] a_10345_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X114 a_6710_5083# a_6292_5167# a_6466_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X115 a_11195_4112# a_11331_4086# a_10776_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X116 a_6375_3605# a_5844_3239# a_6291_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X117 a_2969_6040# a_2853_5648# a_2883_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 a_8288_2340# a_8383_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X119 a_10795_4801# a_10629_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X120 a_7050_4086# a_6305_4112# a_7186_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X121 a_11965_3239# a_10628_3239# a_11856_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X122 a_12102_4296# a_11629_4386# a_12346_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X123 VSS a_2463_4775# a_3170_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X124 a_11970_4112# a_12102_4296# a_11834_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X125 VDD a_3505_4086# x48.Q VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X126 a_8590_3239# comparator_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X127 VDD VSS a_3452_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X128 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_4113_4394# a_3913_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X130 VSS a_11834_4086# a_11769_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X131 a_3807_4801# x27.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X132 a_4790_4801# a_3453_4801# a_4681_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X133 VSS x20.Q_N a_2401_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X134 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X135 a_11564_2366# a_10775_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X136 a_7763_2366# a_6844_2640# a_7317_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_11714_3521# a_11249_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X138 a_11857_4801# a_10629_4801# a_11715_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X139 x4.A a_897_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X140 a_6292_5167# a_5845_4801# a_6199_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X141 VDD a_1207_2340# x51.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X142 a_3983_3605# a_3452_3239# a_3899_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X143 a_2389_5648# a_3258_5648# a_2883_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X144 a_5896_2340# a_5991_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X145 VSS a_6466_4775# a_6400_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X146 a_4658_4086# a_3913_4112# a_4794_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X147 VDD a_2463_4775# a_3170_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X148 a_7481_5083# a_7073_4801# a_7247_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X149 a_9237_2340# D[3] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X150 VDD reset a_621_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X151 a_9173_4112# a_8384_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X152 VDD comparator_out a_2979_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X153 VDD a_11833_2340# a_11766_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X154 VSS VSS a_3452_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X155 VDD a_9442_4086# a_9375_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X156 VDD x30.Q_N a_7049_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X157 a_4317_3521# a_3899_3605# a_4073_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X158 a_6376_5167# a_5845_4801# a_6292_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X159 a_3900_5167# a_3453_4801# a_3807_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X160 VSS a_8383_2340# x60.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X161 a_11249_3213# x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X162 a_1227_4801# a_1061_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 a_4074_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X164 a_8997_3239# x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X165 x5.X a_1338_5674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X166 a_8591_4801# check[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X167 a_11289_4394# a_11089_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X168 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X169 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X170 x75.Q a_5561_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X171 a_11966_4801# a_10629_4801# a_11857_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X172 a_9376_2366# a_9236_2640# a_8938_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X173 eob a_2389_5648# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X174 a_6781_4112# a_5992_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X175 x77.Y eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X176 a_9237_2340# D[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X177 a_11715_5083# a_11250_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X178 x27.Q_N a_4855_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X179 a_3984_5167# a_3453_4801# a_3900_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X180 a_8791_3239# a_8402_3239# a_8683_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X181 a_11089_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X182 a_5991_2340# a_6546_2340# a_6504_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X183 a_11075_3605# a_10794_3239# a_10982_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X184 VDD check[0] a_5372_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X185 VDD a_11629_2340# a_11628_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X186 a_9638_3213# a_9464_3239# a_9754_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X187 a_5088_3521# a_4680_3239# a_4854_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X188 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X189 VDD VDD a_9442_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X190 a_6984_2366# a_6844_2640# a_6546_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X191 VDD x4.X a_4367_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X192 a_7318_4296# a_6846_4086# a_7562_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X193 VSS a_9441_2340# a_9376_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X194 a_4318_5083# a_3900_5167# a_4074_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X195 check[4] a_10346_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X196 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 a_12101_2550# a_11629_2340# a_12345_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 a_12548_4112# a_11629_4386# a_12102_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X199 VSS x5.X a_3453_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X200 a_11250_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X201 a_4453_2340# D[5] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X202 a_3373_5674# a_3258_5648# a_2389_5648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X203 VSS x4.X a_6759_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X204 VSS reset a_621_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X205 a_1762_2340# a_2061_2340# a_1996_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X206 a_9550_3605# a_8402_3239# a_9464_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X207 a_8998_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X208 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 a_7049_2340# a_7317_2550# a_7263_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X210 a_6198_3239# comparator_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X211 VSS comparator_out a_7763_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X212 a_2398_4801# a_1061_4801# a_2289_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X213 VSS a_11629_2340# a_11628_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X214 VDD a_6759_3213# a_7480_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X215 a_3877_5674# a_2853_5648# a_3373_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X216 a_9656_4394# a_8697_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X217 a_7185_2366# a_7317_2550# a_7049_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X218 a_10155_2366# a_9237_2340# a_9709_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X219 a_1926_5083# a_1508_5167# a_1682_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X220 a_9370_4801# a_8858_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X221 a_3504_2340# a_3599_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X222 VDD VDD a_11834_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X223 a_11076_5167# a_10795_4801# a_10983_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X224 a_8792_4801# a_8403_4801# a_8684_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X225 a_5089_5083# a_4681_4801# a_4855_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X226 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 VDD a_2061_2340# a_2060_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X228 a_3671_5674# x48.Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X229 a_4453_2340# D[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X230 a_4657_2340# a_4925_2550# a_4871_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X231 a_3806_3239# VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X232 a_9639_4775# a_9465_4801# a_9755_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X233 VDD a_12030_3213# a_12737_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X234 a_4970_3239# a_4367_3213# a_4854_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X235 a_8857_3213# a_8683_3605# a_8997_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X236 a_3600_4086# a_4155_4086# a_4113_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X237 a_8383_2340# a_8696_2366# a_8802_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X238 VDD a_6465_3213# a_6375_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X239 VSS check[0] a_3877_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X240 VSS a_2463_4775# a_2398_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X241 VSS a_8289_4086# check[1] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X242 x5.A a_1062_5674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X243 VDD check[0] a_3876_6040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X244 a_11390_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X245 VSS a_5991_2340# x57.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X246 a_4590_2732# a_4453_2340# a_4154_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 VDD a_8288_2340# D[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X248 VSS comparator_out a_10155_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X249 a_9953_2732# a_9441_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X250 a_8289_4086# a_8384_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X251 a_2697_5083# a_2289_4801# a_2463_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X252 a_9551_5167# a_8403_4801# a_9465_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 a_9441_2340# a_8696_2366# a_9577_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X254 a_6199_4801# check[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X255 a_11630_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 VSS x4.X a_6760_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X257 a_5170_4112# a_4658_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X258 a_10680_2340# a_10775_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X259 VSS sel_bit[1] a_3258_5648# VSS sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X260 a_9173_4478# a_8384_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X261 VDD sel_bit[1] a_3258_5648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X262 check[6] a_5562_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X263 VDD a_6760_4775# a_7481_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X264 a_4389_4112# a_3600_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X265 a_5372_4112# a_4454_4086# a_4926_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X266 a_9375_4478# a_9238_4086# a_8939_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X267 VSS a_2061_2340# a_2060_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X268 a_6465_3213# a_6291_3605# a_6605_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X269 VSS a_5897_4086# check[0] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X270 a_6399_3239# a_6010_3239# a_6291_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X271 VSS a_3599_2340# x54.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X272 eob a_2389_5648# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X273 VDD x5.X a_1061_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X274 VDD a_5896_2340# D[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X275 VDD x27.Q_N a_3599_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X276 a_11389_3239# a_11543_3213# a_11249_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X277 VDD a_4658_4086# a_4591_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X278 VDD a_9237_2340# a_9236_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X279 a_5897_4086# a_5992_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X280 a_8289_4086# a_8384_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X281 a_6304_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X282 a_3807_4801# x27.D VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X283 a_12146_3239# x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X284 VSS a_12031_4775# a_12738_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X285 a_6781_4478# a_5992_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X286 VSS a_1112_2340# D[7] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X287 a_12146_3239# a_11543_3213# a_12030_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X288 a_6983_4478# a_6846_4086# a_6547_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X289 VDD VDD a_8384_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X290 a_9238_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X291 a_12047_2648# a_11088_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X292 a_6546_2340# a_6844_2640# a_6780_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X293 a_1520_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X294 a_4585_3239# a_4073_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X295 VDD a_6466_4775# a_6376_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X296 VSS a_7049_2340# a_6984_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X297 a_11564_2732# a_10775_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X298 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 a_11766_2732# a_11629_2340# a_11330_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X300 a_11833_2340# a_11088_2366# a_11969_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X301 a_4971_4801# a_4368_4775# a_4855_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X302 a_4155_4086# a_4454_4086# a_4389_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X303 a_10156_4112# a_9237_4386# a_9710_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X304 a_7072_3239# a_6010_3239# a_6977_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X305 a_4007_3239# a_3618_3239# a_3899_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X306 a_8858_4775# a_8684_5167# a_8998_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X307 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VDD x4.X a_11544_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X309 a_6305_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X310 a_4018_2366# a_4154_2340# a_3599_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X311 a_5897_4086# a_5992_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X312 VDD a_12031_4775# a_12738_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X313 a_3912_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X314 a_7158_3605# a_6010_3239# a_7072_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_12346_4112# a_11834_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X316 a_9578_4112# a_9710_4296# a_9442_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X317 a_12548_4112# a_11630_4086# a_12102_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X318 VDD a_8384_4086# x42.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X319 VSS a_9237_2340# a_9236_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X320 a_4925_2550# a_4452_2640# a_5169_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X321 VDD VDD a_5992_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X322 x4.A a_897_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 VSS a_4657_2340# a_4592_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X324 x5.A a_1062_5674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X325 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X326 a_2579_4801# a_1976_4775# a_2463_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X327 VDD x36.Q_N a_10775_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X328 a_4680_3239# a_3618_3239# a_4585_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X329 a_6466_4775# a_6292_5167# a_6606_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X330 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X331 a_3913_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X332 a_1626_2366# a_1762_2340# a_1207_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X333 VSS a_9638_3213# a_10345_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X334 VDD a_9151_3213# a_9101_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X335 a_1112_2340# a_1207_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X336 a_11390_4801# a_11544_4775# a_11250_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X337 VSS a_6846_4086# a_6845_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X338 a_4766_3605# a_3618_3239# a_4680_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 x75.Q_N a_4854_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X340 VDD a_11630_4086# a_11629_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X341 a_2533_2550# a_2060_2640# a_2777_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X342 a_2401_2366# a_2533_2550# a_2265_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X343 a_12147_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X344 VSS check[3] a_12548_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X345 a_12147_4801# a_11544_4775# a_12031_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X346 a_10982_3239# comparator_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X347 a_4586_4801# a_4074_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X348 a_2198_2732# a_2061_2340# a_1762_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X349 a_8857_3213# x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X350 a_8403_4801# a_8237_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X351 a_4008_4801# a_3619_4801# a_3900_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X352 a_7073_4801# a_6011_4801# a_6978_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X353 x66.Q_N a_12030_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X354 VDD a_6759_3213# a_6709_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X355 a_7159_5167# a_6011_4801# a_7073_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X356 a_4454_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X357 VSS a_4454_4086# a_4453_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X358 a_8897_4394# a_8697_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X359 a_12030_3213# x39.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X360 D[1] a_10345_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X361 a_3373_5674# a_2853_5648# a_3648_5972# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X362 a_11331_4086# a_11629_4386# a_11565_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X363 a_11856_3239# a_10794_3239# a_11761_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X364 a_8697_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X365 a_8683_3605# a_8402_3239# a_8590_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X366 D[0] a_7953_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X367 a_6011_4801# a_5845_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X368 VSS x36.Q_N a_11969_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X369 a_4681_4801# a_3619_4801# a_4586_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X370 VDD a_9152_4775# a_9102_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X371 VSS a_3505_4086# x48.Q VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X372 a_4767_5167# a_3619_4801# a_4681_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X373 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X374 VSS VDD a_1976_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X375 a_5170_4478# a_4658_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X376 a_4112_2648# a_3912_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X377 VDD a_3504_2340# D[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X378 VSS a_9639_4775# a_10346_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X379 a_2463_4775# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X380 a_3505_4086# a_3600_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X381 a_4389_4478# a_3600_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X382 VDD comparator_out a_7763_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X383 VSS a_2389_5648# eob VSS sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X384 VDD a_1976_4775# a_2697_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X385 x4.A a_897_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X386 x27.Q_N a_4855_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X387 a_6411_4112# a_6547_4086# a_5992_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X388 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 a_8858_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X390 a_10983_4801# check[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X391 VDD a_6760_4775# a_6710_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X392 a_7318_4296# a_6845_4386# a_7562_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X393 VDD a_9639_4775# a_10346_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X394 a_12031_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X395 a_1720_2648# a_1520_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X396 VSS a_4073_3213# a_4007_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X397 a_3505_4086# a_3600_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X398 VSS a_9638_3213# a_9573_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X399 a_2289_4801# a_1061_4801# a_2147_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X400 a_6845_2340# D[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X401 VDD a_2463_4775# a_2375_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X402 a_7561_2366# a_7049_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X403 a_7763_2366# a_6845_2340# a_7317_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X404 check[4] a_10346_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X405 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X406 VDD a_9441_2340# a_9374_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X407 VSS VDD a_7186_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X408 a_8684_5167# a_8403_4801# a_8591_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X409 a_11857_4801# a_10795_4801# a_11762_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X410 VDD comparator_out a_10155_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X411 a_8938_2340# a_9237_2340# a_9172_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X412 a_6930_3521# a_6465_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X413 VDD a_897_4112# x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 a_3600_4086# a_3913_4112# a_4019_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X415 a_1511_4112# x4.A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X416 VSS VDD a_4019_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X417 a_11288_2648# a_11088_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X418 x75.Q a_5561_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X419 a_12346_4478# a_11834_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X420 x77.Y eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X421 VDD a_9238_4086# a_9237_4386# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X422 a_11493_3521# a_11075_3605# a_11249_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X423 a_3373_5674# sel_bit[1] a_2389_5648# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X424 VDD a_3600_4086# x48.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X425 a_9710_4296# a_9237_4386# a_9954_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X426 a_6845_2340# D[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X427 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 a_6546_2340# a_6845_2340# a_6780_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X429 VSS a_12030_3213# a_11965_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X430 a_11075_3605# a_10628_3239# a_10982_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X431 x69.Q_N a_9638_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X432 a_1415_4801# eob VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X433 VSS a_11249_3213# a_11183_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X434 VDD x5.X a_10629_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X435 x36.Q_N a_12031_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X436 a_5371_2366# a_4452_2640# a_4925_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X437 VDD a_1338_5674# x5.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X438 VSS a_4074_4775# a_4008_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X439 a_2993_5674# sel_bit[0] a_2883_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X440 VSS a_10680_2340# D[3] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VDD check[3] a_12548_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X442 VDD x4.A a_1511_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X443 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 a_12264_3521# a_11856_3239# a_12030_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X445 VSS a_9639_4775# a_9574_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X446 VSS a_2389_5648# eob VSS sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 a_6931_5083# a_6466_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X448 a_10776_4086# a_11089_4112# a_11195_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X449 VDD x4.X a_11543_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X450 a_3619_4801# a_3453_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X451 VSS VDD a_11195_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X452 a_2289_4801# a_1227_4801# a_2194_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X453 check[5] a_7954_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X454 a_11494_5083# a_11076_5167# a_11250_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X455 VDD x27.Q_N a_4657_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X456 a_2979_2366# a_2060_2640# a_2533_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X457 a_11159_3605# a_10628_3239# a_11075_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 check[6] a_5562_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X459 VDD a_7050_4086# a_6983_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X460 a_9754_3239# x42.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X461 a_1508_5167# a_1061_4801# a_1415_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X462 a_9754_3239# a_9151_3213# a_9638_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X463 VSS a_1682_4775# a_1616_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X464 a_9655_2648# a_8696_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X465 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X466 a_8384_4086# a_8939_4086# a_8897_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X467 a_6605_3239# x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X468 a_7764_4112# a_6845_4386# a_7318_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X469 a_3899_3605# a_3618_3239# a_3806_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X470 a_8938_2340# a_9236_2640# a_9172_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X471 a_12547_2366# a_11628_2640# a_12101_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X472 a_9954_4112# a_9442_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X473 x20.Q_N a_2463_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X474 a_11076_5167# a_10629_4801# a_10983_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X475 VSS a_12031_4775# a_11966_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X476 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 VDD x20.Q_N a_2265_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X478 a_1592_5167# a_1061_4801# a_1508_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X479 a_8696_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X480 a_10680_2340# a_10775_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X481 a_5169_2366# a_4657_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X482 a_3599_2340# a_4154_2340# a_4112_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X483 a_12265_5083# a_11857_4801# a_12031_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X484 a_10982_3239# comparator_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X485 a_7246_3213# a_7072_3239# a_7362_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X486 VDD x3.A a_897_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X487 VDD VDD a_7050_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X488 a_4592_2366# a_4452_2640# a_4154_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X489 a_8402_3239# a_8236_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X490 a_4538_3521# a_4073_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X491 a_4926_4296# a_4454_4086# a_5170_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X492 a_10776_4086# a_11331_4086# a_11289_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X493 VDD x36.Q_N a_11833_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X494 a_9709_2550# a_9237_2340# a_9953_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X495 a_2061_2340# D[6] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X496 VSS x5.X a_1061_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X497 a_2777_2366# a_2265_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X498 a_1207_2340# a_1762_2340# a_1720_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X499 a_9755_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X500 a_2979_2366# a_2061_2340# a_2533_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X501 VSS x4.X a_4367_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X502 a_9755_4801# a_9152_4775# a_9639_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X503 a_6606_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X504 a_8802_2366# a_8938_2340# a_8383_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X505 a_11088_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X506 VSS comparator_out a_5371_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X507 VDD a_4657_2340# a_4590_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X508 a_6010_3239# a_5844_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X509 a_11565_4112# a_10776_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X510 VDD a_4367_3213# a_5088_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X511 a_7264_4394# a_6305_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X512 a_8402_3239# a_8236_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X513 VSS x33.Q_N a_8802_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X514 a_9638_3213# x42.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X515 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 VSS a_10775_2340# x63.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X517 x4.X a_1511_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X518 a_11834_4086# a_12102_4296# a_12048_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X519 a_3648_5972# x48.Q VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X520 a_6400_4801# a_6011_4801# a_6292_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X521 a_10983_4801# check[4] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X522 a_6846_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X523 a_11768_2366# a_11628_2640# a_11330_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X524 a_2061_2340# D[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 a_4539_5083# a_4074_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X526 a_2265_2340# a_2533_2550# a_2479_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X527 a_6605_3239# a_6759_3213# a_6465_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X528 a_7247_4775# a_7073_4801# a_7363_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X529 a_11761_3239# a_11249_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X530 a_12102_4296# a_11630_4086# a_12346_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X531 VSS x33.Q_N a_9577_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X532 VDD a_9638_3213# a_10345_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X533 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 a_4872_4394# a_3913_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X535 VSS a_8384_4086# x42.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X536 VDD a_8383_2340# x60.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X537 a_5991_2340# a_6304_2366# a_6410_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X538 a_6010_3239# a_5844_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 VDD a_4073_3213# a_3983_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X540 a_11331_4086# a_11630_4086# a_11565_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X541 VSS x30.Q_N a_6410_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X542 a_9464_3239# a_8236_3239# a_9322_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X543 VDD a_9638_3213# a_9550_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X544 VDD a_897_4112# x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X545 VSS x4.X a_11543_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X546 a_11194_2366# a_11330_2340# a_10775_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X547 a_7561_2732# a_7049_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X548 a_9377_4112# a_9237_4386# a_8939_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X549 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X550 a_7049_2340# a_6304_2366# a_7185_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X551 VSS x4.X a_4368_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X552 a_9238_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_12101_2550# a_11628_2640# a_12345_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X554 eob a_2389_5648# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X555 VDD a_11543_3213# a_12264_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X556 x27.D a_3170_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X557 VDD a_4368_4775# a_5089_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X558 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X559 a_11969_2366# a_12101_2550# a_11833_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X560 VSS a_11833_2340# a_11768_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X561 a_4073_3213# a_3899_3605# a_4213_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X562 a_9639_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X563 VSS a_7246_3213# a_7953_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X564 VSS a_1207_2340# x51.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X565 a_8403_4801# a_8237_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X566 a_6985_4112# a_6845_4386# a_6547_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X567 a_9573_3239# a_8236_3239# a_9464_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X568 a_11942_3605# a_10794_3239# a_11856_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X569 a_4854_3213# a_4680_3239# a_4970_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X570 a_4657_2340# a_3912_2366# a_4793_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X571 x66.Q_N a_12030_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X572 a_1415_4801# eob VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X573 VSS a_9442_4086# a_9377_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X574 VDD a_12030_3213# a_11942_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X575 a_4591_4478# a_4454_4086# a_4155_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X576 a_4154_2340# a_4452_2640# a_4388_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X577 VDD D[1] a_10628_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X578 a_9954_4478# a_9442_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X579 VDD a_10681_4086# check[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X580 a_8896_2648# a_8696_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X581 VDD a_11249_3213# a_11159_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X582 VDD a_4074_4775# a_3984_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X583 a_11762_4801# a_11250_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X584 a_9322_3521# a_8857_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X585 a_9172_2366# a_8383_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X586 a_9465_4801# a_8237_4801# a_9323_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X587 VSS a_4854_3213# a_5561_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X588 VDD a_9639_4775# a_9551_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X589 a_6011_4801# a_5845_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X590 VDD x4.X a_9152_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X591 VSS check[1] a_7764_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X592 D[0] a_7953_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X593 VSS x4.X a_11544_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X594 VSS a_11630_4086# a_11629_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X595 a_1520_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X596 VDD clk_sar a_1062_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X597 x5.X a_1338_5674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X598 a_7186_4112# a_7318_4296# a_7050_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X599 a_10156_4112# a_9238_4086# a_9710_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X600 VDD a_11544_4775# a_12265_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X601 a_3618_3239# a_3452_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X602 VDD a_5992_4086# x45.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X603 a_8683_3605# a_8236_3239# a_8590_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X604 VDD VDD a_3600_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X605 a_11249_3213# a_11075_3605# a_11389_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X606 x72.Q_N a_7246_3213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X607 VSS a_8857_3213# a_8791_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X608 VDD a_1682_4775# a_1592_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X609 x3.A a_621_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X610 a_6780_2366# a_5991_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X611 VSS a_2265_2340# a_2200_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X612 a_4074_4775# a_3900_5167# a_4214_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X613 VSS D[1] a_10628_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X614 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X615 a_4454_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X616 VSS a_7247_4775# a_7954_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X617 a_6547_4086# a_6845_4386# a_6781_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X618 a_10681_4086# a_10776_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X619 a_11943_5167# a_10795_4801# a_11857_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 a_11088_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X621 a_9872_3521# a_9464_3239# a_9638_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X622 a_3876_6040# sel_bit[0] a_3373_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X623 a_11565_4478# a_10776_4086# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X624 VDD a_1511_4112# x4.X VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X625 a_4794_4112# a_4926_4296# a_4658_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X626 a_4855_4775# a_4681_4801# a_4971_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X627 a_9574_4801# a_8237_4801# a_9465_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X628 a_8384_4086# a_8697_4112# a_8803_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X629 a_11767_4478# a_11630_4086# a_11331_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X630 VDD a_12031_4775# a_11943_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X631 x36.Q_N a_12031_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X632 D[2] a_12737_3239# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X633 a_9323_5083# a_8858_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X634 VSS check[2] a_10156_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X635 VDD a_5991_2340# x57.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X636 a_8767_3605# a_8236_3239# a_8683_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X637 a_3618_3239# a_3452_3239# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X638 a_2194_4801# a_1682_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X639 a_1682_4775# a_1508_5167# a_1822_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X640 VDD a_7247_4775# a_7954_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X641 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X642 a_5169_2732# a_4657_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X643 a_6465_3213# x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X644 VSS a_4855_4775# a_5562_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X645 a_10681_4086# a_10776_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X646 a_1616_4801# a_1227_4801# a_1508_5167# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X647 VDD a_4367_3213# a_4317_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X648 VSS a_897_4112# x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X649 a_6505_4394# a_6305_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X650 a_9709_2550# a_9236_2640# a_9953_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X651 a_2463_4775# a_2289_4801# a_2579_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X652 check[5] a_7954_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X653 VDD VDD a_10776_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X654 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X655 VSS a_3600_4086# x48.Q_N VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X656 VDD a_3599_2340# x54.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X657 a_1207_2340# a_1520_2366# a_1626_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X658 a_8684_5167# a_8237_4801# a_8591_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X659 VSS a_8858_4775# a_8792_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X660 VDD a_4855_4775# a_5562_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X661 a_6305_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X662 a_3373_5674# sel_bit[0] a_3671_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X663 a_2777_2732# a_2265_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X664 a_6291_3605# a_6010_3239# a_6198_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X665 a_2883_5674# sel_bit[0] a_2784_5996# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X666 a_9873_5083# a_9465_4801# a_9639_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X667 VSS x5.X a_10629_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X668 a_11629_2340# D[2] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X669 VSS clk_sar a_1062_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X670 a_2375_5167# a_1227_4801# a_2289_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X671 VDD a_1112_2340# D[7] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X672 x69.Q_N a_9638_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X673 VDD a_10776_4086# x39.Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X674 VDD comparator_out a_5371_2366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X675 a_11834_4086# a_11089_4112# a_11970_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X676 x20.Q_N a_2463_4775# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X677 VDD x5.X a_8237_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X678 x3.A a_621_4112# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X679 VDD x33.Q_N a_9441_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X680 a_8768_5167# a_8237_4801# a_8684_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 a_6709_3521# a_6291_3605# a_6465_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X682 a_4019_4112# a_4155_4086# a_3600_4086# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X683 VSS x4.A a_1511_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X684 a_7317_2550# a_6845_2340# a_7561_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X685 a_6466_4775# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X686 a_3913_4112# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X687 a_3619_4801# a_3453_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X688 VSS a_8288_2340# D[4] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X689 VDD a_11543_3213# a_11493_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X690 a_4926_4296# a_4453_4386# a_5170_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X691 VSS a_9238_4086# a_9237_4386# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X692 a_4789_3239# a_3452_3239# a_4680_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X693 VDD a_4368_4775# a_4318_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X694 VSS a_11250_4775# a_11184_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X695 VSS a_4658_4086# a_4593_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X696 a_11629_2340# D[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X697 VSS a_7246_3213# a_7181_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X698 VDD x5.X a_5845_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X699 x30.Q_N a_7247_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X700 VDD a_7049_2340# a_6982_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X701 a_5371_2366# a_4453_2340# a_4925_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X702 a_4388_2366# a_3599_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X703 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X704 VSS VDD a_4794_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X705 a_8383_2340# a_8938_2340# a_8896_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X706 a_10795_4801# a_10629_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X707 VDD check[1] a_7764_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X708 a_9442_4086# a_9710_4296# a_9656_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X709 a_6292_5167# a_6011_4801# a_6199_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X710 VSS a_5896_2340# D[5] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X711 eob a_2389_5648# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X712 VDD a_1976_4775# a_1926_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X713 a_11160_5167# a_10629_4801# a_11076_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X714 a_1511_4112# x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X715 a_8288_2340# a_8383_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X716 VSS a_4854_3213# a_4789_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X717 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X718 a_1996_2366# a_1207_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X719 check[3] a_12738_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X720 a_4073_3213# x77.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X721 a_8997_3239# a_9151_3213# a_8857_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X722 a_3900_5167# a_3619_4801# a_3807_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X723 VDD a_11544_4775# a_11494_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X724 a_4154_2340# a_4453_2340# a_4388_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X725 VSS x3.A a_897_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X726 VDD a_6845_2340# a_6844_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X727 x33.Q_N a_9639_4775# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X728 a_9441_2340# a_9709_2550# a_9655_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X729 VDD a_11834_4086# a_11767_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X730 a_5896_2340# a_5991_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X731 VDD a_9151_3213# a_9872_3521# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X732 a_10775_2340# a_11330_2340# a_11288_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X733 a_12345_2366# a_11833_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X734 VDD check[2] a_10156_4112# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X735 a_9577_2366# a_9709_2550# a_9441_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X736 a_12547_2366# a_11629_2340# a_12101_2550# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X737 VSS a_7247_4775# a_7182_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X738 a_9172_2732# a_8383_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X739 VSS VDD a_11970_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X740 a_9374_2732# a_9237_2340# a_8938_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X741 VDD x4.X a_9151_3213# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X742 a_1227_4801# a_1061_4801# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X743 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X744 VDD a_4453_2340# a_4452_2640# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X745 a_2389_5648# sel_bit[1] a_2883_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X746 VDD a_2389_5648# eob VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X747 x27.D a_3170_4801# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X748 VSS a_6845_2340# a_6844_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X749 a_7362_3239# x45.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X750 a_7263_2648# a_6304_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X751 a_7362_3239# a_6759_3213# a_7246_3213# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X752 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X753 a_5992_4086# a_6547_4086# a_6505_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X754 VDD a_8857_3213# a_8767_3605# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X755 a_4213_3239# x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X756 VSS a_4855_4775# a_4790_4801# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X757 a_6780_2732# a_5991_2340# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X758 a_5372_4112# a_4453_4386# a_4926_4296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X759 VDD x33.Q_N a_8383_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X760 a_11833_2340# a_12101_2550# a_12047_2648# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X761 a_6982_2732# a_6845_2340# a_6546_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X762 a_4925_2550# a_4453_2340# a_5169_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X763 a_11330_2340# a_11629_2340# a_11564_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X764 VSS comparator_out a_12547_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X765 VDD x5.A a_1338_5674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X766 VDD x4.X a_6760_4775# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X767 a_8998_4801# a_9152_4775# a_8858_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X768 a_10155_2366# a_9236_2640# a_9709_2550# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X769 a_7562_4112# a_7050_4086# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X770 VDD a_9152_4775# a_9873_5083# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X771 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 a_7764_4112# a_6846_4086# a_7318_4296# VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X773 VSS a_4453_2340# a_4452_2640# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X774 a_6304_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X775 a_9369_3239# a_8857_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X776 a_4970_3239# x77.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X777 a_4871_2648# a_3912_2366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X778 VSS x5.A a_1338_5674# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X779 VSS a_897_4112# x4.A VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X780 a_8939_4086# a_9238_4086# a_9173_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X781 a_8590_3239# comparator_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X782 VDD a_7246_3213# a_7953_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X783 VDD x30.Q_N a_5991_2340# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X784 a_2533_2550# a_2061_2340# a_2777_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X785 a_1682_4775# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X786 VDD x5.X a_3453_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X787 VDD VDD a_4658_4086# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X788 a_7050_4086# a_7318_4296# a_7264_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X789 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X790 a_2200_2366# a_2060_2640# a_1762_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X791 a_2853_5648# sel_bit[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X792 a_2853_5648# sel_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X793 a_8696_2366# x4.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X794 a_6606_4801# a_6760_4775# a_6466_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X795 VSS a_1511_4112# x4.X VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X796 VSS a_3504_2340# D[6] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X797 a_11630_4086# x5.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X798 a_3912_2366# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X799 a_6977_3239# a_6465_3213# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X800 a_6846_4086# x5.X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X801 a_11389_3239# x39.Q_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X802 VDD a_8858_4775# a_8768_5167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X803 a_7363_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X804 a_8939_4086# a_9237_4386# a_9173_4478# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X805 a_7363_4801# a_6760_4775# a_7247_4775# VSS sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X806 a_6547_4086# a_6846_4086# a_6781_4112# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X807 a_9464_3239# a_8402_3239# a_9369_3239# VSS sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X808 VDD a_4854_3213# a_5561_3239# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X809 a_4214_4801# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X810 x4.X a_1511_4112# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 a_4658_4086# a_4926_4296# a_4872_4394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X812 a_8697_4112# x4.X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X813 VSS comparator_out a_2979_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X814 VDD a_2265_2340# a_2198_2732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X815 a_1508_5167# a_1227_4801# a_1415_4801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X816 a_6410_2366# a_6546_2340# a_5991_2340# VSS sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X817 VSS a_10681_4086# check[2] VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X818 a_7317_2550# a_6844_2640# a_7561_2366# VSS sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X819 a_3504_2340# a_3599_2340# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X820 a_11183_3239# a_10794_3239# a_11075_3605# VSS sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X821 a_7246_3213# x45.Q_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
C0 x5.X a_3258_5648# 0.00256f
C1 a_1338_5674# a_1227_4801# 0.00211f
C2 check[2] a_3877_5674# 8.16e-20
C3 comparator_out a_2265_2340# 0.00311f
C4 a_12031_4775# check[3] 0.0678f
C5 x5.X sel_bit[1] 0.0977f
C6 x27.Q_N a_3912_2366# 0.0928f
C7 a_4926_4296# a_5170_4112# 0.00812f
C8 check[2] a_7050_4086# 4.4e-21
C9 x30.Q_N x60.Q_N 8.43e-20
C10 x48.Q a_4453_4386# 1.14e-19
C11 check[3] a_11564_2366# 2.19e-20
C12 a_6011_4801# a_6305_4112# 9.06e-19
C13 a_6466_4775# a_5992_4086# 4.54e-19
C14 a_4794_4112# a_4854_3213# 4.45e-20
C15 VDD a_3373_5674# 0.353f
C16 a_1976_4775# a_2375_5167# 0.00133f
C17 a_1508_5167# a_1822_4801# 0.0258f
C18 a_1415_4801# a_1592_5167# 8.94e-19
C19 check[1] a_8938_2340# 0.00112f
C20 VDD x63.Q_N 0.0716f
C21 x27.Q_N a_6199_4801# 3.25e-20
C22 a_8938_2340# a_8802_2366# 0.0282f
C23 a_8696_2366# a_9655_2648# 1.21e-20
C24 a_9236_2640# a_9374_2732# 1.09e-19
C25 D[4] a_9376_2366# 7.47e-20
C26 a_10628_3239# a_10775_2340# 8.35e-19
C27 x4.X a_5169_2732# 1.17e-19
C28 x4.X a_8236_3239# 0.0456f
C29 VDD a_5992_4086# 0.716f
C30 x4.X a_6977_3239# 4.96e-19
C31 check[1] a_4074_4775# 5.89e-20
C32 a_8591_4801# x33.Q_N 4.33e-22
C33 check[1] x20.Q_N 8.16e-19
C34 x4.X a_7264_4394# 8.47e-19
C35 comparator_out a_8683_3605# 0.0011f
C36 x45.Q_N x72.Q_N 3.9e-19
C37 x27.Q_N a_6410_2366# 8.39e-20
C38 x45.Q_N a_7764_4112# 8.17e-20
C39 a_3453_4801# a_3505_4086# 6.04e-19
C40 a_6547_4086# a_8384_4086# 1.86e-21
C41 a_6845_4386# a_7186_4112# 0.00118f
C42 a_6846_4086# a_6985_4112# 2.56e-19
C43 a_8289_4086# comparator_out 2.05e-21
C44 check[0] a_6198_3239# 0.00621f
C45 x5.A a_1415_4801# 7.6e-20
C46 a_2061_2340# a_2533_2550# 0.15f
C47 a_2060_2640# x51.Q_N 4.18e-21
C48 check[6] a_7182_4801# 1.13e-20
C49 a_1061_4801# a_3619_4801# 2.9e-21
C50 comparator_out a_8696_2366# 0.00714f
C51 a_1227_4801# a_3453_4801# 5.24e-20
C52 a_1338_5674# check[2] 1.12e-19
C53 check[5] a_7763_2366# 0.0034f
C54 x4.X a_1822_4801# 0.0326f
C55 a_1227_4801# a_2194_4801# 0.00126f
C56 a_1061_4801# a_2697_5083# 1.25e-19
C57 clk_sar a_1338_5674# 6.59e-19
C58 a_1062_5674# x5.A 0.136f
C59 a_4454_4086# x48.Q_N 1.07e-19
C60 a_4658_4086# a_4926_4296# 0.205f
C61 eob reset 4.08e-19
C62 check[0] a_7049_2340# 4.27e-19
C63 VDD eob 2.32f
C64 x36.Q_N a_10680_2340# 3.7e-19
C65 a_4155_4086# x77.Y 0.00176f
C66 x5.X x39.Q_N 0.00647f
C67 a_4214_4801# a_4586_4801# 3.34e-19
C68 a_10795_4801# comparator_out 2.89e-21
C69 D[6] x54.Q_N 0.00317f
C70 a_6465_3213# D[0] 1.23e-20
C71 reset x4.A 0.00101f
C72 x4.X a_11288_2648# 0.00102f
C73 a_12101_2550# a_12345_2366# 0.00812f
C74 VDD x4.A 0.787f
C75 a_11089_4112# a_10628_3239# 2.21e-19
C76 a_10776_4086# a_10794_3239# 3.48e-19
C77 a_11390_4801# a_11762_4801# 3.34e-19
C78 x5.X a_6505_4394# 5.63e-19
C79 x75.Q_N a_6010_3239# 2.12e-19
C80 sel_bit[0] a_2883_5674# 0.0666f
C81 x5.X x75.Q 0.0011f
C82 VDD a_4590_2732# 0.0172f
C83 x4.X a_621_4112# 9.87e-20
C84 a_9237_4386# x39.Q_N 2.03e-19
C85 a_4854_3213# x75.Q 0.0108f
C86 check[0] a_3913_4112# 0.00318f
C87 VDD a_7158_3605# 0.00371f
C88 a_7246_3213# a_7763_2366# 2.38e-19
C89 check[6] a_6400_4801# 1.18e-19
C90 check[4] a_10156_4112# 0.00259f
C91 a_4452_2640# a_6845_2340# 2.9e-21
C92 a_4453_2340# a_6844_2640# 4e-20
C93 a_4925_2550# a_6304_2366# 9.52e-21
C94 a_8236_3239# a_9464_3239# 0.0334f
C95 a_8402_3239# a_9638_3213# 0.0264f
C96 a_8857_3213# a_9151_3213# 0.199f
C97 VDD a_6781_4478# 0.00371f
C98 x72.Q_N a_9151_3213# 2.97e-20
C99 x20.Q_N a_2061_2340# 0.0469f
C100 check[2] a_3453_4801# 9.66e-20
C101 x4.X a_8684_5167# 0.00132f
C102 x5.X a_1592_5167# 4.22e-19
C103 check[0] x4.X 0.245f
C104 x33.Q_N a_11088_2366# 8.24e-20
C105 check[2] a_10629_4801# 0.00307f
C106 check[1] a_7953_3239# 0.00311f
C107 a_7363_4801# a_6845_4386# 8.84e-21
C108 a_6845_2340# a_7561_2732# 0.0018f
C109 a_7049_2340# a_7263_2648# 0.0104f
C110 a_6844_2640# a_7763_2366# 0.159f
C111 a_8402_3239# a_9236_2640# 4.04e-20
C112 a_9151_3213# a_8383_2340# 9.06e-19
C113 a_8857_3213# a_8938_2340# 4.18e-20
C114 a_8236_3239# a_9237_2340# 6.52e-20
C115 a_8683_3605# a_8696_2366# 1.71e-19
C116 a_7481_5083# x30.Q_N 2.02e-20
C117 VDD a_1926_5083# 0.0117f
C118 check[4] check[3] 9.63e-20
C119 x42.Q_N a_10345_3239# 3.23e-19
C120 check[1] a_6931_5083# 4.8e-19
C121 x27.Q_N D[6] 0.00313f
C122 x5.A x5.X 0.00793f
C123 x5.X a_4926_4296# 5.33e-19
C124 x48.Q a_4681_4801# 0.00128f
C125 check[3] a_11629_2340# 0.0405f
C126 a_4926_4296# a_4854_3213# 3.74e-20
C127 a_4658_4086# a_4680_3239# 4.33e-20
C128 x77.Y a_4073_3213# 0.201f
C129 a_8383_2340# a_8938_2340# 0.197f
C130 VDD x48.Q_N 0.0812f
C131 x4.X a_4154_2340# 0.00377f
C132 a_10628_3239# a_12264_3521# 1.25e-19
C133 a_11075_3605# a_11389_3239# 0.0258f
C134 a_10794_3239# a_11761_3239# 0.00126f
C135 a_11543_3213# a_11942_3605# 0.00133f
C136 a_6846_4086# D[0] 3.2e-19
C137 VDD a_11970_4112# 0.0326f
C138 a_5844_3239# a_7953_3239# 1.03e-19
C139 comparator_out a_4657_2340# 0.00586f
C140 x27.Q_N a_5991_2340# 1.43e-19
C141 check[5] a_7246_3213# 0.00432f
C142 x4.X a_4538_3521# 0.00211f
C143 a_3453_4801# a_4074_4775# 0.117f
C144 x20.Q_N a_3453_4801# 0.00252f
C145 a_3170_4801# x27.D 0.0749f
C146 check[2] a_9639_4775# 0.0119f
C147 a_2289_4801# a_2398_4801# 0.00707f
C148 a_10681_4086# a_11630_4086# 7e-20
C149 a_2194_4801# x20.Q_N 1.61e-19
C150 a_1207_2340# a_1996_2732# 7.71e-20
C151 a_1520_2366# a_1720_2648# 0.00185f
C152 a_9237_2340# a_11288_2648# 4.06e-20
C153 x4.X a_7263_2648# 2.86e-19
C154 x4.X a_8791_3239# 6.32e-19
C155 a_10629_4801# a_11250_4775# 0.117f
C156 VDD a_8237_4801# 0.81f
C157 comparator_out D[4] 0.00125f
C158 comparator_out a_11249_3213# 4.81e-19
C159 a_897_4112# a_1207_2340# 6.9e-19
C160 a_3913_4112# a_4389_4478# 0.00133f
C161 comparator_out x69.Q_N 1.46e-19
C162 check[5] a_6844_2640# 0.0314f
C163 a_9639_4775# a_9151_3213# 1.08e-22
C164 a_9152_4775# a_9638_3213# 1.06e-20
C165 x5.X x27.D 0.151f
C166 a_4214_4801# a_3600_4086# 1.08e-19
C167 check[0] a_7186_4112# 3.6e-20
C168 a_8403_4801# a_8697_4112# 9.06e-19
C169 a_8858_4775# a_8384_4086# 4.54e-19
C170 a_3258_5648# a_3373_5674# 0.18f
C171 a_2060_2640# x54.Q_N 1.48e-19
C172 a_6010_3239# a_4970_3239# 7.73e-20
C173 a_6465_3213# a_6375_3605# 6.69e-20
C174 a_6291_3605# a_6198_3239# 0.0367f
C175 a_6759_3213# a_7072_3239# 0.124f
C176 sel_bit[1] a_3373_5674# 0.0439f
C177 a_2883_5674# a_2788_5674# 0.00133f
C178 check[3] a_11834_4086# 8.07e-19
C179 x4.X a_4389_4478# 2.12e-19
C180 comparator_out a_10775_2340# 0.00442f
C181 a_10681_4086# D[1] 0.00123f
C182 a_3452_3239# a_4452_2640# 6.01e-20
C183 a_3899_3605# a_3599_2340# 3.9e-20
C184 a_4073_3213# a_3912_2366# 0.0014f
C185 a_5897_4086# a_6845_4386# 9.02e-21
C186 a_5372_4112# a_6846_4086# 3.65e-21
C187 x5.X a_6760_4775# 0.00141f
C188 x27.Q_N a_6846_4086# 1.92e-21
C189 VDD a_2401_2366# 0.00631f
C190 a_5562_4801# a_5561_3239# 9.85e-20
C191 a_5845_4801# a_6199_4801# 0.0663f
C192 a_6292_5167# a_6760_4775# 0.0633f
C193 a_6011_4801# a_7073_4801# 0.137f
C194 check[0] a_4368_4775# 0.00265f
C195 a_4854_3213# a_4680_3239# 0.197f
C196 a_3899_3605# a_3983_3605# 0.00972f
C197 a_4073_3213# a_4317_3521# 0.0104f
C198 a_3618_3239# a_4538_3521# 1.09e-19
C199 D[0] a_8402_3239# 0.00637f
C200 a_7246_3213# a_6844_2640# 3.43e-19
C201 a_6759_3213# a_6845_2340# 2.19e-19
C202 x72.Q_N a_7953_3239# 0.178f
C203 a_8237_4801# a_10983_4801# 3.65e-21
C204 a_9465_4801# a_10795_4801# 2.57e-20
C205 check[2] a_10794_3239# 0.0351f
C206 VDD a_3806_3239# 0.117f
C207 VDD a_7247_4775# 0.72f
C208 x75.Q a_5896_2340# 0.00129f
C209 x5.X a_9238_4086# 0.261f
C210 x33.Q_N D[3] 0.00525f
C211 VDD a_6780_2732# 0.00371f
C212 check[5] x45.Q_N 5.14e-20
C213 a_10776_4086# a_11565_4478# 7.71e-20
C214 a_11089_4112# a_11289_4394# 0.00185f
C215 eob a_3258_5648# 3.1e-19
C216 eob sel_bit[1] 0.317f
C217 VDD a_9322_3521# 0.0163f
C218 a_9151_3213# a_10794_3239# 1.89e-19
C219 a_9638_3213# a_10628_3239# 0.00116f
C220 a_5991_2340# a_7317_2550# 4.7e-22
C221 a_6304_2366# a_7049_2340# 0.199f
C222 a_6546_2340# a_6845_2340# 0.0334f
C223 a_9151_3213# a_9872_3521# 0.00185f
C224 VDD a_9442_4086# 0.487f
C225 sel_bit[1] x4.A 1.56e-20
C226 x4.X a_9377_4112# 6.75e-19
C227 a_8384_4086# a_8997_3239# 1.16e-20
C228 x42.Q_N a_8590_3239# 8.76e-20
C229 x27.Q_N a_2060_2640# 0.00112f
C230 check[6] a_4454_4086# 0.0339f
C231 x4.X x33.Q_N 0.421f
C232 a_8939_4086# a_9442_4086# 0.00187f
C233 a_8384_4086# x42.Q_N 0.154f
C234 a_9237_4386# a_9238_4086# 0.75f
C235 a_8697_4112# a_9710_4296# 0.0633f
C236 a_11089_4112# comparator_out 2.29e-20
C237 a_4855_4775# a_6199_4801# 8.26e-21
C238 clk_sar x3.A 1.29e-20
C239 x5.X a_9755_4801# 2.07e-19
C240 D[4] a_8696_2366# 8.79e-19
C241 x4.X a_6291_3605# 0.0177f
C242 a_8237_4801# a_9323_5083# 0.00907f
C243 a_8403_4801# a_9102_5083# 2.46e-19
C244 check[3] a_12548_4112# 0.159f
C245 a_2853_5648# a_1976_4775# 1.02e-19
C246 VDD a_2398_4801# 6.04e-19
C247 x48.Q a_3648_5972# 0.00114f
C248 x45.Q_N a_7246_3213# 0.144f
C249 a_7318_4296# a_7072_3239# 2.37e-20
C250 a_5844_3239# a_6198_3239# 0.0708f
C251 comparator_out a_7072_3239# 1.93e-19
C252 x27.Q_N a_5371_2366# 0.0318f
C253 x42.Q_N a_9441_2340# 1.11e-19
C254 VDD a_9574_4801# 7.87e-19
C255 a_5992_4086# a_6505_4394# 0.00945f
C256 a_10795_4801# a_11249_3213# 3.18e-21
C257 a_11076_5167# a_10628_3239# 8.3e-21
C258 check[2] check[5] 7.25e-20
C259 a_11249_3213# a_11194_2366# 5.71e-21
C260 a_8938_2340# a_9577_2366# 0.00316f
C261 a_9236_2640# a_9376_2366# 0.00126f
C262 a_8696_2366# a_10775_2340# 6.25e-21
C263 a_9755_4801# a_9237_4386# 8.84e-21
C264 check[1] a_3913_4112# 9.87e-21
C265 x4.X a_6304_2366# 0.112f
C266 a_7318_4296# a_6845_2340# 6.08e-21
C267 x45.Q_N a_6844_2640# 4.61e-20
C268 sel_bit[0] reset 8.49e-21
C269 a_5844_3239# a_7049_2340# 4.77e-19
C270 comparator_out a_6845_2340# 0.182f
C271 VDD sel_bit[0] 1.26f
C272 a_4074_4775# a_4019_4112# 8.14e-21
C273 check[5] a_9151_3213# 8.29e-21
C274 check[4] a_9953_2366# 5.12e-20
C275 check[2] a_10776_4086# 0.0128f
C276 x5.X a_9954_4478# 1.64e-19
C277 a_3900_5167# a_4214_4801# 0.0258f
C278 a_3619_4801# a_4586_4801# 0.00126f
C279 a_3453_4801# a_5089_5083# 1.25e-19
C280 a_4368_4775# a_4767_5167# 0.00133f
C281 x20.Q_N a_4008_4801# 9.98e-20
C282 x5.X a_8998_4801# 9.4e-19
C283 check[1] x4.X 0.262f
C284 a_11330_2340# a_11564_2732# 0.00976f
C285 a_10775_2340# a_11194_2366# 0.0397f
C286 a_11088_2366# a_11766_2732# 0.00652f
C287 x4.X a_8802_2366# 3.78e-20
C288 a_7481_5083# a_8237_4801# 4.06e-20
C289 check[0] x75.Q_N 4.68e-20
C290 VDD a_10156_4112# 0.109f
C291 x4.X a_11389_3239# 0.00267f
C292 a_1682_4775# a_1511_4112# 0.00416f
C293 a_11076_5167# a_11390_4801# 0.0258f
C294 a_10795_4801# a_11762_4801# 0.00126f
C295 comparator_out a_10155_2366# 0.155f
C296 a_10629_4801# a_12265_5083# 1.25e-19
C297 a_11544_4775# a_11943_5167# 0.00133f
C298 x4.X a_9954_4112# 6.39e-19
C299 a_9578_4112# a_9638_3213# 4.45e-20
C300 a_6011_4801# a_6010_3239# 1.39e-19
C301 a_11970_4112# a_12101_2550# 1.72e-22
C302 a_4454_4086# a_6547_4086# 1.67e-21
C303 a_4926_4296# a_5992_4086# 7.98e-21
C304 a_3600_4086# comparator_out 4.69e-20
C305 x5.X a_5562_4801# 0.0294f
C306 a_9237_4386# a_9954_4478# 4.45e-20
C307 a_9238_4086# a_9656_4394# 0.00276f
C308 a_8384_4086# a_9173_4112# 4.2e-20
C309 x33.Q_N a_9464_3239# 0.00295f
C310 VDD a_2777_2732# 0.00561f
C311 check[6] a_6466_4775# 6.88e-19
C312 check[6] a_4367_3213# 1.13e-19
C313 a_5562_4801# a_4854_3213# 3.19e-20
C314 x5.X a_12738_4801# 0.0161f
C315 sel_bit[0] a_3807_4801# 7.41e-20
C316 a_4452_2640# x54.Q_N 5.46e-21
C317 a_4453_2340# a_4925_2550# 0.15f
C318 a_7246_3213# a_9151_3213# 3.71e-20
C319 a_8858_4775# check[4] 9.03e-21
C320 a_1061_4801# a_1682_4775# 0.113f
C321 a_3877_5674# x4.X 4.83e-20
C322 VDD check[6] 0.503f
C323 eob a_1592_5167# 5.68e-19
C324 x4.X a_7050_4086# 0.00987f
C325 x4.X a_5844_3239# 0.0457f
C326 VDD check[3] 0.745f
C327 a_1338_5674# a_1508_5167# 5.69e-20
C328 x33.Q_N a_9237_2340# 0.0469f
C329 check[0] a_5897_4086# 0.116f
C330 VDD a_4592_2366# 0.00111f
C331 D[5] a_7049_2340# 7e-20
C332 a_8236_3239# D[1] 7.04e-20
C333 a_8402_3239# a_10345_3239# 7.94e-21
C334 a_10795_4801# a_11089_4112# 9.06e-19
C335 a_11250_4775# a_10776_4086# 4.54e-19
C336 a_6199_4801# a_6400_4801# 3.67e-19
C337 a_6760_4775# x30.Q_N 0.00766f
C338 a_7247_4775# a_7481_5083# 0.00945f
C339 a_7073_4801# a_6978_4801# 0.00276f
C340 a_4213_3239# a_4585_3239# 3.34e-19
C341 a_1112_2340# a_2061_2340# 1.03e-19
C342 D[7] a_2060_2640# 1.7e-19
C343 D[0] a_9369_3239# 5.51e-20
C344 x5.A eob 0.0017f
C345 x33.Q_N a_11544_4775# 1.35e-20
C346 a_7186_4112# a_6304_2366# 1.26e-20
C347 a_3373_5674# x27.D 5.58e-20
C348 x5.A x4.A 5.23e-21
C349 check[3] D[2] 0.449f
C350 VDD a_8896_2648# 0.00506f
C351 VDD a_11493_3521# 0.00984f
C352 x30.Q_N a_9238_4086# 1.91e-21
C353 a_12102_4296# a_12346_4112# 0.00812f
C354 x39.Q_N a_11970_4112# 0.00173f
C355 a_10794_3239# a_11075_3605# 0.155f
C356 a_10628_3239# a_11543_3213# 0.126f
C357 a_6844_2640# a_8938_2340# 3.87e-20
C358 a_7317_2550# a_7185_2366# 0.0258f
C359 a_6845_2340# a_8696_2366# 3.1e-19
C360 check[5] a_8591_4801# 0.165f
C361 x4.X a_2061_2340# 0.00458f
C362 check[1] a_7186_4112# 2.11e-19
C363 a_10983_4801# check[3] 1.14e-19
C364 x27.Q_N a_4452_2640# 0.569f
C365 check[2] x45.Q_N 2.88e-21
C366 x5.X a_6305_4112# 0.00598f
C367 x77.Y a_4789_3239# 7.87e-19
C368 x48.Q a_4658_4086# 3.93e-19
C369 a_5845_4801# a_6846_4086# 1.15e-19
C370 a_6292_5167# a_6305_4112# 2.81e-19
C371 a_6466_4775# a_6547_4086# 8.83e-20
C372 a_6760_4775# a_5992_4086# 0.0018f
C373 a_6011_4801# a_6845_4386# 7.24e-20
C374 check[3] a_11969_2366# 4.79e-19
C375 a_3452_3239# comparator_out 6.64e-19
C376 a_2289_4801# a_2375_5167# 0.00976f
C377 a_3618_3239# a_5844_3239# 4e-20
C378 VDD a_2788_5674# 6.52e-19
C379 check[1] a_9237_2340# 1.98e-19
C380 check[4] x42.Q_N 6.27e-20
C381 x27.Q_N a_4971_4801# 0.00139f
C382 x60.Q_N a_8896_2648# 2.02e-20
C383 a_9441_2340# a_9374_2732# 9.46e-19
C384 a_8696_2366# a_10155_2366# 4.94e-21
C385 a_9236_2640# a_9655_2648# 2.46e-19
C386 x4.X a_8857_3213# 0.00506f
C387 a_10794_3239# a_11088_2366# 5.94e-19
C388 a_11249_3213# a_10775_2340# 2.5e-19
C389 VDD a_6547_4086# 0.34f
C390 x4.X D[5] 5.17e-19
C391 x4.X x72.Q_N 0.00455f
C392 eob x27.D 4.69e-19
C393 check[1] a_4368_4775# 1.09e-19
C394 x4.X a_7764_4112# 0.00621f
C395 comparator_out a_9638_3213# 0.00374f
C396 check[5] a_7953_3239# 0.0271f
C397 x45.Q_N a_6781_4112# 0.00138f
C398 a_7050_4086# a_7186_4112# 0.07f
C399 a_6846_4086# a_8384_4086# 2.98e-19
C400 a_6845_4386# a_8697_4112# 1.34e-19
C401 a_3619_4801# a_3600_4086# 6.63e-19
C402 a_3453_4801# a_3913_4112# 3.05e-19
C403 x20.Q_N a_3505_4086# 0.00428f
C404 a_11390_4801# a_11543_3213# 1.61e-20
C405 x36.Q_N a_10628_3239# 2.75e-19
C406 a_1207_2340# a_1996_2366# 4.2e-20
C407 a_1520_2366# a_3504_2340# 9.77e-21
C408 a_10680_2340# a_11629_2340# 1.03e-19
C409 x4.X a_8383_2340# 0.111f
C410 comparator_out a_9236_2640# 0.108f
C411 x4.X a_3453_4801# 0.00472f
C412 x4.X a_2194_4801# 0.00509f
C413 a_1227_4801# x20.Q_N 1.52e-19
C414 check[0] x57.Q_N 0.0113f
C415 x4.X a_10629_4801# 0.00428f
C416 x48.Q a_3170_4801# 0.00244f
C417 a_4454_4086# x77.Y 2.63e-20
C418 VDD a_1520_2366# 0.402f
C419 a_3599_2340# a_4112_2648# 0.00945f
C420 a_4214_4801# x27.Q_N 1.45e-19
C421 a_11769_4112# a_11970_4112# 3.34e-19
C422 a_7246_3213# a_7953_3239# 0.0968f
C423 a_6759_3213# D[0] 4.66e-19
C424 x4.X a_11766_2732# 9.81e-19
C425 check[1] a_8897_4394# 9.73e-20
C426 check[2] a_9151_3213# 2.41e-20
C427 comparator_out a_12345_2732# 8.26e-19
C428 a_11089_4112# a_11249_3213# 0.00148f
C429 a_11629_4386# a_10628_3239# 6.5e-20
C430 a_11331_4086# a_10794_3239# 1.07e-20
C431 a_11390_4801# x36.Q_N 4.02e-20
C432 x5.X a_6983_4478# 7.44e-19
C433 sel_bit[0] a_3258_5648# 0.0205f
C434 x5.X x48.Q 0.203f
C435 a_6466_4775# a_6411_4112# 8.14e-21
C436 VDD a_4871_2648# 0.0102f
C437 sel_bit[0] sel_bit[1] 0.428f
C438 a_9442_4086# x39.Q_N 3.43e-20
C439 a_1926_5083# x27.D 3.95e-22
C440 check[0] a_4453_4386# 0.164f
C441 a_8857_3213# a_9464_3239# 0.00187f
C442 a_8236_3239# a_8767_3605# 0.0018f
C443 a_8402_3239# a_8590_3239# 0.163f
C444 a_8683_3605# a_9638_3213# 4.7e-22
C445 VDD a_6411_4112# 0.00996f
C446 a_6605_3239# a_7181_3239# 2.46e-21
C447 x33.Q_N a_10346_4801# 0.184f
C448 a_8384_4086# a_8402_3239# 3.48e-19
C449 a_8697_4112# a_8236_3239# 2.21e-19
C450 x20.Q_N a_2533_2550# 0.153f
C451 a_11089_4112# a_10775_2340# 5.05e-21
C452 check[2] a_4074_4775# 1.07e-19
C453 a_7318_4296# a_7562_4112# 0.00812f
C454 x4.X a_9639_4775# 0.103f
C455 x5.X a_2147_5083# 4.05e-19
C456 x27.D x48.Q_N 8.11e-20
C457 check[2] x20.Q_N 4.28e-20
C458 a_3619_4801# a_3452_3239# 9.04e-19
C459 a_3453_4801# a_3618_3239# 8.16e-19
C460 x33.Q_N a_11628_2640# 1.12e-20
C461 a_7363_4801# a_7050_4086# 7.76e-20
C462 a_6845_2340# D[4] 0.336f
C463 a_7317_2550# a_7561_2732# 0.00972f
C464 a_7049_2340# a_7763_2366# 6.99e-20
C465 a_10345_3239# a_10628_3239# 8.18e-19
C466 a_9151_3213# a_8938_2340# 2.17e-19
C467 a_8857_3213# a_9237_2340# 0.00199f
C468 a_8402_3239# a_9441_2340# 0.00154f
C469 a_9638_3213# a_8696_2366# 8.4e-19
C470 VDD a_2375_5167# 0.00488f
C471 a_4155_4086# a_4452_2640# 4.75e-21
C472 a_3913_4112# a_4453_2340# 1.4e-21
C473 x77.Y a_3504_2340# 3.35e-21
C474 x27.Q_N a_6759_3213# 8.29e-21
C475 x30.Q_N a_7561_2366# 0.00224f
C476 x48.Q a_3984_5167# 5.76e-19
C477 check[3] a_12101_2550# 9.97e-19
C478 x77.Y a_4367_3213# 0.106f
C479 a_8383_2340# a_9237_2340# 0.0492f
C480 a_8696_2366# a_9236_2640# 0.139f
C481 x4.X a_4453_2340# 0.00242f
C482 a_10794_3239# x66.Q_N 3.85e-21
C483 a_11856_3239# a_11942_3605# 0.00976f
C484 a_9754_3239# a_9573_3239# 4.11e-20
C485 x45.Q_N a_7953_3239# 3.23e-19
C486 VDD x77.Y 0.423f
C487 comparator_out D[0] 0.0253f
C488 comparator_out x54.Q_N 0.00122f
C489 a_11195_4112# a_10794_3239# 4.04e-21
C490 x27.Q_N a_6546_2340# 5.08e-20
C491 x4.X a_4213_3239# 0.00268f
C492 x4.X a_4790_4801# 2.39e-19
C493 a_3453_4801# a_4368_4775# 0.125f
C494 a_3619_4801# a_3900_5167# 0.155f
C495 a_10156_4112# x39.Q_N 8.08e-20
C496 x20.Q_N a_4074_4775# 8.63e-20
C497 x5.X a_8403_4801# 0.0201f
C498 a_10776_4086# a_11331_4086# 0.197f
C499 x30.Q_N a_6305_4112# 1.32e-21
C500 x75.Q_N a_5844_3239# 2.94e-19
C501 a_1520_2366# a_2198_2732# 0.00652f
C502 a_1207_2340# a_1626_2366# 0.0397f
C503 a_1762_2340# a_1996_2732# 0.00976f
C504 a_2853_5648# a_2883_5674# 0.224f
C505 a_6760_4775# a_8237_4801# 1.67e-19
C506 check[0] a_6011_4801# 4.88e-19
C507 a_10155_2366# a_10775_2340# 8.26e-21
C508 a_9236_2640# a_11194_2366# 2.19e-20
C509 x4.X a_7763_2366# 8.68e-20
C510 check[1] a_5897_4086# 1.24e-21
C511 x4.X a_10794_3239# 0.0425f
C512 x33.Q_N a_11630_4086# 1.91e-21
C513 x4.X a_9872_3521# 0.00103f
C514 a_10795_4801# a_11076_5167# 0.155f
C515 a_10629_4801# a_11544_4775# 0.125f
C516 VDD a_8858_4775# 0.488f
C517 a_4155_4086# a_4591_4478# 0.00412f
C518 a_3913_4112# a_4019_4112# 0.0552f
C519 a_4454_4086# a_4113_4394# 1.25e-19
C520 a_4453_4386# a_4389_4478# 2.13e-19
C521 comparator_out a_11543_3213# 6.77e-19
C522 check[5] a_7049_2340# 7.15e-20
C523 a_9639_4775# a_9464_3239# 1.33e-23
C524 a_9465_4801# a_9638_3213# 4.82e-21
C525 a_8403_4801# a_9237_4386# 7.24e-20
C526 a_9152_4775# a_8384_4086# 0.0018f
C527 a_8858_4775# a_8939_4086# 8.83e-20
C528 a_8237_4801# a_9238_4086# 1.15e-19
C529 a_8684_5167# a_8697_4112# 2.81e-19
C530 x36.Q_N a_11183_3239# 6.74e-20
C531 D[6] a_2777_2366# 1.54e-19
C532 a_3504_2340# a_3912_2366# 6.04e-19
C533 a_2200_2366# a_2401_2366# 3.34e-19
C534 a_3373_5674# a_3876_6040# 0.00336f
C535 a_6010_3239# a_6709_3521# 2.46e-19
C536 sel_bit[1] a_2788_5674# 2.36e-19
C537 check[3] x39.Q_N 1.04e-19
C538 x4.X a_4019_4112# 0.00642f
C539 a_5561_3239# a_6010_3239# 6.84e-19
C540 comparator_out a_11330_2340# 0.00103f
C541 a_3618_3239# a_4453_2340# 6.38e-20
C542 a_3452_3239# a_4657_2340# 4.77e-19
C543 a_3899_3605# a_4154_2340# 2.41e-20
C544 a_4367_3213# a_3912_2366# 3.36e-20
C545 a_4073_3213# a_4452_2640# 2.68e-19
C546 a_5992_4086# a_6305_4112# 0.272f
C547 a_5897_4086# a_5844_3239# 5.06e-19
C548 x4.X a_4008_4801# 8.46e-20
C549 a_5372_4112# comparator_out 4.39e-20
C550 x4.X x3.A 2.12e-20
C551 x33.Q_N D[1] 3.29e-19
C552 x5.X a_7073_4801# 0.00115f
C553 x4.X a_11184_4801# 8.46e-20
C554 check[6] x75.Q 0.0149f
C555 VDD a_3912_2366# 0.359f
C556 x27.Q_N comparator_out 0.272f
C557 a_6466_4775# a_6199_4801# 6.99e-20
C558 a_6011_4801# a_6376_5167# 4.45e-20
C559 a_4367_3213# a_4317_3521# 1.21e-20
C560 a_6760_4775# a_7247_4775# 0.273f
C561 x5.A sel_bit[0] 0.0448f
C562 a_3618_3239# a_4213_3239# 0.00118f
C563 check[0] a_4681_4801# 0.00122f
C564 a_7953_3239# a_9151_3213# 5.62e-20
C565 D[0] a_8683_3605# 2.17e-19
C566 a_7246_3213# a_7049_2340# 2.52e-19
C567 a_6759_3213# a_7317_2550# 1.62e-19
C568 x36.Q_N comparator_out 0.267f
C569 a_8289_4086# D[0] 0.00123f
C570 check[2] a_11075_3605# 8.1e-20
C571 VDD a_4317_3521# 0.0107f
C572 VDD a_6199_4801# 0.109f
C573 x39.Q_N a_11493_3521# 0.00136f
C574 x4.X check[5] 0.0317f
C575 x5.X a_9710_4296# 6.08e-19
C576 x30.Q_N a_6605_3239# 6.1e-19
C577 VDD a_6410_2366# 4.84e-19
C578 a_11089_4112# a_11767_4478# 0.00652f
C579 a_10776_4086# a_11195_4112# 0.0397f
C580 a_11331_4086# a_11565_4478# 0.00976f
C581 VDD a_8997_3239# 5.47e-21
C582 D[0] a_8696_2366# 3.91e-20
C583 a_9464_3239# a_10794_3239# 3.48e-20
C584 a_9151_3213# a_11075_3605# 4.38e-20
C585 a_8236_3239# a_10982_3239# 3.65e-21
C586 a_6304_2366# x57.Q_N 0.00553f
C587 a_6844_2640# a_7049_2340# 0.153f
C588 a_9638_3213# x69.Q_N 0.124f
C589 VDD x42.Q_N 0.457f
C590 check[2] a_11088_2366# 0.00327f
C591 x4.X a_10776_4086# 0.1f
C592 x30.Q_N a_8288_2340# 2.02e-19
C593 check[4] a_8402_3239# 1.83e-21
C594 a_4019_4112# a_3618_3239# 4.04e-21
C595 a_9238_4086# a_9442_4086# 0.117f
C596 a_8939_4086# x42.Q_N 0.0287f
C597 a_9237_4386# a_9710_4296# 0.155f
C598 a_11629_4386# comparator_out 2.51e-20
C599 VDD a_10680_2340# 0.189f
C600 a_4855_4775# a_4971_4801# 0.0397f
C601 a_4368_4775# a_4790_4801# 2.87e-21
C602 a_8858_4775# a_8803_4112# 8.14e-21
C603 x5.X a_11494_5083# 3.98e-19
C604 VDD a_4113_4394# 0.00555f
C605 sel_bit[0] x27.D 0.00108f
C606 a_7763_2366# a_9237_2340# 3.65e-21
C607 D[4] a_9236_2640# 3.87e-20
C608 x4.X a_7246_3213# 0.115f
C609 a_621_4112# a_897_4112# 0.00202f
C610 D[1] a_11389_3239# 1.6e-19
C611 a_8858_4775# a_9323_5083# 9.46e-19
C612 a_8403_4801# a_9551_5167# 2.13e-19
C613 a_8237_4801# a_8998_4801# 6.04e-20
C614 check[1] a_2463_4775# 0.00193f
C615 VDD a_4539_5083# 0.0172f
C616 a_5992_4086# a_6605_3239# 1.16e-20
C617 x45.Q_N a_6198_3239# 7.37e-20
C618 x48.Q a_3373_5674# 0.0679f
C619 a_6305_4112# a_6781_4478# 0.00133f
C620 VDD a_11715_5083# 0.0163f
C621 a_1976_4775# a_1511_4112# 0.00824f
C622 a_10795_4801# a_11543_3213# 2.05e-21
C623 a_11076_5167# a_11249_3213# 3.52e-21
C624 a_11250_4775# a_11075_3605# 1.33e-23
C625 eob a_1207_2340# 1.75e-19
C626 a_5845_4801# a_7954_4801# 1.03e-19
C627 a_9755_4801# a_9442_4086# 7.76e-20
C628 x4.X a_6844_2640# 0.00904f
C629 a_9236_2640# a_10775_2340# 3.6e-19
C630 a_9441_2340# a_9376_2366# 9.75e-19
C631 a_9237_2340# a_9577_2366# 6.04e-20
C632 check[1] a_4453_4386# 1.28e-20
C633 a_10346_4801# a_10629_4801# 8.18e-19
C634 x4.A a_1207_2340# 9.28e-20
C635 comparator_out a_10345_3239# 0.00106f
C636 x45.Q_N a_7049_2340# 1.11e-19
C637 a_1227_4801# a_1508_5167# 0.151f
C638 a_1061_4801# a_1976_4775# 0.117f
C639 comparator_out a_7317_2550# 0.00825f
C640 a_3505_4086# a_3913_4112# 6.04e-19
C641 x5.X a_10681_4086# 0.0752f
C642 check[2] a_11331_4086# 3.82e-19
C643 a_2579_4801# a_2398_4801# 4.11e-20
C644 a_3619_4801# x27.Q_N 1.18e-19
C645 a_4681_4801# a_4767_5167# 0.00976f
C646 x5.X a_9370_4801# 2.59e-19
C647 D[6] a_3504_2340# 0.103f
C648 a_2060_2640# a_2777_2366# 0.0019f
C649 x4.X a_9953_2732# 1.17e-19
C650 a_11628_2640# a_11766_2732# 1.09e-19
C651 a_11088_2366# a_12047_2648# 1.21e-20
C652 a_11330_2340# a_11194_2366# 0.0282f
C653 x4.X a_12146_3239# 5.65e-19
C654 x30.Q_N a_8403_4801# 2.26e-19
C655 VDD a_9173_4112# 3.55e-19
C656 x4.X a_11761_3239# 4.96e-19
C657 eob x48.Q 0.0102f
C658 x4.X a_3505_4086# 0.0122f
C659 a_10795_4801# x36.Q_N 2.98e-20
C660 comparator_out D[7] 6.69e-20
C661 a_11857_4801# a_11943_5167# 0.00976f
C662 a_9755_4801# a_9574_4801# 4.11e-20
C663 a_4854_3213# a_6010_3239# 3.57e-19
C664 a_4367_3213# a_6465_3213# 4.53e-20
C665 a_6466_4775# a_6465_3213# 2.59e-19
C666 a_6011_4801# a_6291_3605# 8.52e-21
C667 a_6292_5167# a_6010_3239# 1.65e-21
C668 x4.X a_11565_4478# 2.12e-19
C669 VDD a_9873_5083# 0.00506f
C670 check[5] a_9237_2340# 7.28e-22
C671 a_4454_4086# a_6846_4086# 1.37e-19
C672 a_3913_4112# x45.Q_N 1.22e-20
C673 x48.Q x4.A 1.09e-20
C674 x42.Q_N a_8803_4112# 0.0446f
C675 a_9238_4086# a_10156_4112# 0.0663f
C676 a_8939_4086# a_9173_4112# 0.00707f
C677 a_9442_4086# a_9954_4478# 6.69e-20
C678 a_8697_4112# a_9377_4112# 3.73e-19
C679 a_9237_4386# a_10681_4086# 3.59e-19
C680 x36.Q_N a_11194_2366# 0.0102f
C681 a_4794_4112# x77.Y 7.13e-20
C682 VDD D[6] 0.28f
C683 VDD a_6465_3213# 0.308f
C684 check[6] a_6760_4775# 0.00308f
C685 x33.Q_N a_8697_4112# 7.32e-22
C686 a_6759_3213# a_8590_3239# 3.42e-20
C687 a_7246_3213# a_9464_3239# 1.86e-21
C688 a_1227_4801# x4.X 0.311f
C689 a_9639_4775# a_10346_4801# 0.0968f
C690 a_9152_4775# check[4] 0.00456f
C691 eob a_2147_5083# 0.00298f
C692 a_7186_4112# a_7246_3213# 4.45e-20
C693 x4.X x45.Q_N 0.252f
C694 a_4854_3213# a_4793_2366# 1.2e-20
C695 a_2389_5648# a_1976_4775# 1.09e-19
C696 x33.Q_N a_9709_2550# 0.181f
C697 VDD a_5991_2340# 0.561f
C698 check[0] a_4593_4112# 5.07e-20
C699 D[0] D[4] 0.338f
C700 a_8857_3213# D[1] 1.23e-20
C701 a_7073_4801# x30.Q_N 4.49e-19
C702 D[5] x57.Q_N 0.00107f
C703 a_10795_4801# a_11629_4386# 7.24e-20
C704 a_11544_4775# a_10776_4086# 0.0018f
C705 a_11250_4775# a_11331_4086# 8.83e-20
C706 a_11076_5167# a_11089_4112# 2.81e-19
C707 a_10629_4801# a_11630_4086# 1.15e-19
C708 D[7] a_2265_2340# 2.67e-19
C709 check[2] D[3] 0.194f
C710 a_8998_4801# a_9574_4801# 2.46e-21
C711 x33.Q_N a_11857_4801# 1.75e-20
C712 check[1] a_6011_4801# 4e-19
C713 check[2] a_3913_4112# 1.35e-20
C714 check[2] a_11195_4112# 4.22e-19
C715 x33.Q_N a_11768_2366# 2.75e-20
C716 a_3600_4086# a_3452_3239# 8.29e-19
C717 VDD a_2853_5648# 0.413f
C718 VDD a_9374_2732# 0.0163f
C719 VDD a_11942_3605# 0.00371f
C720 a_11249_3213# a_11543_3213# 0.199f
C721 a_10794_3239# a_12030_3213# 0.0264f
C722 a_10628_3239# a_11856_3239# 0.0334f
C723 a_9638_3213# a_10155_2366# 2.38e-19
C724 a_7317_2550# a_8696_2366# 6.06e-21
C725 a_6845_2340# a_9236_2640# 4e-20
C726 a_6844_2640# a_9237_2340# 2.9e-21
C727 x4.X a_2533_2550# 5.96e-19
C728 check[5] a_7363_4801# 8.69e-20
C729 x69.Q_N a_11543_3213# 2.97e-20
C730 a_4794_4112# a_3912_2366# 1.26e-20
C731 check[1] a_8697_4112# 0.00119f
C732 check[2] x4.X 0.258f
C733 x27.Q_N a_4657_2340# 0.179f
C734 x5.X a_6845_4386# 0.0101f
C735 check[4] a_10628_3239# 0.00655f
C736 a_10629_4801# D[1] 1.99e-20
C737 x48.Q x48.Q_N 0.00314f
C738 a_6466_4775# a_6846_4086# 0.00336f
C739 a_6011_4801# a_7050_4086# 0.00221f
C740 a_6760_4775# a_6547_4086# 3.72e-19
C741 a_7247_4775# a_6305_4112# 0.00161f
C742 a_2463_4775# a_3453_4801# 0.00116f
C743 a_1976_4775# a_3619_4801# 2.05e-19
C744 a_8803_4112# a_9173_4112# 4.11e-20
C745 a_9954_4478# a_10156_4112# 8.94e-19
C746 a_4073_3213# comparator_out 3.96e-19
C747 a_6011_4801# a_5844_3239# 9.04e-19
C748 a_1976_4775# a_2697_5083# 0.00185f
C749 a_1508_5167# x20.Q_N 9.58e-20
C750 x77.Y x75.Q 3.59e-19
C751 VDD a_3671_5674# 7.34e-19
C752 check[1] a_9709_2550# 2.04e-19
C753 x27.Q_N a_4007_3239# 6.74e-20
C754 a_9237_2340# a_9953_2732# 0.0018f
C755 a_9441_2340# a_9655_2648# 0.0104f
C756 a_9236_2640# a_10155_2366# 0.159f
C757 x4.X a_9151_3213# 0.111f
C758 a_10794_3239# a_11628_2640# 4.04e-20
C759 a_11543_3213# a_10775_2340# 9.06e-19
C760 a_11249_3213# a_11330_2340# 4.18e-20
C761 a_10628_3239# a_11629_2340# 6.52e-20
C762 a_11075_3605# a_11088_2366# 1.71e-19
C763 VDD a_6846_4086# 0.805f
C764 check[1] a_4681_4801# 3.58e-20
C765 a_2853_5648# a_3807_4801# 1.57e-19
C766 x4.X a_6781_4112# 8.67e-20
C767 comparator_out a_8590_3239# 0.158f
C768 x20.Q_N a_1112_2340# 4.68e-19
C769 a_7318_4296# a_8384_4086# 7.98e-21
C770 a_6846_4086# a_8939_4086# 1.67e-21
C771 x45.Q_N a_7186_4112# 0.00171f
C772 a_4074_4775# a_3913_4112# 0.0025f
C773 a_3900_5167# a_3600_4086# 4.9e-20
C774 a_3453_4801# a_4453_4386# 9.86e-20
C775 check[4] a_9376_2366# 9.3e-20
C776 a_8384_4086# comparator_out 0.00194f
C777 x20.Q_N a_3913_4112# 7.65e-19
C778 x36.Q_N a_11249_3213# 5.36e-19
C779 check[0] a_5170_4112# 8.39e-20
C780 a_1762_2340# a_1996_2366# 0.00707f
C781 a_1520_2366# a_2200_2366# 3.73e-19
C782 a_2060_2640# a_3504_2340# 6.83e-19
C783 check[0] a_5561_3239# 0.0043f
C784 a_6606_4801# check[5] 1.24e-20
C785 a_11250_4775# a_11195_4112# 8.14e-21
C786 x4.X a_8938_2340# 0.00706f
C787 a_10775_2340# a_11330_2340# 0.197f
C788 check[4] a_11390_4801# 1.64e-19
C789 comparator_out a_9441_2340# 0.00598f
C790 x4.X a_4074_4775# 0.00101f
C791 x4.X x20.Q_N 0.274f
C792 x4.X a_11250_4775# 9.45e-19
C793 x36.Q_N a_10775_2340# 0.142f
C794 a_4926_4296# x77.Y 0.00166f
C795 a_5562_4801# check[6] 0.133f
C796 VDD a_2060_2640# 0.329f
C797 a_3912_2366# a_4388_2732# 0.00133f
C798 a_4586_4801# x27.Q_N 1.61e-19
C799 a_7072_3239# D[0] 5.18e-20
C800 x4.X a_12047_2648# 2.86e-19
C801 check[1] a_9375_4478# 6.38e-20
C802 x5.X a_8236_3239# 9.93e-20
C803 check[6] a_4388_2366# 2.11e-20
C804 a_12738_4801# check[3] 0.175f
C805 a_11630_4086# a_10794_3239# 6.04e-20
C806 a_11834_4086# a_10628_3239# 0.00195f
C807 a_11089_4112# a_11543_3213# 3.33e-20
C808 a_11629_4386# a_11249_3213# 0.0015f
C809 a_11331_4086# a_11075_3605# 1.7e-20
C810 a_11762_4801# x36.Q_N 4.04e-20
C811 x30.Q_N a_6010_3239# 4.02e-19
C812 x5.X a_7264_4394# 3.07e-19
C813 sel_bit[0] a_3876_6040# 0.00262f
C814 VDD a_5371_2366# 0.109f
C815 VDD a_8402_3239# 0.275f
C816 check[0] a_4658_4086# 7.37e-19
C817 VDD a_7480_3521# 0.00506f
C818 D[0] a_6845_2340# 0.0271f
C819 a_8402_3239# a_7362_3239# 1.22e-20
C820 a_8857_3213# a_8767_3605# 6.69e-20
C821 a_8683_3605# a_8590_3239# 0.0367f
C822 a_9151_3213# a_9464_3239# 0.124f
C823 a_4453_2340# x57.Q_N 2.94e-19
C824 VDD a_7562_4478# 0.0042f
C825 check[2] a_9237_2340# 6.22e-19
C826 a_8939_4086# a_8402_3239# 1.07e-20
C827 a_9237_4386# a_8236_3239# 6.5e-20
C828 a_8697_4112# a_8857_3213# 0.00148f
C829 check[2] a_4368_4775# 1.3e-19
C830 a_8289_4086# a_8384_4086# 0.0968f
C831 a_6781_4112# a_7186_4112# 2.46e-21
C832 x4.X a_8591_4801# 2.37e-19
C833 x33.Q_N a_11833_2340# 8.49e-21
C834 a_3619_4801# a_5845_4801# 4e-20
C835 a_3453_4801# a_6011_4801# 2.9e-21
C836 a_3619_4801# a_4073_3213# 3.18e-21
C837 a_3900_5167# a_3452_3239# 8.3e-21
C838 x20.Q_N a_3618_3239# 0.0017f
C839 D[1] a_10794_3239# 0.00642f
C840 a_9638_3213# a_9236_2640# 3.43e-19
C841 a_9151_3213# a_9237_2340# 2.19e-19
C842 a_8237_4801# a_8403_4801# 0.751f
C843 x69.Q_N a_10345_3239# 0.178f
C844 x36.Q_N a_11089_4112# 1.39e-22
C845 a_5992_4086# a_6010_3239# 3.48e-19
C846 x48.Q_N a_3599_2340# 9.38e-21
C847 VDD a_1616_4801# 6e-19
C848 a_4453_4386# a_4453_2340# 7.25e-19
C849 a_4454_4086# a_4452_2640# 7.02e-19
C850 a_3600_4086# x54.Q_N 2.32e-20
C851 a_8697_4112# a_8383_2340# 5.05e-21
C852 VDD a_11564_2732# 0.00371f
C853 x77.Y a_4680_3239# 0.16f
C854 a_11543_3213# a_11965_3239# 2.87e-21
C855 a_12030_3213# a_12146_3239# 0.0397f
C856 x4.X a_7953_3239# 0.00272f
C857 a_8383_2340# a_9709_2550# 4.7e-22
C858 a_8696_2366# a_9441_2340# 0.199f
C859 a_8938_2340# a_9237_2340# 0.0334f
C860 x4.X a_4925_2550# 0.00127f
C861 a_11543_3213# a_12264_3521# 0.00185f
C862 a_11195_4112# a_11075_3605# 1.12e-20
C863 x27.Q_N a_6845_2340# 6.49e-21
C864 x4.X a_4585_3239# 5e-19
C865 a_4074_4775# a_4368_4775# 0.199f
C866 a_3619_4801# a_4855_4775# 0.0265f
C867 a_3453_4801# a_4681_4801# 0.0334f
C868 a_10776_4086# a_11630_4086# 0.0492f
C869 a_11089_4112# a_11629_4386# 0.139f
C870 x45.Q_N x75.Q_N 6.77e-21
C871 x5.X a_8684_5167# 0.00465f
C872 x20.Q_N a_4368_4775# 3e-20
C873 x30.Q_N a_6845_4386# 0.0327f
C874 a_6606_4801# x45.Q_N 2.3e-19
C875 a_2060_2640# a_2198_2732# 1.09e-19
C876 a_1520_2366# a_2479_2648# 1.21e-20
C877 a_1762_2340# a_1626_2366# 0.0282f
C878 a_2853_5648# a_3258_5648# 0.0197f
C879 x5.X check[0] 0.789f
C880 sel_bit[0] x48.Q 0.0566f
C881 a_2853_5648# sel_bit[1] 0.0368f
C882 a_7073_4801# a_8237_4801# 6.38e-20
C883 a_7247_4775# a_8403_4801# 2.64e-19
C884 check[0] a_4854_3213# 0.00313f
C885 D[3] a_11088_2366# 8.67e-19
C886 a_12146_3239# a_11628_2640# 5.05e-21
C887 x4.X a_11075_3605# 0.0178f
C888 a_10795_4801# a_12031_4775# 0.0264f
C889 a_11250_4775# a_11544_4775# 0.199f
C890 a_10629_4801# a_11857_4801# 0.0334f
C891 a_2883_5674# a_1511_4112# 1.46e-20
C892 a_8803_4112# a_8402_3239# 4.04e-21
C893 VDD a_9152_4775# 0.449f
C894 comparator_out a_11856_3239# 1.89e-19
C895 a_4454_4086# a_4591_4478# 0.00907f
C896 a_11195_4112# a_11088_2366# 8.38e-21
C897 x36.Q_N a_10155_2366# 1.34e-20
C898 x36.Q_N a_11965_3239# 1.68e-19
C899 a_9639_4775# a_8697_4112# 0.00161f
C900 a_8403_4801# a_9442_4086# 0.00221f
C901 a_8858_4775# a_9238_4086# 0.00336f
C902 a_9152_4775# a_8939_4086# 3.72e-19
C903 check[4] comparator_out 0.0222f
C904 a_3504_2340# a_4452_2640# 9.65e-21
C905 a_11194_2366# a_11564_2366# 4.11e-20
C906 a_6010_3239# a_7158_3605# 2.13e-19
C907 a_6465_3213# a_6930_3521# 9.46e-19
C908 a_3258_5648# a_3671_5674# 3.58e-19
C909 x4.X a_11088_2366# 0.112f
C910 x4.X a_5170_4478# 9.15e-19
C911 check[6] a_4018_2366# 1.17e-19
C912 comparator_out a_11629_2340# 0.183f
C913 a_4367_3213# a_4452_2640# 5.32e-19
C914 a_4680_3239# a_3912_2366# 2.17e-19
C915 a_3806_3239# a_3599_2340# 2.02e-19
C916 a_5897_4086# x45.Q_N 0.182f
C917 a_5992_4086# a_6845_4386# 0.0264f
C918 a_6305_4112# a_6547_4086# 0.124f
C919 x5.X a_6376_5167# 4.16e-19
C920 VDD a_4452_2640# 0.273f
C921 a_4971_4801# a_4367_3213# 1.05e-20
C922 a_6292_5167# a_6376_5167# 0.00972f
C923 a_5845_4801# a_6710_5083# 0.00276f
C924 a_6760_4775# a_6199_4801# 8.23e-22
C925 a_3899_3605# a_4213_3239# 0.0258f
C926 a_3806_3239# a_3983_3605# 8.94e-19
C927 a_4367_3213# a_4766_3605# 0.00133f
C928 a_7247_4775# a_7073_4801# 0.197f
C929 a_3618_3239# a_4585_3239# 0.00126f
C930 a_3452_3239# a_5088_3521# 1.25e-19
C931 D[0] a_9638_3213# 1.68e-20
C932 a_7072_3239# a_7317_2550# 1.85e-20
C933 a_9639_4775# a_11857_4801# 1.86e-21
C934 VDD a_4766_3605# 0.00394f
C935 VDD a_4971_4801# 0.0111f
C936 x30.Q_N a_8236_3239# 8.92e-20
C937 x39.Q_N a_11942_3605# 3.64e-19
C938 x30.Q_N a_6977_3239# 4.04e-19
C939 VDD a_7561_2732# 0.0042f
C940 VDD a_10628_3239# 0.791f
C941 a_11629_4386# a_11767_4478# 1.09e-19
C942 a_11089_4112# a_12048_4394# 1.21e-20
C943 a_11331_4086# a_11195_4112# 0.0282f
C944 x27.D a_4539_5083# 3.01e-21
C945 check[2] a_10346_4801# 0.0147f
C946 eob a_2993_5674# 9.62e-20
C947 VDD a_9369_3239# 6.2e-19
C948 a_9638_3213# a_11543_3213# 3.71e-20
C949 a_6844_2640# x57.Q_N 4.82e-21
C950 a_6845_2340# a_7317_2550# 0.15f
C951 check[2] a_11628_2640# 3.14e-19
C952 check[2] a_2784_5996# 6.63e-19
C953 a_2389_5648# a_2883_5674# 0.169f
C954 x5.X a_4389_4478# 4.04e-20
C955 x42.Q_N a_9101_3521# 0.00136f
C956 check[2] a_5897_4086# 1.35e-21
C957 x4.X a_11331_4086# 0.00706f
C958 x30.Q_N a_6984_2366# 0.00473f
C959 a_4019_4112# a_3899_3605# 1.12e-20
C960 a_9442_4086# a_9710_4296# 0.205f
C961 a_9238_4086# x42.Q_N 0.00114f
C962 a_11834_4086# comparator_out 4.39e-21
C963 VDD a_9376_2366# 6.2e-19
C964 a_4214_4801# a_4367_3213# 1.61e-20
C965 x27.Q_N a_3452_3239# 2.63e-19
C966 a_4681_4801# a_4790_4801# 0.00707f
C967 VDD a_4591_4478# 0.0172f
C968 x5.X a_11943_5167# 1.78e-19
C969 D[4] a_9441_2340# 6.5e-20
C970 a_10628_3239# D[2] 6.24e-20
C971 a_10794_3239# a_12737_3239# 6.86e-21
C972 D[1] a_12146_3239# 1.57e-20
C973 D[1] a_11761_3239# 5.48e-20
C974 x4.X a_6198_3239# 0.00604f
C975 a_8237_4801# a_9370_4801# 2.56e-19
C976 a_8858_4775# a_8998_4801# 0.07f
C977 a_9152_4775# a_9323_5083# 0.00652f
C978 a_8403_4801# a_8792_4801# 0.0019f
C979 VDD a_4214_4801# 0.035f
C980 x45.Q_N a_4970_3239# 9.58e-21
C981 a_5844_3239# a_6709_3521# 0.00276f
C982 x48.Q a_2788_5674# 1.65e-19
C983 a_6305_4112# a_6411_4112# 0.051f
C984 a_6547_4086# a_6983_4478# 0.00412f
C985 a_6845_4386# a_6781_4478# 2.13e-19
C986 a_6846_4086# a_6505_4394# 1.25e-19
C987 VDD a_11390_4801# 0.0332f
C988 a_2289_4801# a_1511_4112# 0.00374f
C989 check[4] a_8696_2366# 1.1e-20
C990 a_11857_4801# a_10794_3239# 6.75e-21
C991 a_5561_3239# a_5844_3239# 8.18e-19
C992 eob a_1762_2340# 2.19e-19
C993 a_1207_2340# a_1520_2366# 0.273f
C994 a_6011_4801# check[5] 1.26e-20
C995 a_9709_2550# a_9577_2366# 0.0258f
C996 a_9237_2340# a_11088_2366# 3.08e-19
C997 a_9236_2640# a_11330_2340# 4.16e-20
C998 x4.X a_7049_2340# 0.00149f
C999 check[1] a_4658_4086# 4.01e-21
C1000 x5.A a_2853_5648# 2.03e-20
C1001 check[4] a_10795_4801# 0.164f
C1002 x4.A a_1762_2340# 3.45e-19
C1003 VDD a_7954_4801# 0.193f
C1004 a_1227_4801# a_2463_4775# 0.0267f
C1005 a_1682_4775# a_1976_4775# 0.198f
C1006 x4.X a_1508_5167# 0.138f
C1007 a_1061_4801# a_2289_4801# 0.0334f
C1008 a_3505_4086# a_4453_4386# 8.38e-21
C1009 a_1511_4112# a_4454_4086# 7.27e-20
C1010 a_3600_4086# a_4155_4086# 0.197f
C1011 check[0] a_5896_2340# 0.028f
C1012 check[2] a_11630_4086# 1.95e-19
C1013 x36.Q_N a_9236_2640# 0.00112f
C1014 a_3900_5167# x27.Q_N 8.65e-20
C1015 a_4368_4775# a_5089_5083# 0.00185f
C1016 D[6] a_2200_2366# 1.47e-19
C1017 a_2061_2340# a_4112_2648# 4.06e-20
C1018 x5.X x33.Q_N 0.00113f
C1019 a_11628_2640# a_12047_2648# 2.46e-19
C1020 a_11088_2366# a_12547_2366# 4.94e-21
C1021 a_11833_2340# a_11766_2732# 9.46e-19
C1022 a_10775_2340# a_11564_2366# 4.2e-20
C1023 x63.Q_N a_11288_2648# 2.02e-20
C1024 x4.X D[3] 5.34e-19
C1025 x4.X a_1112_2340# 0.0104f
C1026 check[0] x30.Q_N 0.00106f
C1027 VDD a_9578_4112# 0.0326f
C1028 x4.X x66.Q_N 0.00462f
C1029 x4.X a_3913_4112# 0.112f
C1030 check[6] a_3599_2340# 2.38e-20
C1031 a_11544_4775# a_12265_5083# 0.00185f
C1032 a_11076_5167# x36.Q_N 1.74e-20
C1033 a_4854_3213# a_6291_3605# 7.98e-21
C1034 a_4367_3213# a_6759_3213# 3.6e-20
C1035 a_6466_4775# a_6759_3213# 7.57e-21
C1036 a_5845_4801# a_7072_3239# 4.76e-21
C1037 x4.X a_11195_4112# 0.00334f
C1038 a_4453_4386# x45.Q_N 2.05e-19
C1039 a_4454_4086# comparator_out 3.22e-20
C1040 a_8939_4086# a_9578_4112# 0.00316f
C1041 a_9710_4296# a_10156_4112# 0.0367f
C1042 a_9237_4386# a_9377_4112# 0.00126f
C1043 a_12548_4112# comparator_out 4.04e-20
C1044 VDD a_6759_3213# 0.353f
C1045 check[6] a_7073_4801# 4.06e-20
C1046 a_3912_2366# a_4388_2366# 2.87e-21
C1047 x33.Q_N a_9237_4386# 0.0344f
C1048 a_8998_4801# x42.Q_N 2.35e-19
C1049 a_6759_3213# a_7362_3239# 0.0552f
C1050 a_9465_4801# check[4] 1.08e-19
C1051 check[2] D[1] 0.171f
C1052 eob a_1822_4801# 0.00828f
C1053 a_2853_5648# x27.D 3.86e-19
C1054 a_5561_3239# D[5] 0.00127f
C1055 a_2389_5648# a_2289_4801# 0.0019f
C1056 check[0] a_3373_5674# 0.0228f
C1057 check[2] a_2463_4775# 7.62e-20
C1058 a_1822_4801# x4.A 2.88e-19
C1059 VDD a_6546_2340# 0.177f
C1060 check[0] a_5992_4086# 0.0142f
C1061 a_5991_2340# a_6504_2648# 0.00945f
C1062 a_9638_3213# a_10345_3239# 0.0968f
C1063 a_9151_3213# D[1] 4.66e-19
C1064 D[7] x51.Q_N 0.00276f
C1065 a_12031_4775# a_11089_4112# 0.00161f
C1066 a_10795_4801# a_11834_4086# 0.00221f
C1067 a_11250_4775# a_11630_4086# 0.00336f
C1068 a_11544_4775# a_11331_4086# 3.72e-19
C1069 check[1] x5.X 0.767f
C1070 check[1] a_6292_5167# 1.94e-19
C1071 eob a_621_4112# 9.98e-19
C1072 check[2] a_4453_4386# 1.41e-20
C1073 a_1062_5674# a_1338_5674# 0.00104f
C1074 a_3913_4112# a_3618_3239# 4.9e-19
C1075 a_3600_4086# a_4073_3213# 2.45e-19
C1076 VDD a_9655_2648# 0.00984f
C1077 a_4318_5083# check[6] 1.19e-21
C1078 x3.A a_897_4112# 0.3f
C1079 a_621_4112# x4.A 6.66e-19
C1080 reset a_1511_4112# 1.58e-19
C1081 a_11249_3213# a_11856_3239# 0.00187f
C1082 a_10628_3239# a_11159_3605# 0.0018f
C1083 a_10794_3239# a_10982_3239# 0.163f
C1084 a_11075_3605# a_12030_3213# 4.7e-22
C1085 VDD a_1511_4112# 1.55f
C1086 check[5] a_9102_5083# 8.63e-22
C1087 a_8997_3239# a_9573_3239# 2.46e-21
C1088 VDD a_11289_4394# 0.00506f
C1089 check[1] a_9237_4386# 1.6e-19
C1090 comparator_out a_3504_2340# 0.00285f
C1091 a_11494_5083# check[3] 2.79e-19
C1092 x77.Y a_4018_2366# 6.03e-20
C1093 x42.Q_N a_9573_3239# 7.87e-19
C1094 x4.X a_3618_3239# 0.0489f
C1095 x27.Q_N x54.Q_N 4.08e-19
C1096 x5.X a_7050_4086# 9.61e-19
C1097 x30.Q_N a_9172_2366# 1.14e-20
C1098 x5.X a_5844_3239# 8.91e-20
C1099 a_7247_4775# a_6845_4386# 6.17e-19
C1100 a_6760_4775# a_6846_4086# 4.63e-19
C1101 a_6011_4801# x45.Q_N 7.77e-20
C1102 a_9237_4386# a_9954_4112# 0.0019f
C1103 check[4] x69.Q_N 0.00316f
C1104 a_2289_4801# a_3619_4801# 5.38e-20
C1105 a_4367_3213# comparator_out 5.5e-19
C1106 a_4854_3213# a_5844_3239# 0.00116f
C1107 a_6292_5167# a_5844_3239# 8.3e-21
C1108 x48.Q x77.Y 6.96e-20
C1109 a_2463_4775# x20.Q_N 0.129f
C1110 VDD a_1061_4801# 0.901f
C1111 a_9441_2340# a_10155_2366# 6.99e-20
C1112 a_9709_2550# a_9953_2732# 0.00972f
C1113 a_9237_2340# D[3] 0.336f
C1114 reset comparator_out 2.03e-20
C1115 a_12030_3213# a_11088_2366# 8.4e-19
C1116 a_10794_3239# a_11833_2340# 0.00154f
C1117 a_11249_3213# a_11629_2340# 0.00199f
C1118 a_11543_3213# a_11330_2340# 2.17e-19
C1119 VDD a_7318_4296# 0.317f
C1120 x4.X a_9464_3239# 0.00475f
C1121 VDD comparator_out 1.51f
C1122 x4.X a_7186_4112# 0.00311f
C1123 a_8237_4801# a_8236_3239# 6.9e-19
C1124 a_6846_4086# a_9238_4086# 1.37e-19
C1125 a_6305_4112# x42.Q_N 5.52e-21
C1126 check[4] a_10775_2340# 7.18e-21
C1127 a_4074_4775# a_4453_4386# 3.92e-19
C1128 a_3453_4801# a_4658_4086# 6.96e-19
C1129 a_3619_4801# a_4454_4086# 1.18e-19
C1130 a_4368_4775# a_3913_4112# 5.67e-20
C1131 a_3900_5167# a_4155_4086# 2.46e-20
C1132 x20.Q_N a_4453_4386# 1.28e-19
C1133 x36.Q_N a_11543_3213# 0.00494f
C1134 a_2777_2732# a_2979_2366# 8.94e-19
C1135 a_1762_2340# a_2401_2366# 0.00316f
C1136 a_2060_2640# a_2200_2366# 0.00126f
C1137 a_1520_2366# a_3599_2340# 8.34e-21
C1138 a_11088_2366# a_11628_2640# 0.139f
C1139 a_10775_2340# a_11629_2340# 0.0492f
C1140 a_6978_4801# check[5] 1.84e-20
C1141 x4.X a_9237_2340# 0.00274f
C1142 check[4] a_11762_4801# 5.42e-20
C1143 comparator_out D[2] 0.0211f
C1144 check[6] a_6010_3239# 9.27e-20
C1145 comparator_out x60.Q_N 3.61e-19
C1146 x4.X a_4368_4775# 0.101f
C1147 a_1061_4801# a_3807_4801# 3.65e-21
C1148 a_1338_5674# x5.X 0.17f
C1149 x27.Q_N a_5372_4112# 0.0147f
C1150 check[2] a_6011_4801# 1.18e-19
C1151 x4.X a_11544_4775# 0.105f
C1152 x36.Q_N a_11330_2340# 0.16f
C1153 VDD a_2265_2340# 0.326f
C1154 a_3452_3239# a_4073_3213# 0.115f
C1155 D[6] a_4388_2366# 1.34e-19
C1156 a_3912_2366# a_4018_2366# 0.0552f
C1157 a_4154_2340# a_4590_2732# 0.00412f
C1158 a_4452_2640# a_4388_2732# 2.13e-19
C1159 a_4453_2340# a_4112_2648# 1.25e-19
C1160 a_10983_4801# comparator_out 1.78e-20
C1161 x4.X a_12547_2366# 5.99e-20
C1162 VDD a_2389_5648# 0.696f
C1163 a_4970_3239# a_4925_2550# 1.01e-20
C1164 x30.Q_N x33.Q_N 2.51e-20
C1165 check[1] a_9656_4394# 1.56e-20
C1166 x5.X D[5] 3.43e-19
C1167 check[6] a_4793_2366# 4.42e-19
C1168 a_5561_3239# a_4453_2340# 4.83e-19
C1169 a_11089_4112# a_11856_3239# 2.16e-19
C1170 a_11629_4386# a_11543_3213# 5.72e-19
C1171 a_10776_4086# a_10982_3239# 2.44e-19
C1172 x39.Q_N a_10628_3239# 0.0434f
C1173 x30.Q_N a_6291_3605# 0.00193f
C1174 check[2] a_8697_4112# 0.00313f
C1175 x5.X a_7764_4112# 9.62e-19
C1176 x33.Q_N a_9754_3239# 0.00342f
C1177 a_3170_4801# a_3453_4801# 8.18e-19
C1178 VDD a_8683_3605# 0.176f
C1179 a_5896_2340# a_6304_2366# 6.04e-19
C1180 a_4592_2366# a_4793_2366# 3.34e-19
C1181 a_8402_3239# a_9101_3521# 2.46e-19
C1182 a_8236_3239# a_9322_3521# 0.00907f
C1183 VDD a_8289_4086# 0.189f
C1184 a_8939_4086# a_8683_3605# 1.7e-20
C1185 a_9237_4386# a_8857_3213# 0.0015f
C1186 a_8697_4112# a_9151_3213# 3.33e-20
C1187 a_9442_4086# a_8236_3239# 0.00195f
C1188 a_9238_4086# a_8402_3239# 6.04e-20
C1189 x4.X a_8897_4394# 1.75e-19
C1190 a_11089_4112# a_11629_2340# 1.4e-21
C1191 a_11331_4086# a_11628_2640# 4.75e-21
C1192 x30.Q_N a_6304_2366# 0.0928f
C1193 check[2] a_4681_4801# 4.32e-20
C1194 x5.X a_3453_4801# 0.255f
C1195 x4.X a_7363_4801# 0.00557f
C1196 x33.Q_N x63.Q_N 7.78e-20
C1197 a_3619_4801# a_4367_3213# 2.05e-21
C1198 a_4074_4775# a_3899_3605# 1.33e-23
C1199 a_3900_5167# a_4073_3213# 3.52e-21
C1200 VDD a_8696_2366# 0.348f
C1201 x20.Q_N a_3899_3605# 2.96e-20
C1202 x5.X a_10629_4801# 0.27f
C1203 a_10345_3239# a_11543_3213# 5.62e-20
C1204 D[1] a_11075_3605# 2.08e-19
C1205 a_9638_3213# a_9441_2340# 2.52e-19
C1206 a_9151_3213# a_9709_2550# 1.62e-19
C1207 a_8403_4801# a_8858_4775# 0.153f
C1208 a_8237_4801# a_8684_5167# 0.15f
C1209 x36.Q_N a_11629_4386# 0.0351f
C1210 VDD a_3619_4801# 0.617f
C1211 a_11390_4801# x39.Q_N 2.02e-19
C1212 check[2] a_11768_2366# 3.3e-19
C1213 a_6547_4086# a_6010_3239# 1.07e-20
C1214 a_6305_4112# a_6465_3213# 0.00148f
C1215 VDD a_2697_5083# 0.00615f
C1216 a_4926_4296# a_4452_2640# 6.02e-22
C1217 a_4453_4386# a_4925_2550# 6.45e-21
C1218 check[1] x30.Q_N 0.0373f
C1219 x77.Y a_3599_2340# 2.75e-19
C1220 VDD a_10795_4801# 0.593f
C1221 x30.Q_N a_8802_2366# 9.32e-20
C1222 x48.Q a_4113_4394# 5.88e-19
C1223 a_1227_4801# a_897_4112# 4.21e-19
C1224 a_4971_4801# a_4926_4296# 1.9e-20
C1225 x48.Q a_4539_5083# 6.59e-19
C1226 VDD a_11194_2366# 4.84e-19
C1227 D[1] a_11088_2366# 3.91e-20
C1228 a_9236_2640# a_9441_2340# 0.153f
C1229 a_8696_2366# x60.Q_N 0.00553f
C1230 a_11856_3239# a_11965_3239# 0.00707f
C1231 a_12030_3213# x66.Q_N 0.124f
C1232 a_6305_4112# a_5991_2340# 5.05e-21
C1233 a_5844_3239# a_5896_2340# 4.5e-19
C1234 check[4] a_10155_2366# 0.00335f
C1235 check[2] a_9375_4478# 1.05e-20
C1236 x4.X a_6606_4801# 7.25e-19
C1237 x4.X x75.Q_N 0.00464f
C1238 a_3453_4801# a_3984_5167# 0.0018f
C1239 a_3619_4801# a_3807_4801# 0.162f
C1240 a_3900_5167# a_4855_4775# 4.7e-22
C1241 a_4074_4775# a_4681_4801# 0.00187f
C1242 a_2853_5648# a_3876_6040# 0.00747f
C1243 check[2] a_9102_5083# 1.52e-19
C1244 a_1822_4801# a_2398_4801# 2.46e-21
C1245 a_11331_4086# a_11630_4086# 0.0334f
C1246 a_11089_4112# a_11834_4086# 0.199f
C1247 a_10776_4086# a_12102_4296# 4.7e-22
C1248 x5.X a_9639_4775# 0.00985f
C1249 check[1] a_3373_5674# 0.027f
C1250 x20.Q_N a_4681_4801# 2.69e-20
C1251 a_9578_4112# x39.Q_N 5.6e-20
C1252 a_1207_2340# D[6] 3.57e-20
C1253 a_2060_2640# a_2479_2648# 2.46e-19
C1254 a_1520_2366# a_2979_2366# 6.59e-21
C1255 a_2265_2340# a_2198_2732# 9.46e-19
C1256 x51.Q_N a_1720_2648# 2.02e-20
C1257 x30.Q_N a_5844_3239# 2.88e-19
C1258 a_7247_4775# a_8684_5167# 7.98e-21
C1259 a_10155_2366# a_11629_2340# 3.65e-21
C1260 D[3] a_11628_2640# 4.01e-20
C1261 a_12146_3239# a_11833_2340# 3.49e-20
C1262 x4.X a_12030_3213# 0.116f
C1263 check[1] a_5992_4086# 5.87e-20
C1264 a_3258_5648# a_1511_4112# 3.06e-19
C1265 a_11076_5167# a_12031_4775# 4.7e-22
C1266 a_10795_4801# a_10983_4801# 0.162f
C1267 a_11250_4775# a_11857_4801# 0.00187f
C1268 a_10629_4801# a_11160_5167# 0.0018f
C1269 sel_bit[1] a_1511_4112# 3.24e-20
C1270 a_8803_4112# a_8683_3605# 1.12e-20
C1271 VDD a_9465_4801# 0.343f
C1272 a_3600_4086# a_4389_4112# 4.2e-20
C1273 a_4454_4086# a_4872_4394# 0.00276f
C1274 a_4453_4386# a_5170_4478# 4.45e-20
C1275 x4.X a_10346_4801# 0.0067f
C1276 x27.Q_N a_4155_4086# 1.3e-22
C1277 clk_sar a_897_4112# 1.96e-20
C1278 D[6] a_4018_2366# 0.0021f
C1279 a_9152_4775# a_9238_4086# 4.63e-19
C1280 a_9639_4775# a_9237_4386# 6.17e-19
C1281 a_8403_4801# x42.Q_N 7.79e-20
C1282 a_3599_2340# a_3912_2366# 0.273f
C1283 a_3373_5674# a_3877_5674# 5.33e-19
C1284 a_6010_3239# a_6399_3239# 0.0019f
C1285 a_6759_3213# a_6930_3521# 0.00652f
C1286 a_6465_3213# a_6605_3239# 0.07f
C1287 sel_bit[1] a_1061_4801# 7.54e-20
C1288 x4.X a_11628_2640# 0.00712f
C1289 a_6411_4112# a_6010_3239# 4.04e-21
C1290 x4.X a_5897_4086# 0.00454f
C1291 x5.X a_4453_2340# 2.59e-20
C1292 a_8803_4112# a_8696_2366# 8.38e-21
C1293 comparator_out a_12101_2550# 0.00818f
C1294 x75.Q a_6759_3213# 9.18e-20
C1295 a_4854_3213# a_4453_2340# 8.72e-19
C1296 a_4367_3213# a_4657_2340# 0.00144f
C1297 a_4680_3239# a_4452_2640# 1.11e-20
C1298 a_4593_4112# x45.Q_N 3.1e-20
C1299 a_6305_4112# a_6846_4086# 0.125f
C1300 a_6547_4086# a_6845_4386# 0.137f
C1301 a_5992_4086# a_5844_3239# 8.29e-19
C1302 check[1] eob 0.00405f
C1303 VDD a_4657_2340# 0.307f
C1304 D[5] a_5896_2340# 0.0999f
C1305 a_3618_3239# x75.Q_N 1.93e-21
C1306 a_6466_4775# a_6710_5083# 0.0104f
C1307 a_6011_4801# a_6931_5083# 1.09e-19
C1308 a_4680_3239# a_4766_3605# 0.00976f
C1309 D[0] a_8590_3239# 5.04e-19
C1310 a_6605_3239# a_5991_2340# 4.6e-20
C1311 a_9152_4775# a_9755_4801# 0.0552f
C1312 sel_bit[0] a_621_4112# 8.01e-21
C1313 VDD a_6710_5083# 0.00984f
C1314 check[2] a_10982_3239# 0.00707f
C1315 x20.Q_N a_1996_2732# 3.64e-19
C1316 VDD a_4007_3239# 2.82e-19
C1317 x30.Q_N D[5] 0.00272f
C1318 x30.Q_N x72.Q_N 0.0201f
C1319 a_12147_4801# a_11543_3213# 1.05e-20
C1320 VDD D[4] 0.221f
C1321 VDD a_11249_3213# 0.308f
C1322 a_11629_4386# a_12048_4394# 2.46e-19
C1323 a_11834_4086# a_11767_4478# 9.46e-19
C1324 a_10776_4086# a_11565_4112# 4.2e-20
C1325 x39.Q_N a_11289_4394# 2.02e-20
C1326 x30.Q_N a_7764_4112# 0.0147f
C1327 VDD x69.Q_N 0.0716f
C1328 a_9638_3213# a_11856_3239# 1.86e-21
C1329 a_9151_3213# a_10982_3239# 3.42e-20
C1330 a_2853_5648# x48.Q 0.016f
C1331 a_2389_5648# a_3258_5648# 0.0296f
C1332 sel_bit[0] check[0] 0.163f
C1333 check[2] a_11833_2340# 4.61e-19
C1334 a_2389_5648# sel_bit[1] 0.0628f
C1335 x77.Y a_6010_3239# 0.00188f
C1336 x42.Q_N a_9550_3605# 3.64e-19
C1337 x4.X a_11630_4086# 0.0441f
C1338 x30.Q_N a_8383_2340# 1.64e-19
C1339 check[4] a_9638_3213# 0.00527f
C1340 a_9710_4296# x42.Q_N 0.00244f
C1341 x39.Q_N comparator_out 6.03e-19
C1342 VDD a_10775_2340# 0.561f
C1343 x27.Q_N a_4073_3213# 4.88e-19
C1344 x27.Q_N a_5845_4801# 4.37e-19
C1345 D[1] D[3] 0.345f
C1346 x5.X a_11184_4801# 2.88e-19
C1347 VDD a_4872_4394# 0.0102f
C1348 D[4] x60.Q_N 0.00109f
C1349 a_11249_3213# D[2] 1.23e-20
C1350 x4.X a_4970_3239# 5.69e-19
C1351 a_9639_4775# a_9551_5167# 7.71e-20
C1352 a_8858_4775# a_9370_4801# 9.75e-19
C1353 a_9465_4801# a_9323_5083# 0.00412f
C1354 a_8684_5167# a_8792_4801# 0.00812f
C1355 a_9152_4775# a_8998_4801# 0.00943f
C1356 a_8237_4801# x33.Q_N 1.26e-19
C1357 VDD a_4586_4801# 0.00495f
C1358 comparator_out a_4388_2732# 1.8e-19
C1359 x45.Q_N a_6709_3521# 0.00136f
C1360 x48.Q a_3671_5674# 0.0017f
C1361 x77.Y a_4793_2366# 5.33e-22
C1362 x36.Q_N a_12147_4801# 3.8e-19
C1363 x45.Q_N a_5170_4112# 3.4e-20
C1364 a_6846_4086# a_6983_4478# 0.00907f
C1365 VDD a_11762_4801# 0.00445f
C1366 check[4] a_9236_2640# 0.0285f
C1367 a_12031_4775# a_11543_3213# 1.08e-22
C1368 a_11544_4775# a_12030_3213# 1.06e-20
C1369 x45.Q_N a_5561_3239# 1.19e-20
C1370 x5.X check[5] 0.17f
C1371 x75.Q comparator_out 0.00133f
C1372 eob a_2061_2340# 0.00216f
C1373 a_1520_2366# a_1762_2340# 0.124f
C1374 a_1207_2340# a_2060_2640# 0.0264f
C1375 check[0] check[6] 0.45f
C1376 a_6760_4775# a_7954_4801# 6.04e-19
C1377 a_6292_5167# check[5] 7.62e-21
C1378 a_1338_5674# eob 5.41e-19
C1379 a_12030_3213# a_12547_2366# 2.38e-19
C1380 x4.X D[1] 0.0011f
C1381 a_9236_2640# a_11629_2340# 2.9e-21
C1382 a_9237_2340# a_11628_2640# 4e-20
C1383 a_9709_2550# a_11088_2366# 5.19e-21
C1384 x4.X x57.Q_N 0.00786f
C1385 check[4] a_11076_5167# 0.0011f
C1386 a_3373_5674# a_3453_4801# 1.45e-21
C1387 x4.X a_2463_4775# 0.148f
C1388 a_1227_4801# a_1415_4801# 0.163f
C1389 a_1682_4775# a_2289_4801# 0.00187f
C1390 a_1061_4801# a_1592_5167# 0.0018f
C1391 a_2969_6040# x20.Q_N 1.2e-20
C1392 a_1338_5674# x4.A 2.32e-21
C1393 a_3913_4112# a_4453_4386# 0.139f
C1394 a_3600_4086# a_4454_4086# 0.0492f
C1395 a_4855_4775# a_5372_4112# 4.23e-19
C1396 x5.X a_10776_4086# 0.0184f
C1397 check[2] a_12102_4296# 4.54e-20
C1398 a_4855_4775# x27.Q_N 0.128f
C1399 a_2060_2640# a_4018_2366# 2.19e-20
C1400 a_2979_2366# a_3912_2366# 3.42e-20
C1401 D[6] a_3599_2340# 0.0144f
C1402 a_11629_2340# a_12345_2732# 0.0018f
C1403 a_11088_2366# a_11768_2366# 3.73e-19
C1404 a_11833_2340# a_12047_2648# 0.0104f
C1405 a_11330_2340# a_11564_2366# 0.00707f
C1406 a_11628_2640# a_12547_2366# 0.159f
C1407 a_12147_4801# a_11629_4386# 8.84e-21
C1408 VDD a_11089_4112# 0.448f
C1409 check[1] a_8237_4801# 0.00245f
C1410 x4.X a_4453_4386# 0.0483f
C1411 a_12031_4775# x36.Q_N 0.126f
C1412 check[6] a_4154_2340# 1.2e-19
C1413 a_6760_4775# a_6759_3213# 0.00121f
C1414 x4.X a_12346_4478# 9.15e-19
C1415 a_4658_4086# x45.Q_N 3.93e-20
C1416 a_9237_4386# a_10776_4086# 1.52e-19
C1417 a_9442_4086# a_9377_4112# 9.75e-19
C1418 a_9238_4086# a_9578_4112# 6.04e-20
C1419 x42.Q_N a_10681_4086# 1.37e-20
C1420 x36.Q_N a_11564_2366# 9.42e-19
C1421 VDD a_7072_3239# 0.18f
C1422 a_4154_2340# a_4592_2366# 0.00276f
C1423 a_3912_2366# a_4793_2366# 0.00943f
C1424 a_4453_2340# a_5896_2340# 8.18e-19
C1425 a_7072_3239# a_7362_3239# 0.0282f
C1426 a_7246_3213# a_7181_3239# 4.2e-20
C1427 eob a_3453_4801# 5.9e-20
C1428 eob a_2194_4801# 0.00151f
C1429 a_10681_4086# a_10680_2340# 1.07e-20
C1430 x30.Q_N a_4453_2340# 1.57e-19
C1431 check[0] a_6547_4086# 3.86e-19
C1432 VDD a_6845_2340# 0.784f
C1433 a_6304_2366# a_6780_2732# 0.00133f
C1434 a_9464_3239# D[1] 5.18e-20
C1435 a_10795_4801# x39.Q_N 7.79e-20
C1436 a_12031_4775# a_11629_4386# 6.17e-19
C1437 a_11544_4775# a_11630_4086# 4.63e-19
C1438 a_3600_4086# a_3504_2340# 2.97e-20
C1439 check[1] a_7247_4775# 0.0127f
C1440 x33.Q_N a_9574_4801# 7.27e-21
C1441 a_1227_4801# a_3170_4801# 1.76e-19
C1442 x39.Q_N a_11194_2366# 5e-20
C1443 a_1061_4801# x27.D 5.94e-20
C1444 x5.A a_2389_5648# 6.17e-20
C1445 x5.X a_3505_4086# 0.00259f
C1446 check[2] a_4658_4086# 4.4e-21
C1447 a_1062_5674# check[2] 1.82e-20
C1448 x30.Q_N a_7763_2366# 0.0318f
C1449 clk_sar a_1062_5674# 0.185f
C1450 x5.X a_11565_4478# 1.76e-19
C1451 a_4454_4086# a_3452_3239# 6.54e-20
C1452 a_4453_4386# a_3618_3239# 4.11e-20
C1453 a_3600_4086# a_4367_3213# 8.83e-19
C1454 a_4155_4086# a_4073_3213# 1.02e-19
C1455 a_3913_4112# a_3899_3605# 1.61e-19
C1456 VDD a_10155_2366# 0.109f
C1457 VDD a_12264_3521# 0.00506f
C1458 VDD a_3600_4086# 0.741f
C1459 D[1] a_9237_2340# 0.0263f
C1460 a_6845_2340# x60.Q_N 2.94e-19
C1461 a_11543_3213# a_11856_3239# 0.124f
C1462 a_11075_3605# a_10982_3239# 0.0367f
C1463 a_11249_3213# a_11159_3605# 6.69e-20
C1464 a_10794_3239# a_9754_3239# 9.75e-21
C1465 VDD a_11767_4478# 0.0163f
C1466 check[1] a_9442_4086# 1.18e-19
C1467 x5.X a_1227_4801# 0.0165f
C1468 a_11943_5167# check[3] 4.39e-19
C1469 x4.X a_6011_4801# 0.00494f
C1470 x5.X x45.Q_N 0.00731f
C1471 x4.X a_3899_3605# 0.018f
C1472 check[4] a_11543_3213# 8.39e-21
C1473 x4.X a_11966_4801# 2.39e-19
C1474 x45.Q_N a_4854_3213# 1.37e-20
C1475 a_6760_4775# a_7318_4296# 2.85e-19
C1476 a_6292_5167# x45.Q_N 9.97e-20
C1477 a_7247_4775# a_7050_4086# 4.44e-19
C1478 a_4680_3239# comparator_out 1.77e-19
C1479 a_1415_4801# x20.Q_N 5.43e-21
C1480 VDD a_1682_4775# 0.337f
C1481 x27.Q_N a_6400_4801# 2.58e-20
C1482 x33.Q_N a_10156_4112# 0.0147f
C1483 D[2] a_11965_3239# 9.32e-21
C1484 a_12030_3213# a_11628_2640# 3.43e-19
C1485 a_11543_3213# a_11629_2340# 2.19e-19
C1486 x66.Q_N a_12737_3239# 0.178f
C1487 x4.X a_8767_3605# 9.07e-19
C1488 comparator_out a_6504_2648# 1.52e-19
C1489 x45.Q_N a_7181_3239# 7.87e-19
C1490 x4.X a_8697_4112# 0.109f
C1491 a_8403_4801# a_8402_3239# 1.39e-19
C1492 a_4368_4775# a_4453_4386# 7.46e-19
C1493 a_3807_4801# a_3600_4086# 3.44e-19
C1494 a_4681_4801# a_3913_4112# 3.76e-19
C1495 check[2] a_3170_4801# 1.57e-20
C1496 a_2579_4801# a_1511_4112# 3.99e-19
C1497 a_6845_4386# x42.Q_N 1.95e-19
C1498 x20.Q_N a_4658_4086# 2.19e-20
C1499 a_9238_4086# comparator_out 3.21e-20
C1500 check[0] a_6411_4112# 4.09e-19
C1501 x36.Q_N a_11856_3239# 0.00293f
C1502 a_2979_2366# D[6] 6.09e-19
C1503 D[3] a_11768_2366# 7.83e-20
C1504 a_2060_2640# a_3599_2340# 3.6e-19
C1505 a_2265_2340# a_2200_2366# 9.75e-19
C1506 a_2061_2340# a_2401_2366# 6.04e-20
C1507 a_6010_3239# a_6465_3213# 0.153f
C1508 x30.Q_N check[5] 0.902f
C1509 x4.X a_12737_3239# 0.00277f
C1510 a_10775_2340# a_12101_2550# 4.7e-22
C1511 a_11088_2366# a_11833_2340# 0.199f
C1512 a_11330_2340# a_11629_2340# 0.0334f
C1513 x4.X a_9709_2550# 0.00146f
C1514 check[4] x36.Q_N 8.5e-21
C1515 a_3452_3239# a_3504_2340# 4.5e-19
C1516 x4.X a_4681_4801# 0.00584f
C1517 sel_bit[0] check[1] 0.583f
C1518 check[2] x5.X 0.831f
C1519 clk_sar x5.X 0.00891f
C1520 check[0] a_6780_2366# 1.28e-19
C1521 check[2] a_6292_5167# 5.02e-20
C1522 x4.X a_11857_4801# 0.00316f
C1523 x36.Q_N a_11629_2340# 0.0468f
C1524 VDD x51.Q_N 0.085f
C1525 a_3452_3239# a_4367_3213# 0.125f
C1526 a_3618_3239# a_3899_3605# 0.152f
C1527 D[6] a_4793_2366# 4.25e-19
C1528 a_4453_2340# a_4590_2732# 0.00907f
C1529 a_6010_3239# a_5991_2340# 3.73e-19
C1530 a_8237_4801# a_10629_4801# 0.00176f
C1531 VDD a_3452_3239# 0.821f
C1532 check[6] a_6304_2366# 2.39e-20
C1533 a_11630_4086# a_12030_3213# 7.94e-19
C1534 a_11834_4086# a_11543_3213# 0.0014f
C1535 x39.Q_N a_11249_3213# 0.194f
C1536 check[2] a_9237_4386# 0.163f
C1537 x30.Q_N a_7246_3213# 0.0127f
C1538 a_7247_4775# x72.Q_N 4.45e-20
C1539 sel_bit[0] a_3877_5674# 2.93e-19
C1540 x27.D a_3619_4801# 0.159f
C1541 a_7247_4775# a_7764_4112# 4.23e-19
C1542 a_10156_4112# a_9954_4112# 3.67e-19
C1543 x48.Q a_4971_4801# 4.12e-19
C1544 VDD a_9638_3213# 0.569f
C1545 x20.Q_N a_3170_4801# 0.187f
C1546 a_2697_5083# x27.D 7.73e-21
C1547 a_5896_2340# a_6844_2640# 8.38e-21
C1548 check[0] x77.Y 2.24e-20
C1549 a_8857_3213# a_9322_3521# 9.46e-19
C1550 a_8402_3239# a_9550_3605# 2.13e-19
C1551 a_8236_3239# a_8997_3239# 6.04e-20
C1552 VDD a_6985_4112# 0.00445f
C1553 check[1] check[6] 6.18e-20
C1554 eob x3.A 0.00123f
C1555 x4.X a_9375_4478# 0.00114f
C1556 x42.Q_N a_8236_3239# 0.0435f
C1557 a_8697_4112# a_9464_3239# 2.16e-19
C1558 a_9237_4386# a_9151_3213# 5.72e-19
C1559 a_8384_4086# a_8590_3239# 2.44e-19
C1560 x20.Q_N a_1996_2366# 7.87e-19
C1561 a_897_4112# a_1112_2340# 4.64e-19
C1562 x39.Q_N a_10775_2340# 2.2e-19
C1563 a_10776_4086# x63.Q_N 2.32e-20
C1564 a_11630_4086# a_11628_2640# 7.02e-19
C1565 a_11629_4386# a_11629_2340# 7.25e-19
C1566 x30.Q_N a_6844_2640# 0.57f
C1567 x5.X a_4074_4775# 3.66e-19
C1568 a_2389_5648# a_2579_4801# 2.13e-20
C1569 a_8289_4086# a_9238_4086# 7e-20
C1570 x5.X x20.Q_N 0.00434f
C1571 a_4855_4775# a_5845_4801# 0.00116f
C1572 a_4368_4775# a_6011_4801# 1.1e-19
C1573 x3.A x4.A 4.66e-19
C1574 a_4681_4801# a_3618_3239# 6.75e-21
C1575 x5.X a_11250_4775# 0.00324f
C1576 VDD a_9236_2640# 0.269f
C1577 x4.X a_1996_2732# 4.32e-19
C1578 a_8858_4775# a_8684_5167# 0.205f
C1579 a_8403_4801# a_9152_4775# 0.139f
C1580 a_8237_4801# a_9639_4775# 0.0492f
C1581 D[1] a_12030_3213# 1.69e-20
C1582 a_9464_3239# a_9709_2550# 1.85e-20
C1583 VDD a_3900_5167# 0.324f
C1584 check[2] a_12345_2366# 2.05e-20
C1585 a_6547_4086# a_6291_3605# 1.7e-20
C1586 a_6845_4386# a_6465_3213# 0.0015f
C1587 a_6305_4112# a_6759_3213# 3.33e-20
C1588 a_6846_4086# a_6010_3239# 6.04e-20
C1589 a_4658_4086# a_4925_2550# 2.22e-22
C1590 a_12031_4775# a_12147_4801# 0.0397f
C1591 a_11544_4775# a_11966_4801# 2.87e-21
C1592 a_8939_4086# a_9236_2640# 4.75e-21
C1593 a_8697_4112# a_9237_2340# 1.4e-21
C1594 VDD a_11076_5167# 0.317f
C1595 x48.Q a_4591_4478# 6.11e-19
C1596 x77.Y a_4154_2340# 0.00178f
C1597 x4.X a_897_4112# 1.27e-19
C1598 x27.Q_N a_4789_3239# 1.68e-19
C1599 check[4] a_10345_3239# 0.0274f
C1600 x48.Q a_4214_4801# 0.00132f
C1601 check[6] a_5844_3239# 0.00782f
C1602 a_1338_5674# sel_bit[0] 0.0446f
C1603 VDD a_12345_2732# 0.0042f
C1604 x77.Y a_4538_3521# 2.52e-20
C1605 a_9237_2340# a_9709_2550# 0.15f
C1606 a_9236_2640# x60.Q_N 5.14e-21
C1607 check[2] a_9656_4394# 7.77e-21
C1608 check[0] a_3912_2366# 2.06e-21
C1609 x4.X a_6978_4801# 5.55e-19
C1610 a_4074_4775# a_3984_5167# 6.69e-20
C1611 a_3619_4801# a_2579_4801# 7.73e-20
C1612 a_4368_4775# a_4681_4801# 0.124f
C1613 a_3900_5167# a_3807_4801# 0.0367f
C1614 x30.Q_N x45.Q_N 0.0041f
C1615 check[2] a_9551_5167# 1.87e-19
C1616 x5.X a_8591_4801# 0.00545f
C1617 a_2853_5648# a_2993_5674# 1.56e-19
C1618 a_11629_4386# a_11834_4086# 0.153f
C1619 a_11089_4112# x39.Q_N 0.0933f
C1620 a_2060_2640# a_2979_2366# 0.163f
C1621 a_2265_2340# a_2479_2648# 0.0104f
C1622 a_2061_2340# a_2777_2732# 0.0018f
C1623 a_1762_2340# D[6] 2.05e-19
C1624 D[3] a_11833_2340# 6.82e-20
C1625 check[1] a_6547_4086# 7.52e-20
C1626 x4.X a_10982_3239# 0.00531f
C1627 a_11544_4775# a_11857_4801# 0.124f
C1628 a_11076_5167# a_10983_4801# 0.0367f
C1629 a_11250_4775# a_11160_5167# 6.69e-20
C1630 a_10795_4801# a_9755_4801# 4.87e-21
C1631 VDD a_8768_5167# 0.0042f
C1632 a_4454_4086# a_5372_4112# 0.0664f
C1633 a_4155_4086# a_4389_4112# 0.00707f
C1634 a_4658_4086# a_5170_4478# 6.69e-20
C1635 a_3913_4112# a_4593_4112# 3.73e-19
C1636 a_4453_4386# a_5897_4086# 3.56e-19
C1637 check[0] a_6410_2366# 0.00226f
C1638 a_8384_4086# a_9173_4478# 7.71e-20
C1639 a_8697_4112# a_8897_4394# 0.00185f
C1640 x27.Q_N a_4454_4086# 0.0256f
C1641 a_8684_5167# x42.Q_N 9.99e-20
C1642 a_9639_4775# a_9442_4086# 4.44e-19
C1643 a_9152_4775# a_9710_4296# 2.85e-19
C1644 sel_bit[0] a_3453_4801# 4.34e-20
C1645 a_3912_2366# a_4154_2340# 0.124f
C1646 a_3599_2340# a_4452_2640# 0.0264f
C1647 a_3504_2340# x54.Q_N 0.178f
C1648 a_6759_3213# a_6605_3239# 0.00943f
C1649 a_6291_3605# a_6399_3239# 0.00812f
C1650 a_7072_3239# a_6930_3521# 0.00412f
C1651 a_6465_3213# a_6977_3239# 9.75e-19
C1652 a_7246_3213# a_7158_3605# 7.71e-20
C1653 x4.X a_11833_2340# 0.00145f
C1654 sel_bit[1] a_1682_4775# 1.09e-19
C1655 x5.X a_7953_3239# 0.00125f
C1656 x36.Q_N a_12548_4112# 0.0133f
C1657 a_6411_4112# a_6291_3605# 1.12e-20
C1658 x4.X a_4593_4112# 0.0012f
C1659 check[6] D[5] 0.141f
C1660 a_6547_4086# a_7050_4086# 0.00187f
C1661 a_5992_4086# x45.Q_N 0.154f
C1662 a_6845_4386# a_6846_4086# 0.75f
C1663 a_6305_4112# a_7318_4296# 0.0633f
C1664 a_4854_3213# a_4925_2550# 1.66e-21
C1665 a_4680_3239# a_4657_2340# 1.03e-19
C1666 a_6305_4112# comparator_out 2.29e-20
C1667 x5.X a_6931_5083# 5.11e-19
C1668 VDD D[0] 0.301f
C1669 check[2] x30.Q_N 6.73e-21
C1670 VDD x54.Q_N 0.0807f
C1671 a_4925_2550# a_5169_2366# 0.00812f
C1672 a_6199_4801# a_6376_5167# 8.94e-19
C1673 a_6011_4801# a_6606_4801# 0.00118f
C1674 a_6760_4775# a_6710_5083# 1.21e-20
C1675 a_4367_3213# a_5088_3521# 0.00185f
C1676 check[0] a_4539_5083# 4.79e-19
C1677 D[0] a_7362_3239# 8.51e-20
C1678 a_9639_4775# a_9574_4801# 4.2e-20
C1679 a_9465_4801# a_9755_4801# 0.0282f
C1680 a_1511_4112# a_1207_2340# 1.58e-19
C1681 a_6411_4112# a_6304_2366# 8.38e-21
C1682 VDD a_7159_5167# 0.00371f
C1683 VDD a_5088_3521# 0.00529f
C1684 x20.Q_N a_1626_2366# 0.00967f
C1685 x39.Q_N a_11965_3239# 7.87e-19
C1686 x30.Q_N a_9151_3213# 8.28e-21
C1687 x33.Q_N a_9953_2366# 0.00224f
C1688 x39.Q_N a_12264_3521# 2.75e-19
C1689 a_3619_4801# a_5562_4801# 1.64e-20
C1690 a_3453_4801# check[6] 8.06e-20
C1691 VDD a_11543_3213# 0.352f
C1692 eob a_1227_4801# 0.413f
C1693 a_11629_4386# a_12548_4112# 0.163f
C1694 a_11331_4086# a_11565_4112# 0.00707f
C1695 a_11834_4086# a_12048_4394# 0.0104f
C1696 a_11089_4112# a_11769_4112# 3.73e-19
C1697 a_11630_4086# a_12346_4478# 0.0018f
C1698 check[5] a_8237_4801# 0.414f
C1699 a_7954_4801# a_8403_4801# 5.4e-19
C1700 a_6304_2366# a_6780_2366# 2.87e-21
C1701 a_9151_3213# a_9754_3239# 0.0552f
C1702 check[1] a_6411_4112# 1.13e-20
C1703 check[2] a_3373_5674# 0.0404f
C1704 a_10795_4801# a_12738_4801# 8.38e-21
C1705 a_10629_4801# check[3] 0.00126f
C1706 check[4] a_12147_4801# 1.37e-20
C1707 a_1227_4801# x4.A 0.00377f
C1708 check[2] x63.Q_N 0.0121f
C1709 comparator_out a_1207_2340# 6.22e-19
C1710 x27.Q_N a_3504_2340# 3.7e-19
C1711 check[2] a_5992_4086# 3.43e-20
C1712 x5.X a_5170_4478# 1.85e-19
C1713 x4.X a_12102_4296# 0.021f
C1714 x48.Q a_1511_4112# 0.00368f
C1715 x30.Q_N a_8938_2340# 5.93e-20
C1716 a_1508_5167# a_1415_4801# 0.0367f
C1717 a_1976_4775# a_2289_4801# 0.124f
C1718 VDD a_11330_2340# 0.177f
C1719 a_9639_4775# a_10156_4112# 4.23e-19
C1720 x27.Q_N a_4367_3213# 0.00484f
C1721 x27.Q_N a_6466_4775# 1.88e-20
C1722 x4.X a_4112_2648# 0.00102f
C1723 a_8383_2340# a_8896_2648# 0.00945f
C1724 x5.X a_12265_5083# 1.33e-19
C1725 VDD a_5372_4112# 0.11f
C1726 a_11543_3213# D[2] 3.13e-19
C1727 a_12030_3213# a_12737_3239# 0.0968f
C1728 x4.X a_6709_3521# 2.91e-19
C1729 a_8858_4775# x33.Q_N 2.07e-20
C1730 a_9465_4801# a_8998_4801# 0.00316f
C1731 a_9152_4775# a_9370_4801# 3.73e-19
C1732 VDD x27.Q_N 0.452f
C1733 x4.X a_5170_4112# 7.21e-19
C1734 x45.Q_N a_7158_3605# 3.63e-19
C1735 x48.Q a_1061_4801# 4.14e-21
C1736 x4.X a_5561_3239# 0.00286f
C1737 a_6846_4086# a_7264_4394# 0.00276f
C1738 a_6845_4386# a_7562_4478# 4.45e-20
C1739 a_5992_4086# a_6781_4112# 4.2e-20
C1740 VDD x36.Q_N 0.419f
C1741 x48.Q comparator_out 3.3e-20
C1742 check[4] a_9441_2340# 7.03e-20
C1743 a_12031_4775# a_11856_3239# 1.33e-23
C1744 a_11857_4801# a_12030_3213# 4.82e-21
C1745 check[1] a_9953_2366# 2.06e-20
C1746 eob a_2533_2550# 4.21e-20
C1747 a_7247_4775# check[5] 0.0104f
C1748 a_1520_2366# a_2061_2340# 0.125f
C1749 a_1762_2340# a_2060_2640# 0.137f
C1750 check[2] eob 0.0123f
C1751 D[2] a_11330_2340# 2.3e-20
C1752 clk_sar eob 4.74e-20
C1753 check[4] a_12031_4775# 1.91e-20
C1754 comparator_out a_8288_2340# 7.84e-19
C1755 a_1061_4801# a_2147_5083# 0.00907f
C1756 a_1682_4775# a_1592_5167# 6.69e-20
C1757 x4.X a_1415_4801# 9.23e-21
C1758 a_4155_4086# a_4454_4086# 0.0334f
C1759 a_3913_4112# a_4658_4086# 0.199f
C1760 a_3600_4086# a_4926_4296# 4.7e-22
C1761 a_3505_4086# x48.Q_N 0.178f
C1762 check[0] a_5991_2340# 0.0146f
C1763 x5.X a_11331_4086# 8.88e-19
C1764 x36.Q_N D[2] 0.00122f
C1765 a_3807_4801# x27.Q_N 5.03e-21
C1766 a_11195_4112# a_11565_4112# 4.11e-20
C1767 D[6] a_4154_2340# 8.45e-19
C1768 a_12101_2550# a_12345_2732# 0.00972f
C1769 a_11330_2340# a_11969_2366# 0.00316f
C1770 a_11833_2340# a_12547_2366# 6.99e-20
C1771 a_11628_2640# a_11768_2366# 0.00126f
C1772 a_12147_4801# a_11834_4086# 7.76e-20
C1773 VDD a_11629_4386# 0.59f
C1774 x4.X a_4658_4086# 0.0102f
C1775 a_10983_4801# x36.Q_N 5.41e-22
C1776 check[6] a_4453_2340# 0.0409f
C1777 a_10681_4086# a_10628_3239# 5.06e-19
C1778 a_7247_4775# a_7246_3213# 0.00237f
C1779 a_2853_5648# check[0] 0.164f
C1780 a_4854_3213# a_6198_3239# 8.26e-21
C1781 x4.X a_11565_4112# 8.15e-20
C1782 x39.Q_N a_9638_3213# 3.76e-21
C1783 a_2389_5648# x48.Q 0.00138f
C1784 x33.Q_N a_8997_3239# 6.08e-19
C1785 a_9238_4086# a_11089_4112# 5.07e-21
C1786 a_9710_4296# a_9578_4112# 0.0258f
C1787 a_9237_4386# a_11331_4086# 2.53e-20
C1788 x42.Q_N a_9377_4112# 0.00167f
C1789 x36.Q_N a_11969_2366# 0.0403f
C1790 VDD a_6375_3605# 0.0042f
C1791 x77.Y a_5844_3239# 2.13e-19
C1792 a_3452_3239# x75.Q 6.31e-20
C1793 a_3618_3239# a_5561_3239# 3.23e-21
C1794 a_5169_2732# a_5371_2366# 8.94e-19
C1795 x33.Q_N x42.Q_N 0.00395f
C1796 a_8236_3239# a_8402_3239# 0.782f
C1797 a_4154_2340# a_5991_2340# 1.86e-21
C1798 a_4452_2640# a_4793_2366# 0.00118f
C1799 a_4453_2340# a_4592_2366# 2.56e-19
C1800 a_3912_2366# a_6304_2366# 8.41e-21
C1801 a_7480_3521# a_8236_3239# 4.06e-20
C1802 sel_bit[0] x3.A 6.99e-21
C1803 check[5] a_9574_4801# 1.69e-20
C1804 eob x20.Q_N 0.365f
C1805 a_11630_4086# a_12737_3239# 4.72e-19
C1806 x30.Q_N a_7953_3239# 0.00834f
C1807 x5.X a_1508_5167# 0.00288f
C1808 check[0] a_3671_5674# 3.04e-19
C1809 x27.D a_3600_4086# 0.00292f
C1810 x33.Q_N a_10680_2340# 1.87e-19
C1811 check[3] a_10794_3239# 1.56e-21
C1812 x20.Q_N x4.A 5.76e-19
C1813 VDD a_10345_3239# 0.19f
C1814 check[0] a_6846_4086# 2.15e-19
C1815 VDD a_7317_2550# 0.172f
C1816 a_8403_4801# comparator_out 2.9e-21
C1817 a_6304_2366# a_6410_2366# 0.0552f
C1818 a_6546_2340# a_6982_2732# 0.00412f
C1819 a_6844_2640# a_6780_2732# 2.13e-19
C1820 a_6845_2340# a_6504_2648# 1.25e-19
C1821 D[5] a_6780_2366# 3.51e-20
C1822 a_6606_4801# a_6978_4801# 3.34e-19
C1823 a_12031_4775# a_11834_4086# 4.44e-19
C1824 a_11544_4775# a_12102_4296# 2.85e-19
C1825 a_11076_5167# x39.Q_N 1e-19
C1826 a_7362_3239# a_7317_2550# 1.01e-20
C1827 VDD a_1976_4775# 0.489f
C1828 x5.X D[3] 3.43e-19
C1829 a_8289_4086# a_8288_2340# 1.07e-20
C1830 x4.X a_3170_4801# 9.94e-19
C1831 a_1682_4775# x27.D 2.67e-21
C1832 x5.X a_3913_4112# 1.32e-19
C1833 a_4658_4086# a_3618_3239# 2.9e-19
C1834 a_4454_4086# a_4073_3213# 5.04e-19
C1835 a_3913_4112# a_4854_3213# 9.49e-19
C1836 a_4155_4086# a_4367_3213# 2.12e-19
C1837 x48.Q a_3619_4801# 0.0352f
C1838 check[2] a_11970_4112# 3.49e-20
C1839 VDD D[7] 0.225f
C1840 a_6984_2366# a_7185_2366# 3.34e-19
C1841 a_8288_2340# a_8696_2366# 6.04e-19
C1842 VDD a_4155_4086# 0.348f
C1843 a_10628_3239# a_11714_3521# 0.00907f
C1844 a_10794_3239# a_11493_3521# 2.46e-19
C1845 check[5] a_8792_4801# 1.67e-19
C1846 check[1] x42.Q_N 0.0239f
C1847 VDD a_12048_4394# 0.00984f
C1848 x5.X x4.X 0.0429f
C1849 x42.Q_N a_8802_2366# 4.74e-20
C1850 comparator_out a_3599_2340# 0.00328f
C1851 x4.X a_6292_5167# 0.00132f
C1852 x4.X a_4854_3213# 0.117f
C1853 a_10156_4112# a_10776_4086# 8.26e-21
C1854 a_1976_4775# a_3807_4801# 2.23e-21
C1855 a_2463_4775# a_4681_4801# 1.86e-21
C1856 check[2] a_8237_4801# 5.48e-19
C1857 a_7073_4801# a_7318_4296# 3.59e-20
C1858 a_9237_4386# a_11195_4112# 1.71e-20
C1859 x42.Q_N a_9954_4112# 2.4e-19
C1860 a_12030_3213# a_11833_2340# 2.52e-19
C1861 a_11543_3213# a_12101_2550# 1.62e-19
C1862 x4.X a_7181_3239# 1.05e-19
C1863 a_9873_5083# x33.Q_N 2.02e-20
C1864 comparator_out a_6982_2732# 9.43e-19
C1865 x4.X a_9237_4386# 0.048f
C1866 a_8858_4775# a_8857_3213# 2.59e-19
C1867 a_8403_4801# a_8683_3605# 8.52e-21
C1868 a_8684_5167# a_8402_3239# 1.65e-21
C1869 a_9152_4775# a_8236_3239# 9.66e-21
C1870 a_4368_4775# a_4658_4086# 0.00268f
C1871 a_4855_4775# a_4454_4086# 0.00169f
C1872 a_4681_4801# a_4453_4386# 1.96e-20
C1873 a_7050_4086# x42.Q_N 1.92e-20
C1874 check[4] a_11629_2340# 1.57e-21
C1875 x20.Q_N x48.Q_N 0.00138f
C1876 a_3453_4801# x77.Y 9.38e-22
C1877 a_6465_3213# a_6291_3605# 0.205f
C1878 a_6010_3239# a_6759_3213# 0.139f
C1879 a_2060_2640# a_4154_2340# 4.16e-20
C1880 a_2061_2340# a_3912_2366# 3.12e-19
C1881 a_2533_2550# a_2401_2366# 0.0258f
C1882 a_12031_4775# a_12548_4112# 4.23e-19
C1883 check[3] a_10776_4086# 1.93e-20
C1884 a_11088_2366# x63.Q_N 0.00553f
C1885 a_11628_2640# a_11833_2340# 0.153f
C1886 check[0] a_7185_2366# 4.21e-19
C1887 check[2] a_7247_4775# 2.07e-19
C1888 x36.Q_N a_12101_2550# 0.181f
C1889 a_4073_3213# a_4367_3213# 0.198f
C1890 a_5845_4801# a_6466_4775# 0.117f
C1891 a_3452_3239# a_4680_3239# 0.0334f
C1892 a_3618_3239# a_4854_3213# 0.0264f
C1893 a_3912_2366# D[5] 2.89e-20
C1894 a_4452_2640# a_5169_2732# 4.45e-20
C1895 a_4453_2340# a_4871_2648# 0.00276f
C1896 a_6465_3213# a_6304_2366# 0.0014f
C1897 a_6291_3605# a_5991_2340# 3.9e-20
C1898 check[1] a_9173_4112# 1.03e-21
C1899 VDD a_5845_4801# 0.81f
C1900 VDD a_4073_3213# 0.314f
C1901 a_12102_4296# a_12030_3213# 3.74e-20
C1902 a_11834_4086# a_11856_3239# 4.33e-20
C1903 x39.Q_N a_11543_3213# 0.0983f
C1904 VDD a_12147_4801# 0.0101f
C1905 check[2] a_9442_4086# 7.66e-19
C1906 sel_bit[0] a_1227_4801# 2.06e-20
C1907 x27.D a_3900_5167# 8.53e-19
C1908 VDD a_8590_3239# 0.109f
C1909 x75.Q_N a_5561_3239# 0.178f
C1910 D[5] a_6410_2366# 5.42e-19
C1911 a_8236_3239# a_10628_3239# 0.00176f
C1912 a_5991_2340# a_6304_2366# 0.273f
C1913 a_8402_3239# a_8791_3239# 0.0019f
C1914 a_9151_3213# a_9322_3521# 0.00652f
C1915 a_8857_3213# a_8997_3239# 0.07f
C1916 a_8236_3239# a_9369_3239# 2.56e-19
C1917 a_1511_4112# a_2979_2366# 3.09e-20
C1918 VDD a_8384_4086# 0.716f
C1919 x5.X a_9237_2340# 2.59e-20
C1920 a_9442_4086# a_9151_3213# 0.0014f
C1921 a_9238_4086# a_9638_3213# 7.94e-19
C1922 x42.Q_N a_8857_3213# 0.194f
C1923 x4.X a_9656_4394# 8.47e-19
C1924 x20.Q_N a_2401_2366# 0.0313f
C1925 x39.Q_N a_11330_2340# 0.0018f
C1926 a_12102_4296# a_11628_2640# 6.02e-22
C1927 a_11629_4386# a_12101_2550# 6.45e-21
C1928 x30.Q_N a_7049_2340# 0.179f
C1929 x5.X a_4368_4775# 4.59e-19
C1930 a_8384_4086# a_8939_4086# 0.197f
C1931 a_7764_4112# x42.Q_N 5.48e-20
C1932 a_10681_4086# comparator_out 2.05e-21
C1933 a_3453_4801# a_6199_4801# 3.65e-21
C1934 a_4855_4775# a_4367_3213# 1.08e-22
C1935 a_4368_4775# a_4854_3213# 1.06e-20
C1936 a_4681_4801# a_6011_4801# 3.02e-20
C1937 VDD a_9441_2340# 0.304f
C1938 x5.X a_11544_4775# 0.00155f
C1939 x20.Q_N a_3806_3239# 0.00103f
C1940 x4.X a_1626_2366# 3.78e-20
C1941 D[4] a_8288_2340# 0.1f
C1942 D[1] a_10982_3239# 4.96e-19
C1943 a_8403_4801# a_9465_4801# 0.137f
C1944 a_8684_5167# a_9152_4775# 0.0633f
C1945 a_8237_4801# a_8591_4801# 0.0664f
C1946 a_8997_3239# a_8383_2340# 4.6e-20
C1947 VDD a_4855_4775# 0.723f
C1948 x36.Q_N x39.Q_N 0.00386f
C1949 a_6305_4112# a_7072_3239# 2.16e-19
C1950 a_6845_4386# a_6759_3213# 5.72e-19
C1951 a_5992_4086# a_6198_3239# 2.44e-19
C1952 a_5844_3239# a_6465_3213# 0.117f
C1953 comparator_out a_2979_2366# 0.157f
C1954 comparator_out a_6010_3239# 0.149f
C1955 a_11857_4801# a_11966_4801# 0.00707f
C1956 x42.Q_N a_8383_2340# 2.17e-19
C1957 a_9237_4386# a_9237_2340# 7.25e-19
C1958 a_9238_4086# a_9236_2640# 7.02e-19
C1959 a_8384_4086# x60.Q_N 2.32e-20
C1960 VDD a_12031_4775# 0.709f
C1961 x77.Y a_4453_2340# 3.65e-20
C1962 x48.Q a_4872_4394# 1.99e-19
C1963 check[6] x45.Q_N 6.19e-19
C1964 a_2853_5648# check[1] 0.0514f
C1965 x48.Q a_4586_4801# 3.31e-19
C1966 check[2] sel_bit[0] 0.0781f
C1967 clk_sar sel_bit[0] 0.343f
C1968 x77.Y a_4213_3239# 0.0313f
C1969 x4.X a_5896_2340# 0.00507f
C1970 a_6547_4086# a_6844_2640# 4.75e-21
C1971 a_6305_4112# a_6845_2340# 1.4e-21
C1972 a_5844_3239# a_5991_2340# 8.35e-19
C1973 sel_bit[1] a_1976_4775# 8.83e-20
C1974 check[0] a_4452_2640# 2.1e-19
C1975 check[2] a_10156_4112# 0.165f
C1976 x5.X a_8897_4394# 5.64e-19
C1977 x4.X x30.Q_N 0.426f
C1978 a_3453_4801# a_4539_5083# 0.00907f
C1979 a_3619_4801# a_4318_5083# 2.46e-19
C1980 x20.Q_N a_2398_4801# 9.16e-20
C1981 a_11630_4086# a_12102_4296# 0.15f
C1982 x5.X a_7363_4801# 2.04e-19
C1983 a_11629_4386# x39.Q_N 0.00118f
C1984 a_2853_5648# a_3877_5674# 8.24e-20
C1985 check[1] a_3671_5674# 5.38e-19
C1986 a_2061_2340# D[6] 0.338f
C1987 a_2533_2550# a_2777_2732# 0.00972f
C1988 a_2265_2340# a_2979_2366# 6.99e-20
C1989 a_7247_4775# a_8591_4801# 8.26e-21
C1990 D[3] x63.Q_N 0.00107f
C1991 check[1] a_6846_4086# 0.441f
C1992 VDD a_9173_4478# 0.00371f
C1993 x4.X a_9754_3239# 5.61e-19
C1994 a_10629_4801# a_11715_5083# 0.00907f
C1995 comparator_out a_9172_2732# 1.81e-19
C1996 a_10795_4801# a_11494_5083# 2.46e-19
C1997 VDD a_7182_4801# 7.87e-19
C1998 check[5] a_6780_2366# 2.23e-20
C1999 a_4155_4086# a_4794_4112# 0.00316f
C2000 a_4926_4296# a_5372_4112# 0.0367f
C2001 a_4453_4386# a_4593_4112# 0.00126f
C2002 a_11970_4112# a_11088_2366# 1.26e-20
C2003 x33.Q_N a_8402_3239# 3.88e-19
C2004 a_8697_4112# a_9375_4478# 0.00652f
C2005 a_8939_4086# a_9173_4478# 0.00976f
C2006 check[2] check[6] 7.32e-20
C2007 a_8384_4086# a_8803_4112# 0.0397f
C2008 a_4019_4112# x77.Y 1.79e-19
C2009 VDD a_1720_2648# 0.00736f
C2010 x27.Q_N a_4926_4296# 5.7e-19
C2011 a_9465_4801# a_9710_4296# 3.59e-20
C2012 a_6759_3213# a_8236_3239# 3.41e-19
C2013 sel_bit[0] a_4074_4775# 0.00112f
C2014 a_4154_2340# a_4452_2640# 0.137f
C2015 a_3912_2366# a_4453_2340# 0.125f
C2016 a_11564_2366# a_11969_2366# 2.46e-21
C2017 a_12547_2366# a_12345_2366# 3.67e-19
C2018 a_6759_3213# a_6977_3239# 3.73e-19
C2019 a_7072_3239# a_6605_3239# 0.00316f
C2020 sel_bit[0] x20.Q_N 2.7e-20
C2021 a_3373_5674# x4.X 5.96e-20
C2022 x4.X x63.Q_N 0.00782f
C2023 eob a_1508_5167# 0.0514f
C2024 x4.X a_5992_4086# 0.1f
C2025 a_7247_4775# a_7953_3239# 4.94e-20
C2026 a_6845_4386# a_7318_4296# 0.155f
C2027 a_6547_4086# x45.Q_N 0.0285f
C2028 a_6846_4086# a_7050_4086# 0.117f
C2029 a_6845_4386# comparator_out 2.52e-20
C2030 a_6846_4086# a_5844_3239# 6.54e-20
C2031 a_1508_5167# x4.A 0.00373f
C2032 check[0] a_4591_4478# 1.2e-20
C2033 x5.X a_6606_4801# 9.34e-19
C2034 eob a_1112_2340# 3.79e-20
C2035 a_4854_3213# x75.Q_N 0.124f
C2036 a_6760_4775# a_7159_5167# 0.00133f
C2037 a_5845_4801# a_7481_5083# 1.25e-19
C2038 a_6011_4801# a_6978_4801# 0.00126f
C2039 a_6292_5167# a_6606_4801# 0.0258f
C2040 D[5] a_5991_2340# 0.0123f
C2041 a_5371_2366# a_6304_2366# 3.42e-20
C2042 a_1338_5674# a_2853_5648# 5.64e-20
C2043 a_1511_4112# a_1762_2340# 4.16e-20
C2044 a_9873_5083# a_10629_4801# 4.06e-20
C2045 x4.A a_1112_2340# 7.47e-22
C2046 x20.Q_N a_2777_2732# 8.48e-19
C2047 a_4074_4775# check[6] 4.81e-21
C2048 check[1] a_8402_3239# 0.0363f
C2049 a_12102_4296# a_12346_4478# 0.00972f
C2050 a_11331_4086# a_11970_4112# 0.00316f
C2051 a_11834_4086# a_12548_4112# 6.99e-20
C2052 a_11629_4386# a_11769_4112# 0.00126f
C2053 VDD a_11856_3239# 0.18f
C2054 x5.X a_10346_4801# 0.0293f
C2055 eob x4.X 0.22f
C2056 a_6546_2340# a_6984_2366# 0.00276f
C2057 a_6304_2366# a_7185_2366# 0.00943f
C2058 a_6845_2340# a_8288_2340# 8.18e-19
C2059 check[5] a_8858_4775# 6.94e-19
C2060 a_9464_3239# a_9754_3239# 0.0282f
C2061 a_9638_3213# a_9573_3239# 4.2e-20
C2062 a_4019_4112# a_3912_2366# 8.38e-21
C2063 check[2] a_2788_5674# 0.00675f
C2064 a_11250_4775# check[3] 0.00109f
C2065 comparator_out a_1762_2340# 1.88e-19
C2066 a_4658_4086# a_4970_3239# 5.48e-21
C2067 x4.X x4.A 0.00766f
C2068 x42.Q_N a_10794_3239# 9.16e-19
C2069 VDD check[4] 0.5f
C2070 a_4453_4386# a_5170_4112# 0.0019f
C2071 x42.Q_N a_9872_3521# 2.75e-19
C2072 x5.X a_5897_4086# 0.0764f
C2073 x48.Q a_3600_4086# 0.00969f
C2074 x30.Q_N a_9237_2340# 8.11e-21
C2075 VDD a_11629_2340# 0.784f
C2076 VDD a_2883_5674# 0.172f
C2077 x27.Q_N a_6760_4775# 6.16e-21
C2078 x27.Q_N a_4680_3239# 0.0029f
C2079 a_8696_2366# a_9172_2732# 0.00133f
C2080 x4.X a_4590_2732# 9.81e-19
C2081 a_11856_3239# D[2] 5.2e-20
C2082 VDD a_4389_4112# 9.51e-19
C2083 x4.X a_7158_3605# 4.4e-19
C2084 a_9152_4775# x33.Q_N 0.0059f
C2085 a_9639_4775# a_9873_5083# 0.00945f
C2086 a_8591_4801# a_8792_4801# 3.67e-19
C2087 a_9465_4801# a_9370_4801# 0.00276f
C2088 a_2853_5648# a_3453_4801# 7.76e-20
C2089 comparator_out a_5169_2732# 8.25e-19
C2090 a_5844_3239# a_8402_3239# 2.9e-21
C2091 x4.X a_6781_4478# 2.12e-19
C2092 comparator_out a_8236_3239# 0.147f
C2093 x42.Q_N a_9577_2366# 5.33e-22
C2094 x48.Q a_1682_4775# 4.88e-21
C2095 a_5844_3239# a_7480_3521# 1.25e-19
C2096 a_7050_4086# a_7562_4478# 6.69e-20
C2097 a_6846_4086# a_7764_4112# 0.0664f
C2098 x45.Q_N a_6411_4112# 0.0455f
C2099 a_6845_4386# a_8289_4086# 4.36e-19
C2100 a_6547_4086# a_6781_4112# 0.00707f
C2101 a_6305_4112# a_6985_4112# 3.73e-19
C2102 check[0] a_6759_3213# 1.67e-20
C2103 a_1822_4801# a_1511_4112# 1.33e-19
C2104 a_1520_2366# a_2533_2550# 0.0633f
C2105 a_2060_2640# a_2061_2340# 0.783f
C2106 a_1207_2340# x51.Q_N 0.124f
C2107 a_1762_2340# a_2265_2340# 0.00187f
C2108 D[2] a_11629_2340# 0.271f
C2109 a_9237_2340# x63.Q_N 2.94e-19
C2110 check[4] a_10983_4801# 0.164f
C2111 check[5] a_6410_2366# 1.31e-19
C2112 a_1061_4801# a_1822_4801# 6.04e-20
C2113 a_1682_4775# a_2147_5083# 9.46e-19
C2114 a_1227_4801# a_2375_5167# 2.13e-19
C2115 a_4453_4386# a_4658_4086# 0.153f
C2116 a_3913_4112# x48.Q_N 0.00553f
C2117 a_4855_4775# a_4794_4112# 1.79e-20
C2118 check[0] a_6546_2340# 0.00104f
C2119 a_3505_4086# x77.Y 7.15e-21
C2120 x5.X a_11630_4086# 0.26f
C2121 a_621_4112# a_1511_4112# 2.76e-19
C2122 check[5] x42.Q_N 6.88e-19
C2123 D[6] a_4453_2340# 2.08e-19
C2124 a_11628_2640# a_12345_2366# 0.00105f
C2125 a_11833_2340# a_11768_2366# 9.75e-19
C2126 a_11629_2340# a_11969_2366# 6.04e-20
C2127 x30.Q_N a_7363_4801# 0.00129f
C2128 comparator_out a_11288_2648# 1.53e-19
C2129 VDD a_11834_4086# 0.487f
C2130 x4.X x48.Q_N 0.00819f
C2131 check[6] a_4925_2550# 9.23e-19
C2132 a_4367_3213# a_4789_3239# 2.87e-21
C2133 a_4854_3213# a_4970_3239# 0.0397f
C2134 x4.X a_11970_4112# 0.00309f
C2135 x33.Q_N a_10628_3239# 8.92e-20
C2136 VDD a_2777_2366# 8.32e-19
C2137 a_2463_4775# a_3170_4801# 0.0968f
C2138 x48.Q a_3452_3239# 8.21e-19
C2139 x42.Q_N a_10776_4086# 7.84e-21
C2140 a_9237_4386# a_11630_4086# 2.9e-21
C2141 x45.Q_N x77.Y 1.27e-22
C2142 a_1976_4775# x27.D 0.00388f
C2143 x33.Q_N a_9369_3239# 4.04e-19
C2144 a_5845_4801# x75.Q 1.99e-20
C2145 VDD a_4789_3239# 1.15e-19
C2146 check[6] a_6931_5083# 1.5e-21
C2147 a_8402_3239# a_8857_3213# 0.153f
C2148 a_8236_3239# a_8683_3605# 0.15f
C2149 a_621_4112# comparator_out 1.4e-20
C2150 a_4453_2340# a_5991_2340# 0.00116f
C2151 a_4657_2340# a_4793_2366# 0.07f
C2152 a_4452_2640# a_6304_2366# 1.95e-19
C2153 x72.Q_N a_8402_3239# 9.24e-20
C2154 a_7480_3521# x72.Q_N 2.02e-20
C2155 x5.X D[1] 0.00133f
C2156 a_8289_4086# a_8236_3239# 5.06e-19
C2157 x42.Q_N a_7246_3213# 3.76e-21
C2158 a_10776_4086# a_10680_2340# 2.97e-20
C2159 a_10681_4086# a_10775_2340# 1.57e-20
C2160 x20.Q_N a_1520_2366# 0.0983f
C2161 a_7562_4478# a_7764_4112# 8.94e-19
C2162 a_6411_4112# a_6781_4112# 4.11e-20
C2163 x4.X a_8237_4801# 0.0043f
C2164 x5.X a_2463_4775# 0.016f
C2165 x33.Q_N a_9376_2366# 0.00473f
C2166 check[0] a_7318_4296# 4.24e-20
C2167 check[0] comparator_out 0.121f
C2168 a_6845_2340# a_6982_2732# 0.00907f
C2169 D[5] a_7185_2366# 7.82e-20
C2170 a_8402_3239# a_8383_2340# 3.73e-19
C2171 a_8236_3239# a_8696_2366# 1.89e-19
C2172 D[7] a_2200_2366# 3.49e-19
C2173 D[0] a_9573_3239# 1.29e-20
C2174 a_11857_4801# a_12102_4296# 3.59e-20
C2175 a_6606_4801# x30.Q_N 1.33e-19
C2176 a_3600_4086# a_3599_2340# 5.27e-19
C2177 VDD a_2289_4801# 0.203f
C2178 a_9238_4086# a_10345_3239# 4.72e-19
C2179 x33.Q_N a_11390_4801# 6.84e-20
C2180 x5.X a_4453_4386# 0.009f
C2181 check[3] a_11088_2366# 1.09e-20
C2182 a_4454_4086# a_4367_3213# 1.61e-19
C2183 a_4453_4386# a_4854_3213# 3.78e-19
C2184 x48.Q a_3900_5167# 0.00702f
C2185 x27.Q_N a_5562_4801# 0.182f
C2186 a_5089_5083# check[6] 5.84e-21
C2187 a_8288_2340# a_9236_2640# 9.02e-21
C2188 VDD a_4454_4086# 0.809f
C2189 a_11249_3213# a_11714_3521# 9.46e-19
C2190 a_10794_3239# a_11942_3605# 2.13e-19
C2191 a_10628_3239# a_11389_3239# 6.04e-20
C2192 a_5897_4086# a_5896_2340# 1.07e-20
C2193 VDD a_12548_4112# 0.109f
C2194 comparator_out a_4154_2340# 0.00109f
C2195 x27.Q_N a_4388_2366# 9.43e-19
C2196 x36.Q_N a_12738_4801# 0.184f
C2197 a_12265_5083# check[3] 0.0011f
C2198 x4.X a_3806_3239# 0.00861f
C2199 x4.X a_7247_4775# 0.103f
C2200 a_9377_4112# a_9578_4112# 3.34e-19
C2201 a_10681_4086# a_11089_4112# 4.37e-19
C2202 a_6606_4801# a_5992_4086# 1.08e-19
C2203 check[2] a_8858_4775# 5.69e-19
C2204 a_1976_4775# a_2579_4801# 0.0551f
C2205 check[1] a_9376_2366# 3.33e-19
C2206 x4.X a_6780_2732# 4.32e-19
C2207 a_11856_3239# a_12101_2550# 1.85e-20
C2208 x4.X a_9322_3521# 9.99e-19
C2209 x45.Q_N a_6410_2366# 4.18e-20
C2210 comparator_out a_7263_2648# 6.92e-19
C2211 x4.X a_9442_4086# 0.00986f
C2212 check[5] a_5991_2340# 2.6e-20
C2213 a_8858_4775# a_9151_3213# 7.57e-21
C2214 a_8237_4801# a_9464_3239# 4.76e-21
C2215 a_4855_4775# a_4926_4296# 2.97e-21
C2216 a_4681_4801# a_4658_4086# 2.59e-19
C2217 a_4074_4775# x77.Y 5.16e-21
C2218 x20.Q_N x77.Y 0.0156f
C2219 a_6291_3605# a_6759_3213# 0.0633f
C2220 a_6010_3239# a_7072_3239# 0.137f
C2221 sel_bit[0] a_1508_5167# 3.52e-20
C2222 a_2060_2640# a_4453_2340# 2.9e-21
C2223 a_2061_2340# a_4452_2640# 4e-20
C2224 a_2533_2550# a_3912_2366# 6.92e-21
C2225 a_2883_5674# a_3258_5648# 0.014f
C2226 check[3] a_11331_4086# 4.58e-20
C2227 a_11629_2340# a_12101_2550# 0.15f
C2228 a_11628_2640# x63.Q_N 5.46e-21
C2229 a_2883_5674# sel_bit[1] 0.0353f
C2230 check[1] a_7954_4801# 0.0169f
C2231 a_3452_3239# a_3599_2340# 8.35e-19
C2232 a_5897_4086# a_5992_4086# 0.0968f
C2233 a_4389_4112# a_4794_4112# 2.46e-21
C2234 x4.X a_2398_4801# 0.00124f
C2235 x5.X a_6011_4801# 0.0199f
C2236 VDD a_3504_2340# 0.205f
C2237 x4.X a_9574_4801# 2.39e-19
C2238 sel_bit[0] a_3913_4112# 5.05e-19
C2239 a_3899_3605# a_4854_3213# 4.7e-22
C2240 a_4073_3213# a_4680_3239# 0.00187f
C2241 a_6011_4801# a_6292_5167# 0.155f
C2242 a_5845_4801# a_6760_4775# 0.125f
C2243 a_3618_3239# a_3806_3239# 0.159f
C2244 a_3452_3239# a_3983_3605# 0.0018f
C2245 a_4452_2640# D[5] 0.00524f
C2246 a_4657_2340# a_5169_2732# 6.69e-20
C2247 a_4453_2340# a_5371_2366# 0.0708f
C2248 check[0] a_3619_4801# 0.00149f
C2249 x5.X a_11966_4801# 5.38e-20
C2250 a_6291_3605# a_6546_2340# 2.41e-20
C2251 a_6759_3213# a_6304_2366# 3.36e-20
C2252 a_6010_3239# a_6845_2340# 6.38e-20
C2253 a_6465_3213# a_6844_2640# 2.68e-19
C2254 a_6605_3239# D[0] 1.08e-20
C2255 a_9152_4775# a_10629_4801# 1.67e-19
C2256 VDD a_6466_4775# 0.488f
C2257 VDD a_4367_3213# 0.356f
C2258 check[1] a_9578_4112# 3.76e-20
C2259 x39.Q_N a_11856_3239# 0.162f
C2260 VDD reset 0.16f
C2261 x5.X a_8697_4112# 0.00599f
C2262 check[2] x42.Q_N 8.18e-19
C2263 sel_bit[0] x4.X 6.44e-20
C2264 x27.D a_4855_4775# 4.69e-21
C2265 a_7247_4775# a_7186_4112# 1.79e-20
C2266 check[5] a_6846_4086# 0.0346f
C2267 check[1] a_6759_3213# 2.39e-20
C2268 VDD a_7362_3239# 4.88e-19
C2269 D[0] a_8288_2340# 0.00665f
C2270 a_8236_3239# D[4] 5.41e-19
C2271 a_5896_2340# x57.Q_N 0.178f
C2272 a_6304_2366# a_6546_2340# 0.124f
C2273 a_5991_2340# a_6844_2640# 0.0264f
C2274 check[4] x39.Q_N 6.54e-19
C2275 a_8236_3239# x69.Q_N 1.07e-19
C2276 a_9151_3213# a_8997_3239# 0.00943f
C2277 a_8683_3605# a_8791_3239# 0.00812f
C2278 a_9464_3239# a_9322_3521# 0.00412f
C2279 a_8857_3213# a_9369_3239# 9.75e-19
C2280 a_9638_3213# a_9550_3605# 7.71e-20
C2281 VDD a_8939_4086# 0.34f
C2282 check[2] a_10680_2340# 0.027f
C2283 x5.X a_12737_3239# 0.00125f
C2284 a_9442_4086# a_9464_3239# 4.33e-20
C2285 a_9710_4296# a_9638_3213# 3.74e-20
C2286 x42.Q_N a_9151_3213# 0.0983f
C2287 x20.Q_N a_3912_2366# 1.17e-19
C2288 x4.X a_10156_4112# 0.00621f
C2289 a_11834_4086# a_12101_2550# 2.22e-22
C2290 x39.Q_N a_11629_2340# 3.65e-20
C2291 x30.Q_N x57.Q_N 4.08e-19
C2292 a_8697_4112# a_9237_4386# 0.139f
C2293 a_8384_4086# a_9238_4086# 0.0492f
C2294 x5.X a_4681_4801# 1.74e-19
C2295 check[6] a_3913_4112# 7.75e-22
C2296 x4.X a_8792_4801# 8.46e-20
C2297 a_1062_5674# a_897_4112# 9.53e-20
C2298 VDD D[2] 0.29f
C2299 check[3] x66.Q_N 0.00297f
C2300 a_4681_4801# a_4854_3213# 4.82e-21
C2301 a_4855_4775# a_4680_3239# 1.33e-23
C2302 VDD x60.Q_N 0.0716f
C2303 a_7317_2550# a_7561_2366# 0.00812f
C2304 x5.X a_11857_4801# 0.00141f
C2305 x33.Q_N comparator_out 0.263f
C2306 D[1] a_9754_3239# 8.74e-20
C2307 a_9152_4775# a_9639_4775# 0.273f
C2308 a_8858_4775# a_8591_4801# 6.99e-20
C2309 a_8403_4801# a_8768_5167# 4.45e-20
C2310 VDD a_3807_4801# 0.117f
C2311 x45.Q_N a_6465_3213# 0.194f
C2312 a_6846_4086# a_7246_3213# 7.94e-19
C2313 a_7050_4086# a_6759_3213# 0.0014f
C2314 a_5844_3239# a_6759_3213# 0.126f
C2315 comparator_out a_6291_3605# 0.00113f
C2316 a_9710_4296# a_9236_2640# 6.02e-22
C2317 a_9237_4386# a_9709_2550# 6.45e-21
C2318 x42.Q_N a_8938_2340# 0.00179f
C2319 x27.Q_N a_4018_2366# 0.0102f
C2320 x77.Y a_4925_2550# 0.00196f
C2321 x4.X check[6] 0.0328f
C2322 VDD a_10983_4801# 0.109f
C2323 a_10629_4801# a_10628_3239# 6.9e-19
C2324 x4.X check[3] 0.316f
C2325 a_8696_2366# a_9172_2366# 2.87e-21
C2326 x77.Y a_4585_3239# 0.00397f
C2327 check[1] a_1511_4112# 5.91e-22
C2328 a_6845_4386# a_6845_2340# 7.25e-19
C2329 a_5992_4086# x57.Q_N 2.32e-20
C2330 x45.Q_N a_5991_2340# 2.01e-19
C2331 a_6846_4086# a_6844_2640# 7.02e-19
C2332 comparator_out a_6304_2366# 0.00689f
C2333 sel_bit[1] a_2289_4801# 1.47e-20
C2334 a_11970_4112# a_12030_3213# 4.45e-20
C2335 check[5] a_8402_3239# 1.82e-19
C2336 check[2] a_9173_4112# 1.17e-20
C2337 x20.Q_N a_4113_4394# 6.16e-20
C2338 x5.X a_9375_4478# 7.3e-19
C2339 a_4074_4775# a_4539_5083# 9.46e-19
C2340 a_3619_4801# a_4767_5167# 2.13e-19
C2341 a_3453_4801# a_4214_4801# 6.04e-20
C2342 x5.X a_9102_5083# 3.46e-19
C2343 a_11834_4086# x39.Q_N 0.00118f
C2344 check[2] a_9873_5083# 4.31e-19
C2345 a_10775_2340# a_11288_2648# 0.00945f
C2346 a_2533_2550# D[6] 0.00108f
C2347 x4.X a_8896_2648# 0.00102f
C2348 a_7247_4775# a_7363_4801# 0.0397f
C2349 a_6760_4775# a_7182_4801# 2.87e-21
C2350 VDD a_8803_4112# 0.00996f
C2351 check[1] a_7318_4296# 0.0013f
C2352 x4.X a_11493_3521# 2.91e-19
C2353 check[1] comparator_out 0.134f
C2354 a_10795_4801# a_11943_5167# 2.13e-19
C2355 a_11250_4775# a_11715_5083# 9.46e-19
C2356 a_10629_4801# a_11390_4801# 6.04e-20
C2357 a_3452_3239# a_6010_3239# 2.9e-21
C2358 VDD a_9323_5083# 0.0163f
C2359 check[5] a_7185_2366# 4.92e-19
C2360 a_4453_4386# a_5992_4086# 1.24e-19
C2361 a_4658_4086# a_4593_4112# 9.75e-19
C2362 a_4454_4086# a_4794_4112# 6.04e-20
C2363 x33.Q_N a_8683_3605# 0.00192f
C2364 a_9237_4386# a_9375_4478# 1.09e-19
C2365 a_8939_4086# a_8803_4112# 0.0282f
C2366 a_8697_4112# a_9656_4394# 1.21e-20
C2367 x5.X a_897_4112# 0.00452f
C2368 VDD a_2198_2732# 0.0198f
C2369 a_5562_4801# a_5845_4801# 8.18e-19
C2370 check[6] a_3618_3239# 7.95e-22
C2371 a_8998_4801# a_8384_4086# 1.08e-19
C2372 a_4154_2340# a_4657_2340# 0.00187f
C2373 a_4452_2640# a_4453_2340# 0.781f
C2374 a_3912_2366# a_4925_2550# 0.0633f
C2375 a_6759_3213# a_8857_3213# 4.53e-20
C2376 a_7246_3213# a_8402_3239# 1.84e-19
C2377 a_7072_3239# a_8236_3239# 6.38e-20
C2378 a_3599_2340# x54.Q_N 0.124f
C2379 a_8237_4801# a_10346_4801# 1.03e-19
C2380 a_6759_3213# x72.Q_N 0.00553f
C2381 a_7246_3213# a_7480_3521# 0.00945f
C2382 a_6198_3239# a_6399_3239# 3.67e-19
C2383 a_7072_3239# a_6977_3239# 0.00276f
C2384 eob a_2463_4775# 0.00567f
C2385 x4.X a_6547_4086# 0.00727f
C2386 a_7050_4086# a_7318_4296# 0.205f
C2387 a_6846_4086# x45.Q_N 0.00113f
C2388 a_7050_4086# comparator_out 4.39e-21
C2389 x33.Q_N a_8696_2366# 0.0928f
C2390 a_5844_3239# comparator_out 0.147f
C2391 check[0] a_4872_4394# 8.58e-21
C2392 x5.X a_6978_4801# 2.58e-19
C2393 D[5] a_6546_2340# 2.03e-19
C2394 a_7246_3213# a_7185_2366# 1.2e-20
C2395 a_6011_4801# x30.Q_N 1.04e-19
C2396 a_7073_4801# a_7159_5167# 0.00976f
C2397 D[7] a_1207_2340# 0.00629f
C2398 a_1112_2340# a_1520_2366# 6.04e-19
C2399 a_4971_4801# a_4790_4801# 4.11e-20
C2400 check[2] a_2853_5648# 0.112f
C2401 a_2389_5648# check[1] 0.0168f
C2402 a_1511_4112# a_2061_2340# 0.00155f
C2403 x33.Q_N a_10795_4801# 2.19e-19
C2404 x20.Q_N D[6] 0.00261f
C2405 VDD a_7481_5083# 0.00506f
C2406 x33.Q_N a_11194_2366# 8.7e-20
C2407 x48.Q a_1976_4775# 4.67e-19
C2408 a_4855_4775# a_5562_4801# 0.0968f
C2409 a_4368_4775# check[6] 0.00421f
C2410 a_7561_2732# a_7763_2366# 8.94e-19
C2411 x39.Q_N a_12548_4112# 8.27e-20
C2412 check[1] a_8683_3605# 8.21e-20
C2413 a_11629_4386# a_12346_4112# 0.0019f
C2414 a_11834_4086# a_11769_4112# 9.75e-19
C2415 a_11630_4086# a_11970_4112# 6.04e-20
C2416 VDD a_11159_3605# 0.0042f
C2417 a_10628_3239# a_10794_3239# 0.782f
C2418 a_6304_2366# a_8696_2366# 5.35e-21
C2419 a_6845_2340# a_6984_2366# 2.56e-19
C2420 a_6844_2640# a_7185_2366# 0.00118f
C2421 a_6546_2340# a_8383_2340# 1.86e-21
C2422 x4.X a_1520_2366# 0.112f
C2423 check[5] a_9152_4775# 0.00306f
C2424 a_9872_3521# a_10628_3239# 4.06e-20
C2425 check[1] a_8289_4086# 0.125f
C2426 check[2] a_3671_5674# 0.00323f
C2427 a_1338_5674# a_1061_4801# 0.00179f
C2428 a_11544_4775# check[3] 0.00913f
C2429 a_12031_4775# a_12738_4801# 0.0968f
C2430 comparator_out a_2061_2340# 0.188f
C2431 x27.Q_N a_3599_2340# 0.142f
C2432 check[2] a_6846_4086# 2.36e-20
C2433 x77.Y a_6198_3239# 1.34e-20
C2434 x48.Q a_4155_4086# 0.00101f
C2435 a_6011_4801# a_5992_4086# 6.63e-19
C2436 a_5845_4801# a_6305_4112# 3.05e-19
C2437 check[3] a_12547_2366# 0.00323f
C2438 a_1976_4775# a_2147_5083# 0.00652f
C2439 VDD a_3258_5648# 0.116f
C2440 sel_bit[1] reset 1.45e-20
C2441 VDD a_12101_2550# 0.172f
C2442 check[1] a_8696_2366# 0.0033f
C2443 D[4] a_9172_2366# 3.13e-20
C2444 a_9237_2340# a_8896_2648# 1.25e-19
C2445 a_9236_2640# a_9172_2732# 2.13e-19
C2446 a_8938_2340# a_9374_2732# 0.00412f
C2447 a_8696_2366# a_8802_2366# 0.0552f
C2448 VDD sel_bit[1] 0.381f
C2449 x27.Q_N a_7073_4801# 7.65e-21
C2450 a_4214_4801# a_4790_4801# 2.46e-21
C2451 check[4] a_9238_4086# 0.0367f
C2452 a_9639_4775# a_9578_4112# 1.79e-20
C2453 x4.X a_4871_2648# 2.86e-19
C2454 VDD a_4794_4112# 0.0336f
C2455 a_9754_3239# a_9709_2550# 1.01e-20
C2456 x4.X a_6399_3239# 6.32e-19
C2457 check[1] a_3619_4801# 7.46e-20
C2458 a_9465_4801# x33.Q_N 8.55e-20
C2459 a_2853_5648# a_4074_4775# 1.12e-19
C2460 x45.Q_N a_8402_3239# 9.58e-19
C2461 comparator_out D[5] 0.00123f
C2462 comparator_out a_8857_3213# 4.83e-19
C2463 a_2853_5648# x20.Q_N 2.38e-20
C2464 x4.X a_6411_4112# 0.00336f
C2465 x45.Q_N a_7480_3521# 2.75e-19
C2466 comparator_out x72.Q_N 1.49e-19
C2467 a_6845_4386# a_6985_4112# 0.00126f
C2468 a_6547_4086# a_7186_4112# 0.00316f
C2469 a_7318_4296# a_7764_4112# 0.0367f
C2470 a_7764_4112# comparator_out 4.77e-20
C2471 a_9376_2366# a_9577_2366# 3.34e-19
C2472 a_10680_2340# a_11088_2366# 6.04e-19
C2473 check[6] a_7363_4801# 1.16e-20
C2474 a_2060_2640# a_2533_2550# 0.155f
C2475 a_2061_2340# a_2265_2340# 0.117f
C2476 a_1762_2340# x51.Q_N 9.58e-21
C2477 D[2] a_12101_2550# 2.21e-19
C2478 x45.Q_N a_7185_2366# 5.33e-22
C2479 check[4] a_9755_4801# 2.75e-19
C2480 comparator_out a_8383_2340# 0.00434f
C2481 a_1061_4801# a_3453_4801# 0.00176f
C2482 a_1338_5674# a_2389_5648# 0.00356f
C2483 a_1061_4801# a_2194_4801# 2.56e-19
C2484 a_1682_4775# a_1822_4801# 0.07f
C2485 a_1227_4801# a_1616_4801# 0.0019f
C2486 a_4454_4086# a_4926_4296# 0.15f
C2487 a_4453_4386# x48.Q_N 4.82e-21
C2488 check[0] a_6845_2340# 1.9e-19
C2489 a_3913_4112# x77.Y 3.94e-20
C2490 x5.X a_12102_4296# 1.62e-19
C2491 D[6] a_4925_2550# 6.65e-20
C2492 a_6010_3239# D[0] 5.69e-21
C2493 a_12101_2550# a_11969_2366# 0.0258f
C2494 VDD x39.Q_N 0.458f
C2495 comparator_out a_11766_2732# 9.47e-19
C2496 a_4073_3213# a_4018_2366# 5.71e-21
C2497 a_10776_4086# a_10628_3239# 8.29e-19
C2498 a_4680_3239# a_4789_3239# 0.00707f
C2499 x4.X x77.Y 0.07f
C2500 x33.Q_N D[4] 0.00278f
C2501 x5.X a_5561_3239# 0.00125f
C2502 VDD a_4388_2732# 0.00402f
C2503 sel_bit[0] a_2784_5996# 0.00164f
C2504 a_8939_4086# x39.Q_N 1.36e-20
C2505 x33.Q_N x69.Q_N 0.02f
C2506 a_2289_4801# x27.D 1.17e-20
C2507 check[0] a_3600_4086# 9e-20
C2508 a_4854_3213# a_5561_3239# 0.0968f
C2509 a_4367_3213# x75.Q 3.3e-19
C2510 VDD a_6930_3521# 0.0163f
C2511 check[6] a_6606_4801# 1.78e-19
C2512 check[6] x75.Q_N 0.00302f
C2513 a_8857_3213# a_8683_3605# 0.205f
C2514 a_8402_3239# a_9151_3213# 0.139f
C2515 a_8236_3239# a_9638_3213# 0.0492f
C2516 a_4453_2340# a_6546_2340# 6.38e-20
C2517 a_4925_2550# a_5991_2340# 7.98e-21
C2518 a_4657_2340# a_6304_2366# 1.32e-20
C2519 VDD a_6505_4394# 0.00506f
C2520 VDD x75.Q 0.216f
C2521 a_8998_4801# check[4] 1.23e-20
C2522 x39.Q_N D[2] 0.00168f
C2523 x20.Q_N a_2060_2640# 0.351f
C2524 a_6845_4386# a_7562_4112# 0.0019f
C2525 x4.X a_8858_4775# 9.41e-19
C2526 x5.X a_1415_4801# 0.00367f
C2527 x33.Q_N a_10775_2340# 1.5e-19
C2528 check[3] a_12030_3213# 0.00748f
C2529 a_6845_2340# a_7263_2648# 0.00276f
C2530 a_6844_2640# a_7561_2732# 4.45e-20
C2531 a_6304_2366# D[4] 1.86e-20
C2532 a_8857_3213# a_8696_2366# 0.0014f
C2533 a_8683_3605# a_8383_2340# 3.9e-20
C2534 a_8236_3239# a_9236_2640# 6.01e-20
C2535 a_7954_4801# check[5] 0.129f
C2536 a_11390_4801# a_10776_4086# 1.08e-19
C2537 a_6978_4801# x30.Q_N 1.41e-19
C2538 a_4155_4086# a_3599_2340# 1.3e-22
C2539 VDD a_1592_5167# 0.00558f
C2540 a_3913_4112# a_3912_2366# 1.8e-19
C2541 a_8384_4086# a_8288_2340# 2.97e-20
C2542 a_8289_4086# a_8383_2340# 1.57e-20
C2543 x33.Q_N a_11762_4801# 3.57e-20
C2544 check[1] a_6710_5083# 1.55e-19
C2545 x27.Q_N a_2979_2366# 1.34e-20
C2546 x27.Q_N a_6010_3239# 7.07e-20
C2547 x39.Q_N a_11969_2366# 5.33e-22
C2548 a_1062_5674# x5.X 0.00504f
C2549 x5.X a_4658_4086# 4.53e-19
C2550 check[6] a_5897_4086# 0.00265f
C2551 x48.Q a_4855_4775# 0.00105f
C2552 a_4658_4086# a_4854_3213# 2.47e-19
C2553 a_4926_4296# a_4367_3213# 1.71e-19
C2554 check[3] a_11628_2640# 0.0274f
C2555 check[1] D[4] 0.194f
C2556 x77.Y a_3618_3239# 0.528f
C2557 D[4] a_8802_2366# 5.38e-19
C2558 a_8383_2340# a_8696_2366# 0.273f
C2559 x4.X a_3912_2366# 0.105f
C2560 VDD x5.A 0.23f
C2561 a_10628_3239# a_11761_3239# 2.56e-19
C2562 a_11249_3213# a_11389_3239# 0.07f
C2563 a_11543_3213# a_11714_3521# 0.00652f
C2564 a_10794_3239# a_11183_3239# 0.0019f
C2565 VDD a_4926_4296# 0.319f
C2566 a_6846_4086# a_7953_3239# 4.72e-19
C2567 VDD a_11769_4112# 0.00445f
C2568 comparator_out a_4453_2340# 0.181f
C2569 x27.Q_N a_4793_2366# 0.0404f
C2570 check[5] a_6759_3213# 1.11e-19
C2571 a_7954_4801# a_7246_3213# 3.19e-20
C2572 x4.X a_6199_4801# 2.3e-19
C2573 x4.X a_4317_3521# 0.00111f
C2574 a_3453_4801# a_3619_4801# 0.75f
C2575 eob a_1996_2732# 4.16e-20
C2576 a_10681_4086# a_11629_4386# 7.74e-21
C2577 a_10156_4112# a_11630_4086# 3.65e-21
C2578 a_2463_4775# a_2398_4801# 4.2e-20
C2579 a_2289_4801# a_2579_4801# 0.0282f
C2580 a_2697_5083# a_3453_4801# 4.06e-20
C2581 check[2] a_9152_4775# 0.00242f
C2582 a_1207_2340# a_1720_2648# 0.00945f
C2583 a_1616_4801# x20.Q_N 4.31e-20
C2584 a_6011_4801# a_8237_4801# 4e-20
C2585 a_5845_4801# a_8403_4801# 2.9e-21
C2586 D[3] a_10680_2340# 0.0999f
C2587 x4.X a_6410_2366# 3.78e-20
C2588 check[0] a_3452_3239# 2.98e-21
C2589 a_11389_3239# a_10775_2340# 4.6e-20
C2590 x4.X a_8997_3239# 0.00265f
C2591 a_10629_4801# a_10795_4801# 0.751f
C2592 eob a_897_4112# 0.00374f
C2593 comparator_out a_7763_2366# 0.155f
C2594 comparator_out a_10794_3239# 0.148f
C2595 a_3913_4112# a_4113_4394# 0.00185f
C2596 a_3600_4086# a_4389_4478# 7.71e-20
C2597 x4.X x42.Q_N 0.252f
C2598 check[5] a_6546_2340# 1.34e-19
C2599 a_9152_4775# a_9151_3213# 0.00121f
C2600 x5.X a_3170_4801# 0.0367f
C2601 a_897_4112# x4.A 0.238f
C2602 a_8237_4801# a_8697_4112# 3.05e-19
C2603 a_8403_4801# a_8384_4086# 6.63e-19
C2604 check[0] a_6985_4112# 3.21e-20
C2605 sel_bit[0] a_2463_4775# 5.11e-20
C2606 a_3648_5972# a_3373_5674# 0.0156f
C2607 a_6759_3213# a_7246_3213# 0.273f
C2608 a_6465_3213# a_6198_3239# 6.99e-20
C2609 a_6010_3239# a_6375_3605# 4.45e-20
C2610 sel_bit[1] a_3258_5648# 0.259f
C2611 x4.X a_10680_2340# 0.00342f
C2612 check[3] a_11630_4086# 0.223f
C2613 VDD x27.D 0.294f
C2614 x4.X a_4113_4394# 1.78e-19
C2615 a_4073_3213# a_3599_2340# 2.5e-19
C2616 a_3618_3239# a_3912_2366# 5.94e-19
C2617 x33.Q_N a_6845_2340# 1.52e-19
C2618 x5.X a_6292_5167# 0.00462f
C2619 VDD a_2200_2366# 0.00214f
C2620 x3.A comparator_out 2e-20
C2621 a_3618_3239# a_4317_3521# 2.46e-19
C2622 a_3452_3239# a_4538_3521# 0.00907f
C2623 check[0] a_3900_5167# 8.76e-19
C2624 a_4367_3213# a_4680_3239# 0.124f
C2625 a_3899_3605# a_3806_3239# 0.0367f
C2626 a_4073_3213# a_3983_3605# 6.69e-20
C2627 a_6466_4775# a_6760_4775# 0.199f
C2628 a_6011_4801# a_7247_4775# 0.0264f
C2629 a_5845_4801# a_7073_4801# 0.0334f
C2630 a_4925_2550# a_5371_2366# 0.0367f
C2631 D[0] a_8236_3239# 0.348f
C2632 a_7953_3239# a_8402_3239# 3.93e-19
C2633 a_7072_3239# a_6304_2366# 2.17e-19
C2634 a_6198_3239# a_5991_2340# 2.02e-19
C2635 a_6759_3213# a_6844_2640# 5.32e-19
C2636 a_6977_3239# D[0] 1.36e-20
C2637 a_9465_4801# a_10629_4801# 6.38e-20
C2638 a_9639_4775# a_10795_4801# 1.25e-19
C2639 VDD a_6760_4775# 0.449f
C2640 check[2] a_10628_3239# 0.0451f
C2641 VDD a_4680_3239# 0.183f
C2642 x39.Q_N a_11159_3605# 8.48e-19
C2643 x5.X a_9237_4386# 0.00958f
C2644 x33.Q_N a_10155_2366# 0.032f
C2645 VDD a_6504_2648# 0.00506f
C2646 a_10776_4086# a_11289_4394# 0.00945f
C2647 x27.D a_3807_4801# 0.164f
C2648 check[5] comparator_out 0.0221f
C2649 VDD a_9101_3521# 0.00984f
C2650 a_6304_2366# a_6845_2340# 0.125f
C2651 a_6546_2340# a_6844_2640# 0.137f
C2652 a_9151_3213# a_10628_3239# 3.41e-19
C2653 a_9464_3239# a_8997_3239# 0.00316f
C2654 a_9151_3213# a_9369_3239# 3.73e-19
C2655 VDD a_9238_4086# 0.805f
C2656 x42.Q_N a_9464_3239# 0.162f
C2657 x4.X a_9173_4112# 8.4e-20
C2658 x39.Q_N a_12101_2550# 0.00196f
C2659 a_8939_4086# a_9238_4086# 0.0334f
C2660 a_8697_4112# a_9442_4086# 0.199f
C2661 a_8384_4086# a_9710_4296# 4.7e-22
C2662 a_7186_4112# x42.Q_N 4.05e-20
C2663 a_5562_4801# a_4454_4086# 6.67e-19
C2664 check[6] a_4453_4386# 0.0318f
C2665 a_10776_4086# comparator_out 0.00196f
C2666 a_4855_4775# a_7073_4801# 1.86e-21
C2667 a_4368_4775# a_6199_4801# 1.49e-21
C2668 check[0] a_7562_4112# 5.56e-22
C2669 check[1] a_6845_2340# 6.25e-19
C2670 x5.X a_11160_5167# 4.21e-19
C2671 D[4] a_8383_2340# 0.0132f
C2672 a_7763_2366# a_8696_2366# 3.42e-20
C2673 x4.X D[6] 0.00589f
C2674 x4.X a_6465_3213# 0.00499f
C2675 a_8237_4801# a_9102_5083# 0.00276f
C2676 a_9639_4775# a_9465_4801# 0.197f
C2677 a_8684_5167# a_8768_5167# 0.00972f
C2678 a_9152_4775# a_8591_4801# 2.47e-21
C2679 VDD a_2579_4801# 0.0073f
C2680 a_7050_4086# a_7072_3239# 4.33e-20
C2681 a_7318_4296# a_7246_3213# 3.74e-20
C2682 x45.Q_N a_6759_3213# 0.0983f
C2683 comparator_out a_7246_3213# 0.00381f
C2684 a_5844_3239# a_7072_3239# 0.0334f
C2685 x42.Q_N a_9237_2340# 3.65e-20
C2686 a_9442_4086# a_9709_2550# 2.22e-22
C2687 a_2883_5674# x48.Q 0.00144f
C2688 VDD a_9755_4801# 0.0101f
C2689 a_10795_4801# a_10794_3239# 1.39e-19
C2690 check[2] a_7954_4801# 4.53e-20
C2691 a_8696_2366# a_9577_2366# 0.00943f
C2692 a_9237_2340# a_10680_2340# 8.18e-19
C2693 a_8938_2340# a_9376_2366# 0.00276f
C2694 x77.Y x75.Q_N 3.94e-19
C2695 x4.X a_5991_2340# 0.111f
C2696 a_2853_5648# a_3913_4112# 4.72e-21
C2697 a_11389_3239# a_11965_3239# 2.46e-21
C2698 check[1] a_3600_4086# 1.19e-20
C2699 x45.Q_N a_6546_2340# 0.0018f
C2700 a_7318_4296# a_6844_2640# 6.02e-22
C2701 a_6845_4386# a_7317_2550# 6.45e-21
C2702 comparator_out a_6844_2640# 0.108f
C2703 a_5844_3239# a_6845_2340# 6.52e-20
C2704 x27.Q_N a_6984_2366# 2.64e-20
C2705 a_1511_4112# a_3505_4086# 0.0121f
C2706 x20.Q_N a_4591_4478# 6.94e-20
C2707 x5.X a_9656_4394# 2.97e-19
C2708 check[2] a_9578_4112# 1.87e-19
C2709 a_3619_4801# a_4008_4801# 0.0019f
C2710 a_4368_4775# a_4539_5083# 0.00652f
C2711 a_4074_4775# a_4214_4801# 0.07f
C2712 a_3453_4801# a_4586_4801# 2.56e-19
C2713 check[5] a_8289_4086# 0.00275f
C2714 x5.X a_9551_5167# 1.06e-19
C2715 a_1626_2366# a_1996_2366# 4.11e-20
C2716 x20.Q_N a_4214_4801# 1.27e-19
C2717 a_2853_5648# x4.X 5.73e-20
C2718 a_11088_2366# a_11564_2732# 0.00133f
C2719 x4.X a_9374_2732# 9.81e-19
C2720 a_7073_4801# a_7182_4801# 0.00707f
C2721 VDD a_9954_4478# 0.0042f
C2722 x4.X a_11942_3605# 4.4e-19
C2723 comparator_out a_9953_2732# 8.29e-19
C2724 a_1227_4801# a_1511_4112# 0.00301f
C2725 a_11544_4775# a_11715_5083# 0.00652f
C2726 a_10629_4801# a_11762_4801# 2.56e-19
C2727 x5.A sel_bit[1] 0.0425f
C2728 a_10795_4801# a_11184_4801# 0.0019f
C2729 a_11250_4775# a_11390_4801# 0.07f
C2730 VDD a_8998_4801# 0.0332f
C2731 a_5845_4801# a_6010_3239# 8.16e-19
C2732 a_4453_4386# a_6547_4086# 2.47e-20
C2733 a_4926_4296# a_4794_4112# 0.0258f
C2734 a_4454_4086# a_6305_4112# 5.07e-21
C2735 check[5] a_8696_2366# 2.42e-20
C2736 a_3505_4086# comparator_out 2.05e-21
C2737 a_9442_4086# a_9375_4478# 9.46e-19
C2738 x42.Q_N a_8897_4394# 2.02e-20
C2739 x33.Q_N a_9638_3213# 0.0126f
C2740 a_9639_4775# x69.Q_N 4.45e-20
C2741 a_8697_4112# a_10156_4112# 8.23e-22
C2742 a_9237_4386# a_9656_4394# 2.46e-19
C2743 VDD a_2479_2648# 0.0122f
C2744 check[6] a_6011_4801# 0.162f
C2745 a_7246_3213# a_8683_3605# 7.98e-21
C2746 a_6759_3213# a_9151_3213# 3.6e-20
C2747 a_4452_2640# a_4925_2550# 0.145f
C2748 a_4453_2340# a_4657_2340# 0.117f
C2749 a_4154_2340# x54.Q_N 9.58e-21
C2750 a_1061_4801# a_1227_4801# 0.619f
C2751 a_7072_3239# x72.Q_N 9.58e-21
C2752 a_8403_4801# check[4] 1.14e-20
C2753 eob a_1415_4801# 0.151f
C2754 VDD a_5562_4801# 0.192f
C2755 x4.X a_6846_4086# 0.0467f
C2756 VDD a_12738_4801# 0.177f
C2757 a_7318_4296# x45.Q_N 0.00243f
C2758 x45.Q_N comparator_out 0.00129f
C2759 x33.Q_N a_9236_2640# 0.572f
C2760 check[0] a_5372_4112# 0.165f
C2761 VDD a_4388_2366# 1.64e-19
C2762 x5.X x30.Q_N 8.83e-19
C2763 a_6292_5167# x30.Q_N 7.29e-20
C2764 a_6760_4775# a_7481_5083# 0.00185f
C2765 D[5] a_6845_2340# 1.11e-19
C2766 a_8236_3239# a_10345_3239# 1.03e-19
C2767 a_10629_4801# a_11089_4112# 3.05e-19
C2768 D[7] a_1762_2340# 8.38e-19
C2769 a_1112_2340# a_2060_2640# 7.7e-21
C2770 a_10795_4801# a_10776_4086# 6.63e-19
C2771 check[0] x27.Q_N 0.0367f
C2772 D[0] a_8791_3239# 1.27e-19
C2773 a_1062_5674# eob 2.23e-21
C2774 a_1511_4112# a_2533_2550# 6.53e-19
C2775 x33.Q_N a_11076_5167# 1.6e-19
C2776 check[2] a_1511_4112# 5.19e-20
C2777 sel_bit[1] x27.D 4.45e-19
C2778 a_1062_5674# x4.A 8.16e-22
C2779 check[2] a_11289_4394# 9.25e-20
C2780 x30.Q_N a_7181_3239# 1.68e-19
C2781 x48.Q a_2289_4801# 8.99e-20
C2782 check[3] a_12737_3239# 0.0275f
C2783 a_4681_4801# check[6] 4.98e-20
C2784 x39.Q_N a_11769_4112# 0.00167f
C2785 a_12102_4296# a_11970_4112# 0.0258f
C2786 check[5] a_9465_4801# 6.82e-20
C2787 a_6845_2340# a_8383_2340# 0.00116f
C2788 a_7049_2340# a_7185_2366# 0.07f
C2789 a_6844_2640# a_8696_2366# 1.79e-19
C2790 a_10628_3239# a_11075_3605# 0.15f
C2791 a_10794_3239# a_11249_3213# 0.153f
C2792 x4.X a_2060_2640# 0.00821f
C2793 check[1] a_6985_4112# 7.78e-20
C2794 x69.Q_N a_10794_3239# 8.64e-20
C2795 a_9872_3521# x69.Q_N 2.02e-20
C2796 a_2389_5648# a_1227_4801# 3.08e-19
C2797 x5.X a_3373_5674# 1.23e-19
C2798 a_11857_4801# check[3] 0.00257f
C2799 comparator_out a_2533_2550# 0.00698f
C2800 clk_sar a_1061_4801# 1.18e-19
C2801 x5.X a_5992_4086# 0.0202f
C2802 check[2] a_7318_4296# 2.18e-22
C2803 x27.Q_N a_4154_2340# 0.16f
C2804 x77.Y a_4970_3239# 0.00967f
C2805 a_4453_4386# a_6411_4112# 9.75e-21
C2806 check[2] comparator_out 0.125f
C2807 x48.Q a_4454_4086# 2.06e-19
C2808 a_6466_4775# a_6305_4112# 0.0025f
C2809 a_6292_5167# a_5992_4086# 4.9e-20
C2810 a_5845_4801# a_6845_4386# 9.86e-20
C2811 check[3] a_11768_2366# 9.26e-20
C2812 a_3452_3239# a_5844_3239# 0.00176f
C2813 a_1976_4775# a_1822_4801# 0.00943f
C2814 a_1508_5167# a_1616_4801# 0.00812f
C2815 a_2289_4801# a_2147_5083# 0.00412f
C2816 a_2463_4775# a_2375_5167# 7.71e-20
C2817 VDD a_3876_6040# 0.00865f
C2818 check[1] a_9236_2640# 3.18e-19
C2819 D[4] a_9577_2366# 7.47e-20
C2820 a_9237_2340# a_9374_2732# 0.00907f
C2821 x4.X a_5371_2366# 8.28e-20
C2822 VDD a_6305_4112# 0.448f
C2823 sel_bit[0] a_897_4112# 8.65e-21
C2824 a_10628_3239# a_11088_2366# 1.89e-19
C2825 a_10794_3239# a_10775_2340# 3.73e-19
C2826 x4.X a_8402_3239# 0.0429f
C2827 check[1] a_3900_5167# 4.17e-20
C2828 x4.X a_7480_3521# 0.00103f
C2829 eob a_3170_4801# 0.00132f
C2830 x4.X a_7562_4478# 9.15e-19
C2831 comparator_out a_9151_3213# 7.47e-19
C2832 a_7954_4801# a_7953_3239# 9.85e-20
C2833 a_3453_4801# a_3600_4086# 0.00159f
C2834 a_6845_4386# a_8384_4086# 2.16e-19
C2835 a_7050_4086# a_6985_4112# 9.75e-19
C2836 a_6846_4086# a_7186_4112# 6.04e-20
C2837 x45.Q_N a_8289_4086# 8.9e-21
C2838 x20.Q_N a_1511_4112# 0.0407f
C2839 eob a_1996_2366# 1.64e-21
C2840 a_6710_5083# check[5] 3.95e-22
C2841 a_10680_2340# a_11628_2640# 9.65e-21
C2842 a_2265_2340# a_2533_2550# 0.205f
C2843 a_2061_2340# x51.Q_N 1.07e-19
C2844 x5.X eob 0.155f
C2845 a_1227_4801# a_3619_4801# 7.69e-21
C2846 comparator_out a_8938_2340# 0.00103f
C2847 a_2389_5648# check[2] 0.138f
C2848 a_1682_4775# a_2194_4801# 9.75e-19
C2849 a_1061_4801# x20.Q_N 2.14e-19
C2850 check[5] D[4] 0.00424f
C2851 x5.X x4.A 6.17e-19
C2852 check[0] a_7317_2550# 1.78e-19
C2853 x33.Q_N D[0] 1.28e-20
C2854 a_4453_4386# x77.Y 1.11e-20
C2855 VDD a_1207_2340# 0.608f
C2856 x20.Q_N comparator_out 0.0881f
C2857 a_11565_4112# a_11970_4112# 2.46e-21
C2858 a_12548_4112# a_12346_4112# 3.67e-19
C2859 a_6291_3605# D[0] 3.23e-21
C2860 a_6759_3213# a_7953_3239# 6.04e-19
C2861 x4.X a_11564_2732# 4.32e-19
C2862 check[1] a_7562_4112# 1.69e-19
C2863 comparator_out a_12047_2648# 6.95e-19
C2864 a_10776_4086# a_11249_3213# 2.45e-19
C2865 a_11089_4112# a_10794_3239# 4.9e-19
C2866 check[2] a_8289_4086# 1.35e-21
C2867 x5.X a_6781_4478# 3.2e-19
C2868 sel_bit[0] a_3648_5972# 2.6e-19
C2869 x33.Q_N a_11543_3213# 8.28e-21
C2870 VDD a_4018_2366# 0.0028f
C2871 check[0] a_4155_4086# 4.34e-20
C2872 a_9238_4086# x39.Q_N 3.57e-19
C2873 VDD a_6605_3239# 5.47e-21
C2874 check[6] a_6978_4801# 6.18e-20
C2875 D[0] a_6304_2366# 1.92e-21
C2876 check[4] a_10681_4086# 0.00276f
C2877 a_3912_2366# x57.Q_N 8.28e-21
C2878 a_4453_2340# a_6845_2340# 0.00176f
C2879 a_8402_3239# a_9464_3239# 0.137f
C2880 a_8683_3605# a_9151_3213# 0.0633f
C2881 a_8236_3239# a_8590_3239# 0.0708f
C2882 VDD a_6983_4478# 0.0163f
C2883 VDD x48.Q 0.638f
C2884 a_9370_4801# check[4] 9.79e-21
C2885 check[2] a_8696_2366# 1.08e-21
C2886 a_8384_4086# a_8236_3239# 8.29e-19
C2887 a_10776_4086# a_10775_2340# 5.27e-19
C2888 x20.Q_N a_2265_2340# 0.194f
C2889 x30.Q_N a_5896_2340# 3.7e-19
C2890 check[2] a_3619_4801# 6.48e-20
C2891 x4.X a_9152_4775# 0.104f
C2892 a_2389_5648# x20.Q_N 2.12e-20
C2893 x5.X a_1926_5083# 3.49e-19
C2894 x33.Q_N a_11330_2340# 5.36e-20
C2895 a_3453_4801# a_3452_3239# 6.9e-19
C2896 check[1] D[0] 0.169f
C2897 VDD a_8288_2340# 0.189f
C2898 check[2] a_10795_4801# 0.00106f
C2899 a_8591_4801# comparator_out 1.94e-20
C2900 a_6845_2340# a_7763_2366# 0.0708f
C2901 a_7049_2340# a_7561_2732# 6.69e-20
C2902 a_6844_2640# D[4] 0.00557f
C2903 a_8857_3213# a_9236_2640# 2.68e-19
C2904 a_8236_3239# a_9441_2340# 4.77e-19
C2905 a_8402_3239# a_9237_2340# 6.38e-20
C2906 a_9151_3213# a_8696_2366# 3.36e-20
C2907 a_8683_3605# a_8938_2340# 2.41e-20
C2908 a_8997_3239# D[1] 1.13e-20
C2909 check[2] a_11194_2366# 0.00242f
C2910 VDD a_2147_5083# 0.0199f
C2911 a_4453_4386# a_3912_2366# 1.93e-22
C2912 x33.Q_N x36.Q_N 2.37e-20
C2913 check[1] a_7159_5167# 1.92e-19
C2914 x42.Q_N D[1] 0.00176f
C2915 x48.Q a_3807_4801# 0.00791f
C2916 a_4926_4296# a_4680_3239# 2.37e-20
C2917 a_3600_4086# a_4213_3239# 1.16e-20
C2918 check[3] a_11833_2340# 6.99e-20
C2919 x77.Y a_3899_3605# 0.181f
C2920 D[1] a_10680_2340# 0.00635f
C2921 a_10628_3239# D[3] 5.2e-19
C2922 a_8383_2340# a_9236_2640# 0.0264f
C2923 a_8696_2366# a_8938_2340# 0.124f
C2924 a_8288_2340# x60.Q_N 0.178f
C2925 x4.X a_4452_2640# 0.00799f
C2926 a_12030_3213# a_11942_3605# 7.71e-20
C2927 a_11249_3213# a_11761_3239# 9.75e-19
C2928 a_11856_3239# a_11714_3521# 0.00412f
C2929 a_11075_3605# a_11183_3239# 0.00812f
C2930 a_11543_3213# a_11389_3239# 0.00943f
C2931 a_10628_3239# x66.Q_N 1.07e-19
C2932 a_5897_4086# a_5991_2340# 1.57e-20
C2933 a_5992_4086# a_5896_2340# 2.97e-20
C2934 a_5844_3239# D[0] 7.04e-20
C2935 comparator_out a_7953_3239# 0.00109f
C2936 comparator_out a_4925_2550# 0.0087f
C2937 x27.Q_N a_6304_2366# 8.23e-20
C2938 x4.X a_4971_4801# 0.00557f
C2939 x4.X a_4766_3605# 6.48e-19
C2940 a_3619_4801# a_4074_4775# 0.153f
C2941 a_3453_4801# a_3900_5167# 0.15f
C2942 check[2] a_9465_4801# 0.00105f
C2943 x5.X a_8237_4801# 0.27f
C2944 x20.Q_N a_3619_4801# 4.85e-19
C2945 a_10776_4086# a_11089_4112# 0.272f
C2946 a_1520_2366# a_1996_2732# 0.00133f
C2947 a_2697_5083# x20.Q_N 2.02e-20
C2948 a_5088_3521# a_5844_3239# 4.06e-20
C2949 a_2853_5648# a_2784_5996# 0.00105f
C2950 check[0] a_5845_4801# 0.00285f
C2951 a_9709_2550# a_9953_2366# 0.00812f
C2952 x4.X a_7561_2732# 1.17e-19
C2953 x4.X a_10628_3239# 0.0456f
C2954 x4.X a_9369_3239# 4.91e-19
C2955 a_10795_4801# a_11250_4775# 0.153f
C2956 a_10629_4801# a_11076_5167# 0.15f
C2957 check[1] x27.Q_N 3.1e-20
C2958 VDD a_8403_4801# 0.593f
C2959 comparator_out a_11075_3605# 0.0011f
C2960 a_4155_4086# a_4389_4478# 0.00976f
C2961 a_3600_4086# a_4019_4112# 0.0397f
C2962 a_3913_4112# a_4591_4478# 0.00652f
C2963 check[5] a_6845_2340# 0.0379f
C2964 a_7764_4112# a_7562_4112# 3.67e-19
C2965 a_9639_4775# a_9638_3213# 0.00237f
C2966 a_2979_2366# a_2777_2366# 3.67e-19
C2967 a_8858_4775# a_8697_4112# 0.0025f
C2968 a_8684_5167# a_8384_4086# 4.9e-20
C2969 a_8237_4801# a_9237_4386# 9.86e-20
C2970 x36.Q_N a_11389_3239# 6.11e-19
C2971 a_3504_2340# a_3599_2340# 0.0968f
C2972 a_1996_2366# a_2401_2366# 2.46e-21
C2973 a_7246_3213# a_7072_3239# 0.197f
C2974 a_6291_3605# a_6375_3605# 0.00972f
C2975 a_6759_3213# a_6198_3239# 3.79e-20
C2976 a_2061_2340# x54.Q_N 2.94e-19
C2977 check[3] a_12102_4296# 0.00213f
C2978 a_2883_5674# a_2993_5674# 0.00857f
C2979 x4.X a_4591_4478# 0.00114f
C2980 comparator_out a_11088_2366# 0.00716f
C2981 a_5897_4086# a_6846_4086# 7e-20
C2982 a_4367_3213# a_3599_2340# 9.06e-19
C2983 a_4073_3213# a_4154_2340# 4.18e-20
C2984 a_3899_3605# a_3912_2366# 1.71e-19
C2985 a_3618_3239# a_4452_2640# 4.04e-20
C2986 a_3452_3239# a_4453_2340# 6.52e-20
C2987 x4.X a_4214_4801# 7.25e-19
C2988 x33.Q_N a_10345_3239# 0.0101f
C2989 x5.X a_7247_4775# 0.00983f
C2990 x27.Q_N a_5844_3239# 8.96e-20
C2991 check[6] a_5561_3239# 0.027f
C2992 x4.X a_11390_4801# 7.25e-19
C2993 VDD a_3599_2340# 0.58f
C2994 a_6466_4775# a_7073_4801# 0.00187f
C2995 a_6292_5167# a_7247_4775# 4.7e-22
C2996 a_1062_5674# sel_bit[0] 0.0419f
C2997 a_6011_4801# a_6199_4801# 0.162f
C2998 a_5845_4801# a_6376_5167# 0.0018f
C2999 a_3452_3239# a_4213_3239# 6.04e-20
C3000 a_3618_3239# a_4766_3605# 2.13e-19
C3001 a_4073_3213# a_4538_3521# 9.46e-19
C3002 check[0] a_4855_4775# 0.0127f
C3003 D[0] a_8857_3213# 8.87e-20
C3004 a_7072_3239# a_6844_2640# 1.11e-20
C3005 a_6759_3213# a_7049_2340# 0.00144f
C3006 a_7246_3213# a_6845_2340# 8.72e-19
C3007 x72.Q_N D[0] 2.5e-19
C3008 a_9639_4775# a_11076_5167# 7.98e-21
C3009 VDD a_3983_3605# 0.00494f
C3010 VDD a_7073_4801# 0.343f
C3011 check[2] x69.Q_N 4.68e-20
C3012 x4.X a_7954_4801# 0.00672f
C3013 x5.X a_9442_4086# 9.38e-19
C3014 VDD a_6982_2732# 0.0163f
C3015 a_11089_4112# a_11565_4478# 0.00133f
C3016 eob a_3373_5674# 1.33e-19
C3017 VDD a_9550_3605# 0.00371f
C3018 D[0] a_8383_2340# 0.00127f
C3019 a_6304_2366# a_7317_2550# 0.0633f
C3020 a_6844_2640# a_6845_2340# 0.781f
C3021 a_5991_2340# x57.Q_N 0.124f
C3022 a_6546_2340# a_7049_2340# 0.00187f
C3023 a_9464_3239# a_10628_3239# 6.38e-20
C3024 a_9638_3213# a_10794_3239# 1.69e-19
C3025 a_9151_3213# a_11249_3213# 4.53e-20
C3026 a_9464_3239# a_9369_3239# 0.00276f
C3027 a_8590_3239# a_8791_3239# 3.67e-19
C3028 a_9638_3213# a_9872_3521# 0.00945f
C3029 VDD a_9710_4296# 0.317f
C3030 a_9151_3213# x69.Q_N 0.00553f
C3031 check[2] a_10775_2340# 0.0128f
C3032 x27.Q_N a_2061_2340# 1.55e-19
C3033 x42.Q_N a_8767_3605# 8.48e-19
C3034 x4.X a_9578_4112# 0.0031f
C3035 check[4] a_8236_3239# 1.94e-20
C3036 a_9237_4386# a_9442_4086# 0.153f
C3037 a_8697_4112# x42.Q_N 0.0927f
C3038 a_4368_4775# a_4971_4801# 0.0552f
C3039 x5.X a_9574_4801# 5.36e-20
C3040 D[4] a_8938_2340# 1.94e-19
C3041 a_9638_3213# a_9577_2366# 1.2e-20
C3042 x4.X a_6759_3213# 0.111f
C3043 a_8403_4801# a_9323_5083# 1.09e-19
C3044 a_8858_4775# a_9102_5083# 0.0104f
C3045 VDD a_4318_5083# 0.0104f
C3046 a_2853_5648# a_2463_4775# 9.54e-20
C3047 x45.Q_N a_7072_3239# 0.162f
C3048 x48.Q a_3258_5648# 0.00631f
C3049 comparator_out a_6198_3239# 0.158f
C3050 a_5844_3239# a_6375_3605# 0.0018f
C3051 sel_bit[1] x48.Q 0.173f
C3052 a_6305_4112# a_6505_4394# 0.00185f
C3053 a_5992_4086# a_6781_4478# 7.71e-20
C3054 x42.Q_N a_9709_2550# 0.00196f
C3055 x27.Q_N D[5] 0.00536f
C3056 VDD a_11494_5083# 0.00984f
C3057 a_1508_5167# a_1511_4112# 3.47e-19
C3058 a_11250_4775# a_11249_3213# 2.59e-19
C3059 a_10795_4801# a_11075_3605# 8.52e-21
C3060 a_11076_5167# a_10794_3239# 1.65e-21
C3061 a_11544_4775# a_10628_3239# 9.66e-21
C3062 sel_bit[0] x5.X 0.0739f
C3063 a_9953_2732# a_10155_2366# 8.94e-19
C3064 a_8696_2366# a_11088_2366# 4.59e-21
C3065 a_9237_2340# a_9376_2366# 2.56e-19
C3066 a_8938_2340# a_10775_2340# 1.86e-21
C3067 a_9236_2640# a_9577_2366# 0.00118f
C3068 a_12146_3239# a_11965_3239# 4.11e-20
C3069 x4.X a_6546_2340# 0.00704f
C3070 eob x4.A 0.0197f
C3071 x45.Q_N a_6845_2340# 3.65e-20
C3072 a_7050_4086# a_7317_2550# 2.22e-22
C3073 comparator_out a_7049_2340# 0.00589f
C3074 a_1061_4801# a_1508_5167# 0.138f
C3075 a_3505_4086# a_3600_4086# 0.0968f
C3076 a_1511_4112# a_3913_4112# 1e-19
C3077 x5.X a_10156_4112# 9.37e-19
C3078 check[2] a_11089_4112# 0.00131f
C3079 a_4855_4775# a_4767_5167# 7.71e-20
C3080 a_4074_4775# a_4586_4801# 9.75e-19
C3081 a_4681_4801# a_4539_5083# 0.00412f
C3082 a_3900_5167# a_4008_4801# 0.00812f
C3083 a_4368_4775# a_4214_4801# 0.00943f
C3084 a_3453_4801# x27.Q_N 2.36e-19
C3085 x5.X a_8792_4801# 2.86e-19
C3086 x20.Q_N a_4586_4801# 5.69e-20
C3087 a_11088_2366# a_11194_2366# 0.0552f
C3088 a_11330_2340# a_11766_2732# 0.00412f
C3089 a_11628_2640# a_11564_2732# 2.13e-19
C3090 a_11629_2340# a_11288_2648# 1.25e-19
C3091 x4.X a_9655_2648# 2.86e-19
C3092 x30.Q_N a_8237_4801# 3.15e-19
C3093 x4.X a_11183_3239# 6.32e-19
C3094 VDD a_10681_4086# 0.189f
C3095 x4.X a_1511_4112# 1.74f
C3096 a_12031_4775# a_11943_5167# 7.71e-20
C3097 a_11857_4801# a_11715_5083# 0.00412f
C3098 a_10629_4801# x36.Q_N 1.22e-19
C3099 comparator_out D[3] 0.00125f
C3100 a_11250_4775# a_11762_4801# 9.75e-19
C3101 a_11076_5167# a_11184_4801# 0.00812f
C3102 a_11544_4775# a_11390_4801# 0.00943f
C3103 comparator_out a_1112_2340# 1.42e-19
C3104 a_6011_4801# a_6465_3213# 3.18e-21
C3105 a_4367_3213# a_6010_3239# 2.89e-19
C3106 VDD a_9370_4801# 0.00445f
C3107 x4.X a_11289_4394# 1.75e-19
C3108 comparator_out x66.Q_N 2.08e-20
C3109 a_4453_4386# a_6846_4086# 2.9e-21
C3110 a_3913_4112# comparator_out 2.29e-20
C3111 x5.X check[6] 0.168f
C3112 a_9237_4386# a_10156_4112# 0.162f
C3113 a_9442_4086# a_9656_4394# 0.0104f
C3114 a_8697_4112# a_9173_4112# 2.87e-21
C3115 a_9238_4086# a_9954_4478# 0.0018f
C3116 VDD a_2979_2366# 0.117f
C3117 VDD a_6010_3239# 0.274f
C3118 check[6] a_4854_3213# 0.00397f
C3119 check[6] a_6292_5167# 0.00105f
C3120 x5.X check[3] 0.285f
C3121 a_4453_2340# x54.Q_N 1.07e-19
C3122 a_4657_2340# a_4925_2550# 0.205f
C3123 a_1061_4801# x4.X 0.0131f
C3124 a_8684_5167# check[4] 4.29e-21
C3125 a_9152_4775# a_10346_4801# 6.04e-19
C3126 a_1227_4801# a_1682_4775# 0.145f
C3127 eob a_1926_5083# 0.00171f
C3128 check[6] a_5169_2366# 5.24e-20
C3129 x4.X a_7318_4296# 0.0211f
C3130 x4.X comparator_out 0.797f
C3131 x33.Q_N a_9441_2340# 0.179f
C3132 check[0] a_4389_4112# 8.48e-21
C3133 VDD a_4793_2366# 9.91e-19
C3134 a_7953_3239# D[4] 0.00127f
C3135 a_10629_4801# a_11629_4386# 9.86e-20
C3136 a_11250_4775# a_11089_4112# 0.0025f
C3137 a_11076_5167# a_10776_4086# 4.9e-20
C3138 a_8402_3239# D[1] 5.69e-21
C3139 D[5] a_7317_2550# 1.96e-20
C3140 a_7247_4775# x30.Q_N 0.126f
C3141 D[7] a_2061_2340# 1.85e-19
C3142 check[1] a_5845_4801# 5.4e-19
C3143 check[2] a_3600_4086# 1.65e-20
C3144 a_3505_4086# a_3452_3239# 5.06e-19
C3145 check[2] a_11767_4478# 5.02e-20
C3146 x33.Q_N a_11564_2366# 1e-20
C3147 VDD a_9172_2732# 0.00371f
C3148 x39.Q_N a_12346_4112# 2.43e-19
C3149 VDD a_11714_3521# 0.0163f
C3150 check[1] a_8590_3239# 0.00666f
C3151 x4.X a_2265_2340# 0.00118f
C3152 a_6845_2340# a_8938_2340# 6.38e-20
C3153 a_7317_2550# a_8383_2340# 7.98e-21
C3154 a_7049_2340# a_8696_2366# 8.4e-21
C3155 a_10628_3239# a_12030_3213# 0.0492f
C3156 a_10794_3239# a_11543_3213# 0.139f
C3157 a_11249_3213# a_11075_3605# 0.205f
C3158 check[1] a_8384_4086# 0.0126f
C3159 a_2389_5648# x4.X 0.00219f
C3160 a_11160_5167# check[3] 1.13e-19
C3161 x42.Q_N a_10982_3239# 1.34e-20
C3162 a_9442_4086# a_9754_3239# 5.48e-21
C3163 x27.Q_N a_4453_2340# 0.0462f
C3164 x5.X a_6547_4086# 0.00115f
C3165 x48.Q a_4926_4296# 1.36e-19
C3166 a_1976_4775# a_3453_4801# 1.75e-19
C3167 a_6466_4775# a_6845_4386# 3.92e-19
C3168 a_6292_5167# a_6547_4086# 2.46e-20
C3169 a_6760_4775# a_6305_4112# 5.67e-20
C3170 a_6011_4801# a_6846_4086# 1.18e-19
C3171 a_5845_4801# a_7050_4086# 6.96e-19
C3172 a_5845_4801# a_5844_3239# 6.9e-19
C3173 check[3] a_12345_2366# 5.09e-20
C3174 a_3618_3239# comparator_out 4.91e-19
C3175 a_1976_4775# a_2194_4801# 3.73e-19
C3176 a_2289_4801# a_1822_4801# 0.00316f
C3177 VDD a_2993_5674# 4.34e-19
C3178 x77.Y a_5561_3239# 3.29e-19
C3179 check[1] a_9441_2340# 4.56e-19
C3180 x27.Q_N a_4790_4801# 8.36e-20
C3181 x27.Q_N a_4213_3239# 6.11e-19
C3182 a_9237_2340# a_9655_2648# 0.00276f
C3183 a_9236_2640# a_9953_2732# 4.45e-20
C3184 a_8696_2366# D[3] 1.61e-20
C3185 VDD a_6845_4386# 0.59f
C3186 a_11249_3213# a_11088_2366# 0.0014f
C3187 a_11075_3605# a_10775_2340# 3.9e-20
C3188 a_10628_3239# a_11628_2640# 6.01e-20
C3189 x4.X a_8683_3605# 0.0177f
C3190 check[1] a_4855_4775# 1.73e-19
C3191 x4.X a_8289_4086# 0.00368f
C3192 comparator_out a_9464_3239# 1.93e-19
C3193 a_5844_3239# a_8590_3239# 3.65e-21
C3194 check[5] D[0] 0.417f
C3195 check[4] a_9172_2366# 2.2e-20
C3196 a_3619_4801# a_3913_4112# 9.06e-19
C3197 a_4074_4775# a_3600_4086# 4.54e-19
C3198 a_6845_4386# a_8939_4086# 3.16e-20
C3199 a_6846_4086# a_8697_4112# 5.07e-21
C3200 a_7318_4296# a_7186_4112# 0.0258f
C3201 x45.Q_N a_6985_4112# 0.00166f
C3202 a_7363_4801# a_6759_3213# 1.05e-20
C3203 x20.Q_N a_3600_4086# 0.00304f
C3204 x36.Q_N a_10794_3239# 3.85e-19
C3205 a_1520_2366# a_1996_2366# 2.87e-21
C3206 D[3] a_11194_2366# 5.39e-19
C3207 a_10775_2340# a_11088_2366# 0.273f
C3208 x4.X a_8696_2366# 0.112f
C3209 comparator_out a_9237_2340# 0.184f
C3210 x4.X a_3619_4801# 0.00737f
C3211 a_1682_4775# x20.Q_N 1.32e-19
C3212 a_9639_4775# a_10345_3239# 4.94e-20
C3213 x27.Q_N a_4019_4112# 2.89e-22
C3214 x4.X a_10795_4801# 0.00496f
C3215 a_4658_4086# x77.Y 1.87e-21
C3216 x48.Q x27.D 0.0333f
C3217 VDD a_1762_2340# 0.201f
C3218 a_4008_4801# x27.Q_N 4.32e-20
C3219 a_3912_2366# a_4112_2648# 0.00185f
C3220 a_3599_2340# a_4388_2732# 7.71e-20
C3221 a_7246_3213# D[0] 0.0116f
C3222 x4.X a_11194_2366# 3.78e-20
C3223 a_4970_3239# a_4452_2640# 5.05e-21
C3224 check[2] a_9638_3213# 0.0022f
C3225 check[6] a_5896_2340# 0.00282f
C3226 comparator_out a_12547_2366# 0.155f
C3227 a_11629_4386# a_10794_3239# 4.11e-20
C3228 a_10776_4086# a_11543_3213# 8.83e-19
C3229 a_11331_4086# a_11249_3213# 1.02e-19
C3230 a_11630_4086# a_10628_3239# 6.54e-20
C3231 a_11089_4112# a_11075_3605# 1.61e-19
C3232 a_6606_4801# a_6759_3213# 1.61e-20
C3233 x75.Q_N a_6759_3213# 2.97e-20
C3234 sel_bit[0] a_3373_5674# 0.0563f
C3235 VDD a_5169_2732# 0.00436f
C3236 a_2147_5083# x27.D 2.85e-21
C3237 VDD a_8236_3239# 0.791f
C3238 a_9710_4296# x39.Q_N 1.29e-19
C3239 check[0] a_4454_4086# 0.44f
C3240 VDD a_6977_3239# 6.2e-19
C3241 check[6] x30.Q_N 1.48e-21
C3242 D[0] a_6844_2640# 6.76e-19
C3243 a_7953_3239# a_6845_2340# 4.83e-19
C3244 a_9151_3213# a_9638_3213# 0.273f
C3245 a_8857_3213# a_8590_3239# 6.99e-20
C3246 a_8402_3239# a_8767_3605# 4.45e-20
C3247 a_4452_2640# x57.Q_N 1.53e-19
C3248 VDD a_7264_4394# 0.00984f
C3249 x33.Q_N check[4] 0.842f
C3250 eob a_2398_4801# 2.92e-19
C3251 check[2] a_9236_2640# 8.03e-20
C3252 a_8384_4086# a_8857_3213# 2.45e-19
C3253 a_8697_4112# a_8402_3239# 4.9e-19
C3254 a_11331_4086# a_10775_2340# 1.3e-22
C3255 a_11089_4112# a_11088_2366# 1.8e-19
C3256 x20.Q_N x51.Q_N 4.6e-19
C3257 a_7764_4112# a_8384_4086# 8.26e-21
C3258 x45.Q_N a_7562_4112# 2.38e-19
C3259 check[2] a_3900_5167# 5.02e-20
C3260 a_6845_4386# a_8803_4112# 3.66e-20
C3261 x4.X a_9465_4801# 0.00321f
C3262 x33.Q_N a_11629_2340# 7.03e-21
C3263 x5.X a_2375_5167# 1.58e-19
C3264 a_3453_4801# a_5845_4801# 0.00176f
C3265 a_3619_4801# a_3618_3239# 1.39e-19
C3266 VDD a_6984_2366# 6.2e-19
C3267 a_7363_4801# a_7318_4296# 1.9e-20
C3268 x20.Q_N a_3452_3239# 0.00411f
C3269 a_3170_4801# x77.Y 5.69e-20
C3270 a_10345_3239# a_10794_3239# 3.74e-19
C3271 D[1] a_10628_3239# 0.348f
C3272 a_7317_2550# a_7763_2366# 0.0367f
C3273 a_9464_3239# a_8696_2366# 2.17e-19
C3274 a_8590_3239# a_8383_2340# 2.02e-19
C3275 a_9151_3213# a_9236_2640# 5.32e-19
C3276 a_9369_3239# D[1] 1.36e-20
C3277 a_4454_4086# a_4154_2340# 3.47e-21
C3278 a_4453_4386# a_4452_2640# 1.32e-20
C3279 a_4658_4086# a_3912_2366# 7.14e-22
C3280 VDD a_1822_4801# 0.00544f
C3281 a_8384_4086# a_8383_2340# 5.27e-19
C3282 sel_bit[0] eob 0.294f
C3283 check[6] a_5992_4086# 0.00385f
C3284 x48.Q a_2579_4801# 1.65e-19
C3285 VDD a_11288_2648# 0.00506f
C3286 a_4971_4801# a_4453_4386# 8.84e-21
C3287 sel_bit[0] x4.A 1.17e-20
C3288 x77.Y a_4854_3213# 0.142f
C3289 x4.X a_4657_2340# 0.0013f
C3290 a_8696_2366# a_9237_2340# 0.125f
C3291 a_8938_2340# a_9236_2640# 0.137f
C3292 a_11543_3213# a_12146_3239# 0.0552f
C3293 a_11856_3239# a_11389_3239# 0.00316f
C3294 a_11543_3213# a_11761_3239# 3.73e-19
C3295 x45.Q_N D[0] 0.00168f
C3296 reset a_621_4112# 0.197f
C3297 a_11195_4112# a_11249_3213# 3.34e-20
C3298 x27.Q_N a_6844_2640# 1.07e-20
C3299 VDD a_621_4112# 0.255f
C3300 check[4] a_8802_2366# 1.3e-19
C3301 x4.X a_4007_3239# 6.32e-19
C3302 a_4074_4775# a_3900_5167# 0.205f
C3303 a_3619_4801# a_4368_4775# 0.139f
C3304 a_3453_4801# a_4855_4775# 0.0492f
C3305 x30.Q_N a_6547_4086# 1.3e-22
C3306 a_10776_4086# a_11629_4386# 0.0264f
C3307 a_11089_4112# a_11331_4086# 0.124f
C3308 x5.X a_8858_4775# 0.00316f
C3309 x20.Q_N a_3900_5167# 2.13e-19
C3310 a_10681_4086# x39.Q_N 0.181f
C3311 x75.Q_N comparator_out 1.48e-19
C3312 a_2853_5648# a_3648_5972# 0.00271f
C3313 a_1520_2366# a_1626_2366# 0.0552f
C3314 a_1762_2340# a_2198_2732# 0.00412f
C3315 a_2060_2640# a_1996_2732# 2.13e-19
C3316 a_2061_2340# a_1720_2648# 1.25e-19
C3317 a_6760_4775# a_8403_4801# 1.55e-19
C3318 a_7247_4775# a_8237_4801# 0.00116f
C3319 check[1] a_2883_5674# 0.195f
C3320 a_2853_5648# a_2969_6040# 0.00149f
C3321 x4.X D[4] 5.2e-19
C3322 a_10155_2366# a_11088_2366# 3.42e-20
C3323 D[3] a_10775_2340# 0.0131f
C3324 check[0] a_4367_3213# 2.58e-20
C3325 x4.X a_11249_3213# 0.00509f
C3326 x4.X x69.Q_N 0.00454f
C3327 a_10629_4801# a_12031_4775# 0.0492f
C3328 a_10795_4801# a_11544_4775# 0.139f
C3329 a_11250_4775# a_11076_5167# 0.205f
C3330 comparator_out a_12030_3213# 0.00336f
C3331 VDD a_8684_5167# 0.317f
C3332 VDD check[0] 0.685f
C3333 a_4155_4086# a_4019_4112# 0.0282f
C3334 a_3913_4112# a_4872_4394# 1.21e-20
C3335 a_4453_4386# a_4591_4478# 1.09e-19
C3336 check[5] a_7317_2550# 0.00103f
C3337 x36.Q_N a_12146_3239# 0.00341f
C3338 x36.Q_N a_11761_3239# 4.03e-19
C3339 a_8684_5167# a_8939_4086# 2.46e-20
C3340 a_9152_4775# a_8697_4112# 5.67e-20
C3341 a_8403_4801# a_9238_4086# 1.18e-19
C3342 a_8237_4801# a_9442_4086# 6.96e-19
C3343 a_8858_4775# a_9237_4386# 3.92e-19
C3344 a_6465_3213# a_6709_3521# 0.0104f
C3345 a_6010_3239# a_6930_3521# 1.09e-19
C3346 x4.X a_10775_2340# 0.11f
C3347 sel_bit[1] a_2993_5674# 4.44e-19
C3348 x4.X a_4872_4394# 8.47e-19
C3349 x75.Q a_6010_3239# 0.00207f
C3350 a_4854_3213# a_3912_2366# 8.4e-19
C3351 a_4073_3213# a_4453_2340# 0.00199f
C3352 a_4367_3213# a_4154_2340# 2.17e-19
C3353 comparator_out a_11628_2640# 0.108f
C3354 a_3618_3239# a_4657_2340# 0.00154f
C3355 a_5992_4086# a_6547_4086# 0.197f
C3356 a_5372_4112# x45.Q_N 8.9e-20
C3357 a_5897_4086# comparator_out 2.05e-21
C3358 x4.X a_4586_4801# 5.55e-19
C3359 x27.Q_N x45.Q_N 2.8e-20
C3360 x5.X a_6199_4801# 0.00541f
C3361 VDD a_4154_2340# 0.182f
C3362 x4.X a_11762_4801# 5.55e-19
C3363 a_3452_3239# a_4585_3239# 2.56e-19
C3364 a_3618_3239# a_4007_3239# 0.0019f
C3365 a_6760_4775# a_7073_4801# 0.124f
C3366 a_4073_3213# a_4213_3239# 0.07f
C3367 a_4367_3213# a_4538_3521# 0.00652f
C3368 a_6011_4801# a_4971_4801# 1.71e-20
C3369 a_6466_4775# a_6376_5167# 6.69e-20
C3370 a_6292_5167# a_6199_4801# 0.0367f
C3371 a_4018_2366# a_4388_2366# 4.11e-20
C3372 sel_bit[0] x48.Q_N 3.83e-20
C3373 D[0] a_9151_3213# 1.24e-19
C3374 a_7246_3213# a_7317_2550# 1.66e-21
C3375 a_7072_3239# a_7049_2340# 1.03e-19
C3376 check[2] a_11543_3213# 1.77e-20
C3377 VDD a_6376_5167# 0.0042f
C3378 VDD a_4538_3521# 0.0174f
C3379 x39.Q_N a_11714_3521# 0.00203f
C3380 x30.Q_N a_6399_3239# 6.75e-20
C3381 x5.X x42.Q_N 0.00729f
C3382 VDD a_7263_2648# 0.00984f
C3383 x30.Q_N a_6411_4112# 2.89e-22
C3384 x27.D a_4318_5083# 3.45e-21
C3385 a_11089_4112# a_11195_4112# 0.051f
C3386 a_11331_4086# a_11767_4478# 0.00412f
C3387 a_11629_4386# a_11565_4478# 2.13e-19
C3388 a_11630_4086# a_11289_4394# 1.25e-19
C3389 eob a_2788_5674# 1.71e-19
C3390 a_9638_3213# a_11075_3605# 7.98e-21
C3391 a_9151_3213# a_11543_3213# 3.6e-20
C3392 a_6844_2640# a_7317_2550# 0.145f
C3393 a_6845_2340# a_7049_2340# 0.117f
C3394 a_6546_2340# x57.Q_N 9.58e-21
C3395 a_9464_3239# x69.Q_N 9.58e-21
C3396 check[2] a_11330_2340# 0.00111f
C3397 a_2389_5648# a_2784_5996# 0.0102f
C3398 x20.Q_N x54.Q_N 1.47e-19
C3399 x4.X a_11089_4112# 0.109f
C3400 x30.Q_N a_6780_2366# 9.42e-19
C3401 a_4019_4112# a_4073_3213# 3.34e-20
C3402 check[2] x27.Q_N 3.57e-20
C3403 a_9237_4386# x42.Q_N 0.00118f
C3404 a_9238_4086# a_9710_4296# 0.15f
C3405 a_11630_4086# comparator_out 3e-20
C3406 a_4855_4775# a_4790_4801# 4.2e-20
C3407 a_4681_4801# a_4971_4801# 0.0282f
C3408 a_10628_3239# a_12737_3239# 1.03e-19
C3409 VDD a_4389_4478# 0.00402f
C3410 x5.X a_11715_5083# 6.65e-19
C3411 check[2] x36.Q_N 0.0011f
C3412 D[4] a_9237_2340# 1.09e-19
C3413 D[1] a_11183_3239# 1.22e-19
C3414 x4.X a_7072_3239# 0.00457f
C3415 a_8591_4801# a_8768_5167# 8.94e-19
C3416 a_8403_4801# a_8998_4801# 0.00118f
C3417 a_9152_4775# a_9102_5083# 1.21e-20
C3418 VDD a_4767_5167# 0.00394f
C3419 x45.Q_N a_6375_3605# 8.49e-19
C3420 a_11390_4801# a_11966_4801# 2.46e-21
C3421 a_6305_4112# a_6983_4478# 0.00652f
C3422 a_5992_4086# a_6411_4112# 0.0397f
C3423 a_6547_4086# a_6781_4478# 0.00976f
C3424 VDD a_11943_5167# 0.00371f
C3425 a_2463_4775# a_1511_4112# 0.0111f
C3426 check[4] a_8383_2340# 2.57e-20
C3427 a_11250_4775# a_11543_3213# 7.57e-21
C3428 a_10629_4801# a_11856_3239# 4.76e-21
C3429 eob a_1520_2366# 1.2e-19
C3430 a_5845_4801# check[5] 8.72e-20
C3431 a_6011_4801# a_7954_4801# 8.38e-21
C3432 a_9755_4801# a_9710_4296# 1.9e-20
C3433 a_9236_2640# a_11088_2366# 1.89e-19
C3434 a_9441_2340# a_9577_2366# 0.07f
C3435 a_9237_2340# a_10775_2340# 0.00116f
C3436 x4.X a_6845_2340# 0.00277f
C3437 check[1] a_4454_4086# 2.15e-20
C3438 a_10346_4801# a_10795_4801# 3.41e-19
C3439 check[4] a_10629_4801# 0.413f
C3440 x4.A a_1520_2366# 6.86e-19
C3441 a_12264_3521# x66.Q_N 2.02e-20
C3442 x45.Q_N a_7317_2550# 0.00196f
C3443 comparator_out D[1] 0.025f
C3444 comparator_out x57.Q_N 2.04e-19
C3445 a_1061_4801# a_2463_4775# 0.0492f
C3446 a_1682_4775# a_1508_5167# 0.205f
C3447 a_1227_4801# a_1976_4775# 0.132f
C3448 a_3600_4086# a_3913_4112# 0.273f
C3449 check[2] a_11629_4386# 1.44e-19
C3450 a_4681_4801# a_4214_4801# 0.00316f
C3451 a_4368_4775# a_4586_4801# 3.73e-19
C3452 a_4074_4775# x27.Q_N 1.34e-19
C3453 check[5] a_8384_4086# 0.0042f
C3454 D[6] a_1996_2366# 3.71e-20
C3455 x20.Q_N x27.Q_N 1.21e-20
C3456 a_11629_2340# a_11766_2732# 0.00907f
C3457 x4.X a_10155_2366# 7.73e-20
C3458 x4.X a_11965_3239# 1.05e-19
C3459 x4.X a_12264_3521# 0.00103f
C3460 VDD a_9377_4112# 0.00445f
C3461 x4.X a_3600_4086# 0.106f
C3462 a_11250_4775# x36.Q_N 2.08e-20
C3463 a_11857_4801# a_11390_4801# 0.00316f
C3464 a_11544_4775# a_11762_4801# 3.73e-19
C3465 a_6292_5167# a_6465_3213# 3.52e-21
C3466 a_6466_4775# a_6291_3605# 1.33e-23
C3467 a_6011_4801# a_6759_3213# 2.05e-21
C3468 a_4680_3239# a_6010_3239# 5.35e-20
C3469 a_4367_3213# a_6291_3605# 4.38e-20
C3470 a_3452_3239# a_6198_3239# 3.65e-21
C3471 VDD x33.Q_N 0.446f
C3472 x4.X a_11767_4478# 0.00114f
C3473 a_4155_4086# x45.Q_N 1.43e-20
C3474 a_4453_4386# comparator_out 2.5e-20
C3475 a_9442_4086# a_10156_4112# 6.99e-20
C3476 a_8939_4086# a_9377_4112# 0.00276f
C3477 a_9710_4296# a_9954_4478# 0.00972f
C3478 a_8697_4112# a_9578_4112# 0.00943f
C3479 a_9238_4086# a_10681_4086# 2.08e-19
C3480 sel_bit[1] a_621_4112# 1.03e-20
C3481 VDD a_6291_3605# 0.176f
C3482 check[6] a_7247_4775# 2.19e-20
C3483 a_3599_2340# a_4388_2366# 4.2e-20
C3484 a_3912_2366# a_5896_2340# 1.34e-20
C3485 a_7953_3239# D[0] 0.0968f
C3486 x33.Q_N a_8939_4086# 1.3e-22
C3487 a_7246_3213# a_8590_3239# 8.26e-21
C3488 a_9639_4775# check[4] 0.0122f
C3489 a_1682_4775# x4.X 0.176f
C3490 check[2] a_10345_3239# 0.00302f
C3491 eob a_2375_5167# 5.84e-19
C3492 a_9578_4112# a_9709_2550# 1.72e-22
C3493 a_2389_5648# a_2463_4775# 0.00225f
C3494 check[2] a_1976_4775# 0.00168f
C3495 x33.Q_N x60.Q_N 4.08e-19
C3496 check[0] a_4794_4112# 1.51e-19
C3497 VDD a_6304_2366# 0.348f
C3498 a_8683_3605# D[1] 3.23e-21
C3499 a_9151_3213# a_10345_3239# 6.04e-19
C3500 a_11076_5167# a_11331_4086# 2.46e-20
C3501 a_11544_4775# a_11089_4112# 5.67e-20
C3502 a_10795_4801# a_11630_4086# 1.18e-19
C3503 a_11250_4775# a_11629_4386# 3.92e-19
C3504 a_6199_4801# x30.Q_N 4.57e-21
C3505 a_1112_2340# x51.Q_N 0.178f
C3506 D[7] a_2533_2550# 6.45e-20
C3507 a_10629_4801# a_11834_4086# 6.96e-19
C3508 a_2853_5648# x5.X 6.24e-19
C3509 x33.Q_N a_10983_4801# 1e-19
C3510 check[1] a_6466_4775# 5.74e-19
C3511 eob x77.Y 0.05f
C3512 x30.Q_N a_6410_2366# 0.0102f
C3513 check[2] a_12048_4394# 1.36e-20
C3514 a_3913_4112# a_3452_3239# 2.21e-19
C3515 a_3600_4086# a_3618_3239# 3.48e-19
C3516 VDD check[1] 0.762f
C3517 VDD a_8802_2366# 4.84e-19
C3518 VDD a_11389_3239# 5.47e-21
C3519 x30.Q_N x42.Q_N 1.63e-20
C3520 D[1] a_8696_2366# 1.64e-21
C3521 a_6845_2340# a_9237_2340# 0.00176f
C3522 a_6304_2366# x60.Q_N 5.09e-21
C3523 a_10794_3239# a_11856_3239# 0.137f
C3524 a_11075_3605# a_11543_3213# 0.0633f
C3525 a_10628_3239# a_10982_3239# 0.0708f
C3526 x4.X x51.Q_N 0.0098f
C3527 check[5] a_7182_4801# 1.11e-20
C3528 check[1] a_8939_4086# 3.29e-19
C3529 a_4454_4086# D[5] 1.26e-20
C3530 x42.Q_N a_9754_3239# 0.00969f
C3531 x27.Q_N a_4925_2550# 0.181f
C3532 x4.X a_3452_3239# 0.0477f
C3533 x5.X a_6846_4086# 0.261f
C3534 check[4] a_10794_3239# 1.18e-19
C3535 a_2289_4801# a_3453_4801# 6.38e-20
C3536 a_2463_4775# a_3619_4801# 3.31e-19
C3537 a_6199_4801# a_5992_4086# 3.44e-19
C3538 a_7073_4801# a_6305_4112# 3.76e-19
C3539 a_6760_4775# a_6845_4386# 7.46e-19
C3540 a_5845_4801# x45.Q_N 3.67e-20
C3541 a_4367_3213# a_5844_3239# 3.41e-19
C3542 a_3899_3605# comparator_out 1.95e-19
C3543 a_6011_4801# comparator_out 2.9e-21
C3544 a_2289_4801# a_2194_4801# 0.00276f
C3545 a_1415_4801# a_1616_4801# 3.67e-19
C3546 a_2463_4775# a_2697_5083# 0.00945f
C3547 a_1976_4775# x20.Q_N 0.0094f
C3548 VDD a_3877_5674# 3.02e-19
C3549 check[1] x60.Q_N 0.0122f
C3550 x33.Q_N a_8803_4112# 2.89e-22
C3551 x27.Q_N a_4585_3239# 4.03e-19
C3552 a_9237_2340# a_10155_2366# 0.0708f
C3553 a_9441_2340# a_9953_2732# 6.69e-20
C3554 a_9236_2640# D[3] 0.00531f
C3555 a_11075_3605# a_11330_2340# 2.41e-20
C3556 a_11543_3213# a_11088_2366# 3.36e-20
C3557 a_10794_3239# a_11629_2340# 6.38e-20
C3558 a_10628_3239# a_11833_2340# 4.77e-19
C3559 a_11249_3213# a_11628_2640# 2.68e-19
C3560 VDD a_7050_4086# 0.487f
C3561 a_11389_3239# D[2] 1.3e-20
C3562 x4.X a_9638_3213# 0.116f
C3563 VDD a_5844_3239# 0.791f
C3564 a_8998_4801# a_9370_4801# 3.34e-19
C3565 x45.Q_N a_8590_3239# 1.34e-20
C3566 a_7050_4086# a_7362_3239# 5.48e-21
C3567 x4.X a_6985_4112# 6.8e-19
C3568 x20.Q_N D[7] 5.48e-19
C3569 a_3619_4801# a_4453_4386# 7.24e-20
C3570 a_4368_4775# a_3600_4086# 0.0018f
C3571 a_3900_5167# a_3913_4112# 2.81e-19
C3572 a_3453_4801# a_4454_4086# 1.15e-19
C3573 a_4074_4775# a_4155_4086# 8.83e-20
C3574 check[4] a_9577_2366# 4.82e-19
C3575 a_6845_4386# a_9238_4086# 2.9e-21
C3576 x45.Q_N a_8384_4086# 5.27e-21
C3577 a_8697_4112# comparator_out 2.29e-20
C3578 x20.Q_N a_4155_4086# 2.32e-19
C3579 x36.Q_N a_11075_3605# 0.00192f
C3580 check[0] a_6505_4394# 9.42e-20
C3581 a_1626_2366# D[6] 3.23e-20
C3582 a_1762_2340# a_2200_2366# 0.00276f
C3583 a_1520_2366# a_2401_2366# 0.00943f
C3584 a_2061_2340# a_3504_2340# 8.18e-19
C3585 check[0] x75.Q 0.0176f
C3586 a_6400_4801# check[5] 5.31e-21
C3587 a_11088_2366# a_11330_2340# 0.124f
C3588 a_10775_2340# a_11628_2640# 0.0264f
C3589 a_10680_2340# x63.Q_N 0.178f
C3590 x4.X a_9236_2640# 0.00898f
C3591 check[4] a_11184_4801# 9.44e-20
C3592 comparator_out a_12737_3239# 1.9e-19
C3593 comparator_out a_9709_2550# 0.00825f
C3594 a_4019_4112# a_4389_4112# 4.11e-20
C3595 a_5170_4478# a_5372_4112# 8.94e-19
C3596 x4.X a_3900_5167# 0.00135f
C3597 check[2] a_5845_4801# 1.76e-19
C3598 x4.X a_11076_5167# 0.00135f
C3599 x36.Q_N a_11088_2366# 0.0928f
C3600 a_3452_3239# a_3618_3239# 0.638f
C3601 VDD a_2061_2340# 0.853f
C3602 a_3912_2366# a_4590_2732# 0.00652f
C3603 a_4154_2340# a_4388_2732# 0.00976f
C3604 a_3599_2340# a_4018_2366# 0.0397f
C3605 a_5089_5083# x27.Q_N 2.02e-20
C3606 a_4970_3239# a_4657_2340# 3.49e-20
C3607 VDD a_1338_5674# 0.255f
C3608 x4.X a_12345_2732# 1.17e-19
C3609 check[1] a_8803_4112# 4.26e-19
C3610 a_4854_3213# a_5371_2366# 2.38e-19
C3611 check[6] a_4592_2366# 8.47e-20
C3612 a_11331_4086# a_11543_3213# 2.12e-19
C3613 a_11089_4112# a_12030_3213# 9.49e-19
C3614 a_11834_4086# a_10794_3239# 2.9e-19
C3615 a_11630_4086# a_11249_3213# 5.04e-19
C3616 a_12265_5083# x36.Q_N 2.02e-20
C3617 x5.X a_7562_4478# 1.85e-19
C3618 check[2] a_8384_4086# 6.25e-20
C3619 x30.Q_N a_6465_3213# 5.84e-19
C3620 a_4213_3239# a_4789_3239# 2.46e-21
C3621 sel_bit[0] a_2788_5674# 3.68e-19
C3622 VDD D[5] 0.221f
C3623 a_5371_2366# a_5169_2366# 3.67e-19
C3624 VDD a_8857_3213# 0.308f
C3625 check[0] a_4926_4296# 0.00111f
C3626 VDD x72.Q_N 0.0716f
C3627 a_4388_2366# a_4793_2366# 2.46e-21
C3628 a_5896_2340# a_5991_2340# 0.0968f
C3629 check[4] a_10776_4086# 0.00416f
C3630 a_9638_3213# a_9464_3239# 0.197f
C3631 a_8683_3605# a_8767_3605# 0.00972f
C3632 a_8236_3239# a_9101_3521# 0.00276f
C3633 a_9151_3213# a_8590_3239# 3.79e-20
C3634 VDD a_7764_4112# 0.109f
C3635 a_8697_4112# a_8683_3605# 1.61e-19
C3636 a_9238_4086# a_8236_3239# 6.54e-20
C3637 a_8939_4086# a_8857_3213# 1.02e-19
C3638 a_8384_4086# a_9151_3213# 8.83e-19
C3639 a_9237_4386# a_8402_3239# 4.11e-20
C3640 x4.X a_7562_4112# 6.4e-19
C3641 a_11629_4386# a_11088_2366# 1.93e-22
C3642 x30.Q_N a_5991_2340# 0.142f
C3643 a_6985_4112# a_7186_4112# 3.34e-19
C3644 a_8289_4086# a_8697_4112# 4.37e-19
C3645 check[2] a_4855_4775# 2.07e-19
C3646 a_897_4112# a_1511_4112# 9.05e-20
C3647 a_4368_4775# a_3452_3239# 9.66e-21
C3648 a_3900_5167# a_3618_3239# 1.65e-21
C3649 a_4074_4775# a_4073_3213# 2.59e-19
C3650 a_3619_4801# a_3899_3605# 8.52e-21
C3651 VDD a_8383_2340# 0.561f
C3652 x20.Q_N a_4073_3213# 8.02e-21
C3653 D[1] a_11249_3213# 8.77e-20
C3654 a_8237_4801# a_8858_4775# 0.117f
C3655 a_9464_3239# a_9236_2640# 1.11e-20
C3656 a_9151_3213# a_9441_2340# 0.00144f
C3657 a_9638_3213# a_9237_2340# 8.72e-19
C3658 x69.Q_N D[1] 2.5e-19
C3659 VDD a_3453_4801# 0.841f
C3660 x36.Q_N a_11331_4086# 1.3e-22
C3661 check[2] a_11564_2366# 1.34e-19
C3662 a_5992_4086# a_6465_3213# 2.45e-19
C3663 a_6305_4112# a_6010_3239# 4.9e-19
C3664 a_4454_4086# a_4453_2340# 1.55e-19
C3665 a_4453_4386# a_4657_2340# 1.26e-21
C3666 VDD a_2194_4801# 0.00214f
C3667 a_8697_4112# a_8696_2366# 1.8e-19
C3668 a_8939_4086# a_8383_2340# 1.3e-22
C3669 VDD a_10629_4801# 0.81f
C3670 check[1] a_7481_5083# 4.45e-19
C3671 a_1061_4801# a_897_4112# 0.00384f
C3672 a_897_4112# comparator_out 7.09e-20
C3673 VDD a_11766_2732# 0.0163f
C3674 x48.Q a_4318_5083# 4.61e-19
C3675 a_4971_4801# a_4658_4086# 7.76e-20
C3676 x77.Y a_3806_3239# 0.0112f
C3677 D[1] a_10775_2340# 0.00122f
C3678 x4.X D[0] 0.0011f
C3679 a_8696_2366# a_9709_2550# 0.0633f
C3680 a_9236_2640# a_9237_2340# 0.781f
C3681 a_8383_2340# x60.Q_N 0.124f
C3682 a_8938_2340# a_9441_2340# 0.00187f
C3683 a_11856_3239# a_12146_3239# 0.0282f
C3684 a_12030_3213# a_11965_3239# 4.2e-20
C3685 x4.X x54.Q_N 0.00996f
C3686 a_10982_3239# a_11183_3239# 3.67e-19
C3687 a_11856_3239# a_11761_3239# 0.00276f
C3688 a_11543_3213# x66.Q_N 0.00553f
C3689 a_12030_3213# a_12264_3521# 0.00945f
C3690 a_5992_4086# a_5991_2340# 5.27e-19
C3691 x27.Q_N a_7049_2340# 8.08e-21
C3692 x4.X a_5088_3521# 0.0012f
C3693 a_3619_4801# a_4681_4801# 0.137f
C3694 a_3900_5167# a_4368_4775# 0.0633f
C3695 a_3453_4801# a_3807_4801# 0.0662f
C3696 eob D[6] 8.49e-20
C3697 x30.Q_N a_6846_4086# 0.0258f
C3698 a_9377_4112# x39.Q_N 2.88e-20
C3699 x5.X a_9152_4775# 0.00142f
C3700 a_11089_4112# a_11630_4086# 0.125f
C3701 a_11331_4086# a_11629_4386# 0.137f
C3702 check[1] a_3258_5648# 0.0414f
C3703 a_2853_5648# a_3373_5674# 0.394f
C3704 a_2061_2340# a_2198_2732# 0.00907f
C3705 D[3] a_11330_2340# 1.99e-19
C3706 check[1] sel_bit[1] 0.26f
C3707 a_5845_4801# a_8591_4801# 3.65e-21
C3708 a_7073_4801# a_8403_4801# 4e-20
C3709 x33.Q_N x39.Q_N 2.41e-20
C3710 x4.X a_11543_3213# 0.111f
C3711 a_10629_4801# a_10983_4801# 0.0665f
C3712 a_11076_5167# a_11544_4775# 0.0633f
C3713 a_10795_4801# a_11857_4801# 0.137f
C3714 a_8803_4112# a_8857_3213# 3.34e-20
C3715 comparator_out a_10982_3239# 0.157f
C3716 VDD a_9639_4775# 0.72f
C3717 x48.Q_N a_4113_4394# 2.02e-20
C3718 a_4658_4086# a_4591_4478# 9.46e-19
C3719 a_3913_4112# a_5372_4112# 1.65e-21
C3720 a_4453_4386# a_4872_4394# 2.46e-19
C3721 x27.Q_N a_3913_4112# 1.32e-21
C3722 x36.Q_N D[3] 0.00274f
C3723 a_9152_4775# a_9237_4386# 7.46e-19
C3724 a_8237_4801# x42.Q_N 3.67e-20
C3725 a_8591_4801# a_8384_4086# 3.44e-19
C3726 a_9465_4801# a_8697_4112# 3.76e-19
C3727 x36.Q_N x66.Q_N 0.02f
C3728 a_3504_2340# a_4453_2340# 1.03e-19
C3729 a_12345_2732# a_12547_2366# 8.94e-19
C3730 a_3373_5674# a_3671_5674# 0.00489f
C3731 a_6010_3239# a_6605_3239# 0.00118f
C3732 a_6198_3239# a_6375_3605# 8.94e-19
C3733 a_6759_3213# a_6709_3521# 1.21e-20
C3734 x4.X a_11330_2340# 0.0071f
C3735 x36.Q_N a_11195_4112# 2.89e-22
C3736 x4.X a_5372_4112# 0.00623f
C3737 a_5561_3239# a_6759_3213# 5.62e-20
C3738 comparator_out a_11833_2340# 0.00593f
C3739 a_4367_3213# a_4453_2340# 2.19e-19
C3740 a_4854_3213# a_4452_2640# 3.43e-19
C3741 a_6305_4112# a_6845_4386# 0.139f
C3742 a_5992_4086# a_6846_4086# 0.0492f
C3743 x4.X x27.Q_N 0.425f
C3744 a_2853_5648# eob 0.00163f
C3745 VDD a_4453_2340# 0.788f
C3746 x4.X x36.Q_N 0.278f
C3747 a_4452_2640# a_5169_2366# 0.00105f
C3748 a_4854_3213# a_4766_3605# 7.71e-20
C3749 a_4073_3213# a_4585_3239# 9.75e-19
C3750 a_4680_3239# a_4538_3521# 0.00412f
C3751 a_3899_3605# a_4007_3239# 0.00812f
C3752 a_4367_3213# a_4213_3239# 0.00943f
C3753 a_6011_4801# a_6710_5083# 2.46e-19
C3754 a_5845_4801# a_6931_5083# 0.00907f
C3755 a_3452_3239# x75.Q_N 1.07e-19
C3756 D[0] a_9464_3239# 3.72e-20
C3757 a_9639_4775# a_10983_4801# 8.26e-21
C3758 x5.X a_10628_3239# 9.1e-20
C3759 x20.Q_N a_1720_2648# 2.75e-19
C3760 VDD a_4790_4801# 9.01e-19
C3761 VDD a_4213_3239# 0.00187f
C3762 a_11834_4086# a_12146_3239# 5.48e-21
C3763 x30.Q_N a_5371_2366# 1.34e-20
C3764 x39.Q_N a_11389_3239# 0.0314f
C3765 x30.Q_N a_8402_3239# 3.97e-20
C3766 VDD a_7763_2366# 0.109f
C3767 check[2] check[4] 0.347f
C3768 a_11630_4086# a_11767_4478# 0.00907f
C3769 VDD a_10794_3239# 0.274f
C3770 x39.Q_N a_9954_4112# 2.57e-20
C3771 VDD a_9872_3521# 0.00506f
C3772 D[0] a_9237_2340# 1.09e-20
C3773 a_6845_2340# x57.Q_N 1.07e-19
C3774 a_7049_2340# a_7317_2550# 0.205f
C3775 check[2] a_11629_2340# 1.99e-19
C3776 a_2389_5648# a_2969_6040# 0.00342f
C3777 a_1338_5674# sel_bit[1] 0.0421f
C3778 check[2] a_2883_5674# 0.0516f
C3779 x42.Q_N a_9322_3521# 0.00203f
C3780 x5.X a_4591_4478# 1.55e-19
C3781 x4.X a_11629_4386# 0.0479f
C3782 x30.Q_N a_7185_2366# 0.0403f
C3783 check[4] a_9151_3213# 1.06e-19
C3784 a_10346_4801# a_9638_3213# 3.19e-20
C3785 a_9442_4086# x42.Q_N 0.00116f
C3786 a_1508_5167# a_1976_4775# 0.0627f
C3787 check[6] x77.Y 3.89e-20
C3788 x27.Q_N a_3618_3239# 3.65e-19
C3789 a_5089_5083# a_5845_4801# 4.06e-20
C3790 a_10345_3239# D[3] 0.00127f
C3791 a_10794_3239# D[2] 5.71e-21
C3792 D[1] a_11965_3239# 1.23e-20
C3793 D[4] a_9709_2550# 1.83e-20
C3794 x5.X a_11390_4801# 9.46e-19
C3795 VDD a_4019_4112# 0.0124f
C3796 x4.X a_6375_3605# 9.07e-19
C3797 a_8684_5167# a_8998_4801# 0.0258f
C3798 a_8403_4801# a_9370_4801# 0.00126f
C3799 a_8237_4801# a_9873_5083# 1.25e-19
C3800 a_9152_4775# a_9551_5167# 0.00133f
C3801 reset x3.A 0.00364f
C3802 comparator_out a_4112_2648# 1.53e-19
C3803 VDD a_4008_4801# 2.82e-19
C3804 VDD x3.A 0.203f
C3805 x48.Q a_2993_5674# 1.96e-19
C3806 a_5844_3239# a_6930_3521# 0.00907f
C3807 a_6845_4386# a_6983_4478# 1.09e-19
C3808 a_6305_4112# a_7264_4394# 1.21e-20
C3809 a_6547_4086# a_6411_4112# 0.0282f
C3810 check[4] a_8938_2340# 1.33e-19
C3811 a_11544_4775# a_11543_3213# 0.00121f
C3812 x75.Q a_5844_3239# 0.335f
C3813 a_5561_3239# comparator_out 0.00108f
C3814 x5.X a_7954_4801# 0.0293f
C3815 eob a_2060_2640# 1.44e-19
C3816 a_6466_4775# check[5] 1.71e-20
C3817 a_1207_2340# a_1762_2340# 0.197f
C3818 check[0] a_5562_4801# 0.0162f
C3819 a_9441_2340# a_11088_2366# 7.2e-21
C3820 a_9237_2340# a_11330_2340# 6.38e-20
C3821 a_9709_2550# a_10775_2340# 7.98e-21
C3822 x4.X a_10345_3239# 0.00275f
C3823 a_1112_2340# D[7] 0.0786f
C3824 x4.X a_7317_2550# 0.00147f
C3825 check[1] a_4926_4296# 1.97e-22
C3826 check[4] a_11250_4775# 6.31e-19
C3827 VDD check[5] 0.493f
C3828 a_1061_4801# a_1415_4801# 0.0708f
C3829 x4.X a_1976_4775# 0.0979f
C3830 a_1227_4801# a_2289_4801# 0.137f
C3831 sel_bit[1] a_3453_4801# 0.00123f
C3832 a_3505_4086# a_4454_4086# 1.03e-19
C3833 a_3600_4086# a_4453_4386# 0.0264f
C3834 a_3913_4112# a_4155_4086# 0.124f
C3835 a_2883_5674# x20.Q_N 5.75e-20
C3836 check[2] a_11834_4086# 1.08e-19
C3837 x36.Q_N a_9237_2340# 1.55e-19
C3838 a_4681_4801# a_4586_4801# 0.00276f
C3839 a_3807_4801# a_4008_4801# 3.67e-19
C3840 a_4855_4775# a_5089_5083# 0.00945f
C3841 a_4368_4775# x27.Q_N 0.00773f
C3842 D[6] a_2401_2366# 5.27e-19
C3843 a_2979_2366# a_3599_2340# 8.26e-21
C3844 a_2533_2550# a_2777_2366# 0.00812f
C3845 a_11088_2366# a_11564_2366# 2.87e-21
C3846 a_11629_2340# a_12047_2648# 0.00276f
C3847 a_11628_2640# a_12345_2732# 4.45e-20
C3848 x4.X D[7] 0.00353f
C3849 VDD a_10776_4086# 0.716f
C3850 x4.X a_4155_4086# 0.00873f
C3851 a_1062_5674# a_1061_4801# 0.00165f
C3852 check[6] a_3912_2366# 1.31e-20
C3853 a_11544_4775# x36.Q_N 0.0059f
C3854 a_12031_4775# a_12265_5083# 0.00945f
C3855 a_10983_4801# a_11184_4801# 3.67e-19
C3856 a_11857_4801# a_11762_4801# 0.00276f
C3857 a_7073_4801# a_6010_3239# 6.75e-21
C3858 a_4854_3213# a_6759_3213# 3.71e-20
C3859 x4.X a_12048_4394# 8.47e-19
C3860 check[0] a_7561_2366# 1.87e-20
C3861 a_4454_4086# x45.Q_N 3.85e-19
C3862 a_4658_4086# comparator_out 4.39e-21
C3863 x36.Q_N a_12547_2366# 0.0317f
C3864 x42.Q_N a_10156_4112# 8.23e-20
C3865 a_9238_4086# a_9377_4112# 2.56e-19
C3866 a_9237_4386# a_9578_4112# 0.00118f
C3867 a_8939_4086# a_10776_4086# 1.86e-21
C3868 VDD a_7246_3213# 0.569f
C3869 check[6] a_6199_4801# 0.165f
C3870 a_4154_2340# a_4388_2366# 0.00707f
C3871 a_3912_2366# a_4592_2366# 3.73e-19
C3872 a_4452_2640# a_5896_2340# 6.96e-19
C3873 x33.Q_N a_9238_4086# 0.026f
C3874 a_7246_3213# a_7362_3239# 0.0397f
C3875 a_6759_3213# a_7181_3239# 2.87e-21
C3876 a_6605_3239# a_6977_3239# 3.34e-19
C3877 check[1] x27.D 1.12e-20
C3878 eob a_1616_4801# 4.1e-19
C3879 x75.Q D[5] 9.96e-19
C3880 x30.Q_N a_4452_2640# 0.00116f
C3881 check[0] a_3876_6040# 2.26e-19
C3882 a_3170_4801# a_1511_4112# 5.42e-19
C3883 check[0] a_6305_4112# 0.00126f
C3884 VDD a_6844_2640# 0.269f
C3885 a_5991_2340# a_6780_2732# 7.71e-20
C3886 a_6304_2366# a_6504_2648# 0.00185f
C3887 a_8236_3239# a_8288_2340# 4.5e-19
C3888 a_9638_3213# D[1] 0.0115f
C3889 a_11857_4801# a_11089_4112# 3.76e-19
C3890 a_10983_4801# a_10776_4086# 3.44e-19
C3891 a_11544_4775# a_11629_4386# 7.46e-19
C3892 a_10629_4801# x39.Q_N 3.68e-20
C3893 a_7362_3239# a_6844_2640# 5.05e-21
C3894 a_5088_3521# x75.Q_N 2.02e-20
C3895 a_3505_4086# a_3504_2340# 1.07e-20
C3896 a_7186_4112# a_7317_2550# 1.72e-22
C3897 x33.Q_N a_9755_4801# 3.78e-19
C3898 check[1] a_6760_4775# 0.00254f
C3899 a_1062_5674# a_2389_5648# 1.61e-20
C3900 a_1061_4801# a_3170_4801# 1.03e-19
C3901 x5.A a_1338_5674# 0.263f
C3902 check[2] a_4454_4086# 2.36e-20
C3903 x5.X a_1511_4112# 2.24e-19
C3904 a_3913_4112# a_4073_3213# 0.00148f
C3905 a_4155_4086# a_3618_3239# 1.07e-20
C3906 a_4453_4386# a_3452_3239# 6.5e-20
C3907 x5.X a_11289_4394# 4.41e-19
C3908 VDD a_9953_2732# 0.0042f
C3909 a_4539_5083# check[6] 1.43e-21
C3910 VDD a_12146_3239# 4.88e-19
C3911 VDD a_11761_3239# 6.2e-19
C3912 D[1] a_9236_2640# 5.41e-19
C3913 a_10345_3239# a_9237_2340# 4.83e-19
C3914 VDD a_3505_4086# 0.212f
C3915 a_6844_2640# x60.Q_N 1.38e-19
C3916 a_11543_3213# a_12030_3213# 0.273f
C3917 a_11249_3213# a_10982_3239# 6.99e-20
C3918 a_10794_3239# a_11159_3605# 4.45e-20
C3919 check[1] a_9238_4086# 2.12e-19
C3920 VDD a_11565_4478# 0.00371f
C3921 x5.X a_1061_4801# 0.265f
C3922 a_11715_5083# check[3] 9.55e-19
C3923 x4.X a_4073_3213# 0.00798f
C3924 x4.X a_5845_4801# 0.00422f
C3925 x30.Q_N a_9376_2366# 2.98e-20
C3926 x5.X a_7318_4296# 6.4e-19
C3927 x5.X comparator_out 6.13e-20
C3928 a_2463_4775# a_3900_5167# 7.98e-21
C3929 a_7247_4775# a_6846_4086# 0.00169f
C3930 a_6466_4775# x45.Q_N 2.19e-19
C3931 a_6760_4775# a_7050_4086# 0.00268f
C3932 x45.Q_N a_4367_3213# 3.74e-20
C3933 a_7073_4801# a_6845_4386# 1.96e-20
C3934 a_4854_3213# comparator_out 0.00379f
C3935 a_4680_3239# a_5844_3239# 6.38e-20
C3936 a_6760_4775# a_5844_3239# 9.66e-21
C3937 x4.X a_12147_4801# 0.00557f
C3938 a_2289_4801# x20.Q_N 8.79e-19
C3939 VDD a_1227_4801# 0.34f
C3940 D[2] a_12146_3239# 9.48e-20
C3941 x27.Q_N a_6606_4801# 1.93e-20
C3942 x27.Q_N x75.Q_N 0.02f
C3943 a_9709_2550# a_10155_2366# 0.0367f
C3944 a_11543_3213# a_11628_2640# 5.32e-19
C3945 a_10982_3239# a_10775_2340# 2.02e-19
C3946 a_11856_3239# a_11088_2366# 2.17e-19
C3947 x4.X a_8590_3239# 0.0062f
C3948 a_11761_3239# D[2] 1.36e-20
C3949 VDD x45.Q_N 0.458f
C3950 a_8998_4801# x33.Q_N 4.01e-20
C3951 x45.Q_N a_7362_3239# 0.00968f
C3952 x4.X a_8384_4086# 0.101f
C3953 a_8237_4801# a_8402_3239# 8.16e-19
C3954 a_8403_4801# a_8236_3239# 9.04e-19
C3955 a_2389_5648# a_3170_4801# 1.39e-19
C3956 a_4855_4775# a_3913_4112# 0.00161f
C3957 a_4368_4775# a_4155_4086# 3.72e-19
C3958 a_4074_4775# a_4454_4086# 0.00336f
C3959 a_3619_4801# a_4658_4086# 0.00221f
C3960 check[4] a_11088_2366# 2.47e-20
C3961 a_6547_4086# x42.Q_N 7.23e-21
C3962 a_9237_4386# comparator_out 2.49e-20
C3963 x20.Q_N a_4454_4086# 1.21e-19
C3964 a_12031_4775# x66.Q_N 4.45e-20
C3965 x36.Q_N a_12030_3213# 0.0126f
C3966 check[0] a_6983_4478# 6.27e-20
C3967 x48.Q check[0] 0.0102f
C3968 a_2061_2340# a_2200_2366# 2.56e-19
C3969 a_2060_2640# a_2401_2366# 0.00118f
C3970 a_1762_2340# a_3599_2340# 1.86e-21
C3971 D[3] a_11564_2366# 3.38e-20
C3972 a_1520_2366# a_3912_2366# 6.12e-21
C3973 x30.Q_N a_7954_4801# 0.182f
C3974 a_7481_5083# check[5] 1.93e-21
C3975 a_11330_2340# a_11628_2640# 0.137f
C3976 a_11088_2366# a_11629_2340# 0.125f
C3977 x4.X a_9441_2340# 0.00148f
C3978 x4.X a_4855_4775# 0.102f
C3979 a_1227_4801# a_3807_4801# 3.07e-21
C3980 a_2389_5648# x5.X 0.00112f
C3981 sel_bit[0] a_2853_5648# 1.09f
C3982 sel_bit[1] x3.A 1.43e-20
C3983 check[2] a_6466_4775# 1.08e-19
C3984 x4.X a_12031_4775# 0.0991f
C3985 x36.Q_N a_11628_2640# 0.572f
C3986 a_3618_3239# a_4073_3213# 0.149f
C3987 a_3452_3239# a_3899_3605# 0.141f
C3988 VDD a_2533_2550# 0.194f
C3989 a_4452_2640# a_4590_2732# 1.09e-19
C3990 a_3912_2366# a_4871_2648# 1.21e-20
C3991 a_4154_2340# a_4018_2366# 0.0282f
C3992 D[6] a_4592_2366# 3.35e-19
C3993 VDD check[2] 0.713f
C3994 clk_sar reset 1.31e-20
C3995 VDD clk_sar 0.114f
C3996 check[6] a_5991_2340# 1.42e-21
C3997 x39.Q_N a_10794_3239# 0.348f
C3998 a_11630_4086# a_11543_3213# 1.61e-19
C3999 a_11629_4386# a_12030_3213# 3.78e-19
C4000 x5.X a_8289_4086# 0.0767f
C4001 check[2] a_8939_4086# 5.79e-20
C4002 x30.Q_N a_6759_3213# 0.00506f
C4003 a_3170_4801# a_3619_4801# 6.24e-19
C4004 x27.D a_3453_4801# 0.412f
C4005 x33.Q_N a_9573_3239# 1.68e-19
C4006 VDD a_9151_3213# 0.353f
C4007 a_8857_3213# a_9101_3521# 0.0104f
C4008 a_8402_3239# a_9322_3521# 1.09e-19
C4009 VDD a_6781_4112# 3.56e-19
C4010 check[1] a_5562_4801# 3.76e-20
C4011 a_9238_4086# a_8857_3213# 5.04e-19
C4012 a_9442_4086# a_8402_3239# 2.9e-19
C4013 a_8697_4112# a_9638_3213# 9.49e-19
C4014 a_8939_4086# a_9151_3213# 2.12e-19
C4015 x4.X a_9173_4478# 2.12e-19
C4016 x20.Q_N a_3504_2340# 6.66e-19
C4017 a_11629_4386# a_11628_2640# 1.32e-20
C4018 a_11630_4086# a_11330_2340# 3.47e-21
C4019 a_11834_4086# a_11088_2366# 7.14e-22
C4020 x5.X a_3619_4801# 0.0076f
C4021 x30.Q_N a_6546_2340# 0.16f
C4022 a_7764_4112# a_9238_4086# 3.65e-21
C4023 a_8289_4086# a_9237_4386# 9.65e-21
C4024 x5.X a_2697_5083# 3.53e-19
C4025 x4.X a_7182_4801# 2.39e-19
C4026 a_4368_4775# a_5845_4801# 1.72e-19
C4027 a_3453_4801# a_4680_3239# 4.76e-21
C4028 a_4074_4775# a_4367_3213# 7.57e-21
C4029 x5.X a_10795_4801# 0.0203f
C4030 VDD a_8938_2340# 0.177f
C4031 a_6410_2366# a_6780_2366# 4.11e-20
C4032 x20.Q_N a_4367_3213# 1.25e-21
C4033 x4.X a_1720_2648# 0.00102f
C4034 D[1] a_11543_3213# 1.24e-19
C4035 a_8237_4801# a_9152_4775# 0.125f
C4036 a_8403_4801# a_8684_5167# 0.155f
C4037 a_9638_3213# a_9709_2550# 1.66e-21
C4038 a_9464_3239# a_9441_2340# 1.03e-19
C4039 VDD a_4074_4775# 0.494f
C4040 x36.Q_N a_11630_4086# 0.0255f
C4041 a_6305_4112# a_6291_3605# 1.61e-19
C4042 a_6547_4086# a_6465_3213# 1.02e-19
C4043 a_5992_4086# a_6759_3213# 8.83e-19
C4044 a_6845_4386# a_6010_3239# 4.11e-20
C4045 VDD x20.Q_N 1.29f
C4046 check[2] a_11969_2366# 4.38e-19
C4047 a_4926_4296# a_4453_2340# 6.08e-21
C4048 a_9237_4386# a_8696_2366# 1.93e-22
C4049 a_11544_4775# a_12147_4801# 0.0552f
C4050 VDD a_11250_4775# 0.488f
C4051 x77.Y a_3912_2366# 7.49e-20
C4052 x48.Q a_4389_4478# 3.17e-19
C4053 x27.Q_N a_4970_3239# 0.00341f
C4054 a_10346_4801# a_10345_3239# 9.85e-20
C4055 check[6] a_6846_4086# 2.07e-22
C4056 x48.Q a_4767_5167# 1.31e-19
C4057 VDD a_12047_2648# 0.00984f
C4058 x77.Y a_4317_3521# 4.28e-20
C4059 a_9237_2340# a_9441_2340# 0.117f
C4060 a_9236_2640# a_9709_2550# 0.145f
C4061 a_8938_2340# x60.Q_N 9.58e-21
C4062 a_11856_3239# x66.Q_N 9.58e-21
C4063 a_6305_4112# a_6304_2366# 1.8e-19
C4064 a_6547_4086# a_5991_2340# 1.3e-22
C4065 comparator_out a_5896_2340# 7.85e-19
C4066 x27.Q_N x57.Q_N 7.46e-20
C4067 check[4] D[3] 0.00432f
C4068 x4.X a_6400_4801# 8.46e-20
C4069 check[2] a_8803_4112# 1.27e-20
C4070 a_4074_4775# a_3807_4801# 6.99e-20
C4071 a_4368_4775# a_4855_4775# 0.273f
C4072 a_3619_4801# a_3984_5167# 4.45e-20
C4073 x36.Q_N D[1] 1.36e-20
C4074 x20.Q_N a_3807_4801# 1.92e-19
C4075 x5.X a_9465_4801# 0.00117f
C4076 check[2] a_9323_5083# 4.69e-19
C4077 a_10776_4086# x39.Q_N 0.155f
C4078 a_11331_4086# a_11834_4086# 0.00187f
C4079 a_11629_4386# a_11630_4086# 0.782f
C4080 a_11089_4112# a_12102_4296# 0.0633f
C4081 x30.Q_N a_7318_4296# 5.71e-19
C4082 x30.Q_N comparator_out 0.274f
C4083 a_2061_2340# a_2479_2648# 0.00276f
C4084 a_2060_2640# a_2777_2732# 4.45e-20
C4085 a_1520_2366# D[6] 6.36e-20
C4086 D[3] a_11629_2340# 1.1e-19
C4087 check[1] a_6305_4112# 0.00312f
C4088 a_12146_3239# a_12101_2550# 1.01e-20
C4089 x4.X a_11856_3239# 0.00481f
C4090 sel_bit[1] a_3505_4086# 1.09e-19
C4091 a_10795_4801# a_11160_5167# 4.45e-20
C4092 a_11250_4775# a_10983_4801# 6.99e-20
C4093 a_11544_4775# a_12031_4775# 0.273f
C4094 VDD a_8591_4801# 0.109f
C4095 a_4454_4086# a_5170_4478# 0.0018f
C4096 a_3913_4112# a_4389_4112# 2.87e-21
C4097 a_4658_4086# a_4872_4394# 0.0104f
C4098 a_4453_4386# a_5372_4112# 0.162f
C4099 a_8384_4086# a_8897_4394# 0.00945f
C4100 x4.X check[4] 0.037f
C4101 x27.Q_N a_4453_4386# 0.0318f
C4102 a_9465_4801# a_9237_4386# 1.96e-20
C4103 a_9152_4775# a_9442_4086# 0.00268f
C4104 a_9639_4775# a_9238_4086# 0.00169f
C4105 a_8858_4775# x42.Q_N 2.19e-19
C4106 a_3599_2340# a_4154_2340# 0.197f
C4107 a_6010_3239# a_8236_3239# 4e-20
C4108 a_6759_3213# a_7158_3605# 0.00133f
C4109 a_6010_3239# a_6977_3239# 0.00126f
C4110 a_6291_3605# a_6605_3239# 0.0258f
C4111 sel_bit[1] a_1227_4801# 3.62e-20
C4112 x4.X a_11629_2340# 0.00254f
C4113 x4.X a_4389_4112# 3.84e-19
C4114 a_6411_4112# a_6465_3213# 3.34e-20
C4115 check[6] a_5371_2366# 0.00326f
C4116 comparator_out x63.Q_N 2.11e-19
C4117 a_4367_3213# a_4925_2550# 1.62e-19
C4118 a_4854_3213# a_4657_2340# 2.52e-19
C4119 a_6547_4086# a_6846_4086# 0.0334f
C4120 a_6305_4112# a_7050_4086# 0.199f
C4121 a_5992_4086# a_7318_4296# 4.7e-22
C4122 a_4794_4112# x45.Q_N 5.94e-20
C4123 a_6305_4112# a_5844_3239# 2.21e-19
C4124 a_5992_4086# comparator_out 0.00201f
C4125 x33.Q_N a_8288_2340# 3.7e-19
C4126 x5.X a_6710_5083# 3.44e-19
C4127 VDD a_7953_3239# 0.19f
C4128 VDD a_4925_2550# 0.174f
C4129 a_4453_2340# a_6504_2648# 4.06e-20
C4130 a_5845_4801# a_6606_4801# 6.04e-20
C4131 a_6011_4801# a_7159_5167# 2.13e-19
C4132 a_6466_4775# a_6931_5083# 9.46e-19
C4133 check[0] a_4318_5083# 1.54e-19
C4134 a_4367_3213# a_4585_3239# 3.73e-19
C4135 a_4680_3239# a_4213_3239# 0.00316f
C4136 eob a_1511_4112# 0.0585f
C4137 x5.X D[4] 3.43e-19
C4138 a_9639_4775# a_9755_4801# 0.0397f
C4139 a_9152_4775# a_9574_4801# 2.87e-21
C4140 VDD a_6931_5083# 0.0163f
C4141 VDD a_4585_3239# 0.00112f
C4142 x20.Q_N a_2198_2732# 0.00203f
C4143 x39.Q_N a_12146_3239# 0.00968f
C4144 x4.A a_1511_4112# 0.619f
C4145 x39.Q_N a_11761_3239# 0.00399f
C4146 a_3453_4801# a_5562_4801# 1.03e-19
C4147 eob a_1061_4801# 0.514f
C4148 a_11089_4112# a_11565_4112# 2.87e-21
C4149 a_11630_4086# a_12048_4394# 0.00276f
C4150 a_11629_4386# a_12346_4478# 4.45e-20
C4151 VDD a_11075_3605# 0.176f
C4152 a_6304_2366# a_8288_2340# 8.55e-21
C4153 a_5991_2340# a_6780_2366# 4.2e-20
C4154 a_7954_4801# a_8237_4801# 8.18e-19
C4155 a_10345_3239# D[1] 0.0968f
C4156 check[1] a_6983_4478# 9.03e-21
C4157 a_9638_3213# a_10982_3239# 8.26e-21
C4158 check[2] a_3258_5648# 0.0201f
C4159 eob comparator_out 3.93e-19
C4160 a_2389_5648# a_3373_5674# 0.176f
C4161 check[1] x48.Q 0.0512f
C4162 check[2] sel_bit[1] 0.393f
C4163 a_1061_4801# x4.A 0.00353f
C4164 check[2] a_12101_2550# 2.02e-19
C4165 a_10629_4801# a_12738_4801# 9.94e-20
C4166 clk_sar sel_bit[1] 0.329f
C4167 x5.X a_4872_4394# 1.11e-19
C4168 x77.Y D[6] 4.91e-19
C4169 x42.Q_N a_8997_3239# 0.0309f
C4170 x4.X a_11834_4086# 0.00986f
C4171 a_5845_4801# a_5897_4086# 6.04e-19
C4172 x30.Q_N a_8696_2366# 8.85e-20
C4173 x4.A comparator_out 1.12e-19
C4174 a_1976_4775# a_2463_4775# 0.271f
C4175 x27.Q_N a_6011_4801# 1.48e-19
C4176 VDD a_11088_2366# 0.348f
C4177 check[1] a_8288_2340# 0.027f
C4178 x27.Q_N a_3899_3605# 0.00192f
C4179 a_4855_4775# x75.Q_N 4.45e-20
C4180 VDD a_5170_4478# 0.00436f
C4181 x5.X a_11762_4801# 2.61e-19
C4182 a_11543_3213# a_12737_3239# 6.04e-19
C4183 a_11075_3605# D[2] 3.24e-21
C4184 x4.X a_4789_3239# 1.05e-19
C4185 a_9465_4801# a_9551_5167# 0.00976f
C4186 a_7363_4801# a_7182_4801# 4.11e-20
C4187 a_8403_4801# x33.Q_N 2.97e-20
C4188 comparator_out a_4590_2732# 9.45e-19
C4189 VDD a_5089_5083# 0.00529f
C4190 x48.Q a_3877_5674# 4.02e-19
C4191 x45.Q_N a_6930_3521# 0.00203f
C4192 a_5844_3239# a_6605_3239# 6.04e-20
C4193 x36.Q_N a_11966_4801# 7.29e-21
C4194 a_6305_4112# a_7764_4112# 1.65e-21
C4195 a_6845_4386# a_7264_4394# 2.46e-19
C4196 x45.Q_N a_6505_4394# 2.02e-20
C4197 a_7050_4086# a_6983_4478# 9.46e-19
C4198 VDD a_12265_5083# 0.00506f
C4199 check[0] a_6010_3239# 0.0252f
C4200 check[4] a_9237_2340# 0.0399f
C4201 x45.Q_N x75.Q 9.42e-21
C4202 a_12031_4775# a_12030_3213# 0.00237f
C4203 eob a_2265_2340# 9.03e-20
C4204 a_6760_4775# check[5] 0.00406f
C4205 a_7247_4775# a_7954_4801# 0.0968f
C4206 a_1520_2366# a_2060_2640# 0.139f
C4207 a_1207_2340# a_2061_2340# 0.0492f
C4208 D[2] a_11088_2366# 5.92e-20
C4209 a_2389_5648# eob 0.222f
C4210 a_9237_2340# a_11629_2340# 0.00176f
C4211 a_8696_2366# x63.Q_N 4.29e-21
C4212 check[4] a_11544_4775# 0.00302f
C4213 a_1227_4801# a_1592_5167# 4.45e-20
C4214 a_1682_4775# a_1415_4801# 6.99e-20
C4215 x4.X a_2289_4801# 0.167f
C4216 a_1061_4801# a_1926_5083# 0.00276f
C4217 a_4155_4086# a_4453_4386# 0.137f
C4218 a_3913_4112# a_4454_4086# 0.125f
C4219 sel_bit[1] x20.Q_N 3.57e-20
C4220 x5.X a_11089_4112# 0.00571f
C4221 check[2] x39.Q_N 0.0223f
C4222 x36.Q_N a_12737_3239# 0.0107f
C4223 a_4681_4801# x27.Q_N 5.04e-19
C4224 check[5] a_9238_4086# 6.24e-22
C4225 D[6] a_3912_2366# 0.00221f
C4226 a_11629_2340# a_12547_2366# 0.0708f
C4227 a_11088_2366# a_11969_2366# 0.00943f
C4228 a_11330_2340# a_11768_2366# 0.00276f
C4229 a_11833_2340# a_12345_2732# 6.69e-20
C4230 a_6606_4801# a_7182_4801# 2.46e-21
C4231 VDD a_11331_4086# 0.34f
C4232 x4.X a_4454_4086# 0.0468f
C4233 x5.A a_1227_4801# 6.32e-21
C4234 a_11857_4801# x36.Q_N 8.57e-20
C4235 check[1] a_8403_4801# 0.00119f
C4236 check[6] a_4452_2640# 0.0327f
C4237 x39.Q_N a_9151_3213# 3.3e-20
C4238 x4.X a_12548_4112# 0.00434f
C4239 a_4854_3213# a_7072_3239# 1.86e-21
C4240 a_4367_3213# a_6198_3239# 3.42e-20
C4241 a_6760_4775# a_7246_3213# 1.06e-20
C4242 a_7247_4775# a_6759_3213# 1.08e-22
C4243 a_4926_4296# x45.Q_N 1.43e-19
C4244 a_9237_4386# a_11089_4112# 9.95e-20
C4245 x42.Q_N a_9173_4112# 0.00139f
C4246 a_9442_4086# a_9578_4112# 0.07f
C4247 a_9238_4086# a_10776_4086# 2.98e-19
C4248 x36.Q_N a_11768_2366# 0.00473f
C4249 a_3452_3239# a_5561_3239# 1.03e-19
C4250 VDD a_6198_3239# 0.109f
C4251 check[6] a_4971_4801# 8.4e-20
C4252 a_6465_3213# a_6410_2366# 5.71e-21
C4253 a_4154_2340# a_4793_2366# 0.00316f
C4254 a_4452_2640# a_4592_2366# 0.00126f
C4255 a_3912_2366# a_5991_2340# 1.15e-20
C4256 x33.Q_N a_9710_4296# 5.71e-19
C4257 a_7072_3239# a_7181_3239# 0.00707f
C4258 check[5] a_9755_4801# 1.85e-20
C4259 eob a_3619_4801# 9.05e-22
C4260 eob a_2697_5083# 4.29e-19
C4261 x5.X a_6845_2340# 2.59e-20
C4262 x27.D a_3505_4086# 5.09e-21
C4263 check[3] a_10628_3239# 1.99e-20
C4264 check[0] a_6845_4386# 1.56e-19
C4265 VDD a_7049_2340# 0.304f
C4266 a_6546_2340# a_6780_2732# 0.00976f
C4267 a_5991_2340# a_6410_2366# 0.0397f
C4268 a_6304_2366# a_6982_2732# 0.00652f
C4269 a_7362_3239# a_7049_2340# 3.49e-20
C4270 a_11857_4801# a_11629_4386# 1.96e-20
C4271 a_11544_4775# a_11834_4086# 0.00268f
C4272 a_12031_4775# a_11630_4086# 0.00169f
C4273 a_11250_4775# x39.Q_N 2.02e-19
C4274 VDD a_1508_5167# 0.197f
C4275 check[1] a_7073_4801# 0.00111f
C4276 a_1227_4801# x27.D 4.24e-20
C4277 x5.X a_3600_4086# 1.13e-19
C4278 check[2] a_4926_4296# 2.18e-22
C4279 x5.A check[2] 0.00137f
C4280 x30.Q_N D[4] 0.005f
C4281 clk_sar x5.A 0.00356f
C4282 check[2] a_11769_4112# 3.17e-20
C4283 x48.Q a_3453_4801# 0.0505f
C4284 x5.X a_11767_4478# 4e-19
C4285 a_4155_4086# a_3899_3605# 1.7e-20
C4286 a_4453_4386# a_4073_3213# 0.0015f
C4287 a_3913_4112# a_4367_3213# 3.33e-20
C4288 a_4658_4086# a_3452_3239# 0.00195f
C4289 a_4454_4086# a_3618_3239# 6.04e-20
C4290 VDD a_1112_2340# 0.227f
C4291 VDD D[3] 0.221f
C4292 a_7763_2366# a_7561_2366# 3.67e-19
C4293 VDD x66.Q_N 0.0716f
C4294 a_8288_2340# a_8383_2340# 0.0968f
C4295 a_6780_2366# a_7185_2366# 2.46e-21
C4296 VDD a_3913_4112# 0.46f
C4297 x4.X a_3504_2340# 0.0105f
C4298 check[5] a_8998_4801# 2.15e-19
C4299 a_11543_3213# a_10982_3239# 3.79e-20
C4300 a_10628_3239# a_11493_3521# 0.00276f
C4301 a_11075_3605# a_11159_3605# 0.00972f
C4302 a_12030_3213# a_11856_3239# 0.197f
C4303 check[1] a_9710_4296# 3.53e-20
C4304 VDD a_11195_4112# 0.00996f
C4305 a_4794_4112# a_4925_2550# 1.72e-22
C4306 x5.X a_1682_4775# 0.00283f
C4307 a_11390_4801# check[3] 1.02e-20
C4308 x4.X a_4367_3213# 0.112f
C4309 x4.X a_6466_4775# 9.39e-19
C4310 a_6760_4775# x45.Q_N 9.66e-21
C4311 a_7073_4801# a_7050_4086# 2.59e-19
C4312 a_7247_4775# a_7318_4296# 2.97e-21
C4313 a_9710_4296# a_9954_4112# 0.00812f
C4314 x45.Q_N a_4680_3239# 1.74e-21
C4315 VDD x4.X 5.74f
C4316 x27.Q_N a_6978_4801# 1.15e-20
C4317 x4.X a_7362_3239# 5.65e-19
C4318 a_11856_3239# a_11628_2640# 1.11e-20
C4319 a_11543_3213# a_11833_2340# 0.00144f
C4320 a_12030_3213# a_11629_2340# 8.72e-19
C4321 a_10346_4801# check[4] 0.13f
C4322 x66.Q_N D[2] 2.25e-19
C4323 comparator_out a_6780_2732# 1.8e-19
C4324 a_9370_4801# x33.Q_N 4.03e-20
C4325 x4.X a_8939_4086# 0.00731f
C4326 a_8403_4801# a_8857_3213# 3.18e-21
C4327 a_8684_5167# a_8236_3239# 8.3e-21
C4328 check[2] x27.D 1.63e-20
C4329 a_6846_4086# x42.Q_N 2.42e-19
C4330 a_4855_4775# a_4453_4386# 6.17e-19
C4331 a_4368_4775# a_4454_4086# 4.63e-19
C4332 a_9442_4086# comparator_out 4.39e-21
C4333 a_8237_4801# a_8289_4086# 6.04e-19
C4334 check[0] a_7264_4394# 1.47e-20
C4335 D[3] a_11969_2366# 7.69e-20
C4336 a_2061_2340# a_3599_2340# 0.00116f
C4337 a_2265_2340# a_2401_2366# 0.07f
C4338 a_6010_3239# a_6291_3605# 0.155f
C4339 a_2060_2640# a_3912_2366# 1.9e-19
C4340 x4.X D[2] 4e-19
C4341 a_11330_2340# a_11833_2340# 0.00187f
C4342 a_11088_2366# a_12101_2550# 0.0633f
C4343 a_11628_2640# a_11629_2340# 0.781f
C4344 a_10775_2340# x63.Q_N 0.124f
C4345 x4.X x60.Q_N 0.00784f
C4346 a_2784_5996# a_2883_5674# 0.00134f
C4347 check[6] a_6759_3213# 8.24e-21
C4348 check[5] a_7561_2366# 5.2e-20
C4349 x4.X a_3807_4801# 2.51e-19
C4350 check[0] a_6984_2366# 3.17e-19
C4351 x5.X a_3452_3239# 3.24e-20
C4352 check[2] a_6760_4775# 1.3e-19
C4353 x4.X a_10983_4801# 2.36e-19
C4354 a_5845_4801# a_6011_4801# 0.751f
C4355 x36.Q_N a_11833_2340# 0.179f
C4356 sel_bit[0] a_1511_4112# 3.42e-19
C4357 a_3618_3239# a_4367_3213# 0.139f
C4358 a_3452_3239# a_4854_3213# 0.0492f
C4359 a_4073_3213# a_3899_3605# 0.205f
C4360 x54.Q_N a_4112_2648# 2.02e-20
C4361 a_4657_2340# a_4590_2732# 9.46e-19
C4362 a_3912_2366# a_5371_2366# 9.06e-21
C4363 a_4452_2640# a_4871_2648# 2.46e-19
C4364 a_6010_3239# a_6304_2366# 5.94e-19
C4365 a_6465_3213# a_5991_2340# 2.5e-19
C4366 a_8237_4801# a_10795_4801# 2.9e-21
C4367 a_8403_4801# a_10629_4801# 4e-20
C4368 VDD a_3618_3239# 0.291f
C4369 a_12147_4801# a_11966_4801# 4.11e-20
C4370 x39.Q_N a_11075_3605# 0.152f
C4371 a_12102_4296# a_11543_3213# 1.71e-19
C4372 a_11834_4086# a_12030_3213# 2.47e-19
C4373 check[2] a_9238_4086# 0.439f
C4374 x30.Q_N a_7072_3239# 0.00298f
C4375 sel_bit[0] a_1061_4801# 5.2e-20
C4376 x27.D a_4074_4775# 6.07e-19
C4377 check[5] a_6305_4112# 7.68e-22
C4378 VDD a_9464_3239# 0.18f
C4379 x20.Q_N x27.D 0.0032f
C4380 x48.Q a_4790_4801# 6.64e-20
C4381 check[4] a_11630_4086# 1.46e-21
C4382 a_5896_2340# a_6845_2340# 1.03e-19
C4383 VDD a_7186_4112# 0.0326f
C4384 a_9151_3213# a_9101_3521# 1.21e-20
C4385 a_8590_3239# a_8767_3605# 8.94e-19
C4386 a_8402_3239# a_8997_3239# 0.00118f
C4387 x20.Q_N a_2200_2366# 0.00397f
C4388 x42.Q_N a_8402_3239# 0.345f
C4389 a_9237_4386# a_9638_3213# 3.78e-19
C4390 a_9238_4086# a_9151_3213# 1.61e-19
C4391 x4.X a_8803_4112# 0.00332f
C4392 a_11630_4086# a_11629_2340# 1.55e-19
C4393 a_11629_4386# a_11833_2340# 1.26e-21
C4394 x39.Q_N a_11088_2366# 6.35e-20
C4395 a_897_4112# D[7] 3.76e-20
C4396 check[2] a_2579_4801# 1.13e-21
C4397 a_8384_4086# a_8697_4112# 0.272f
C4398 x5.X a_3900_5167# 1.6e-19
C4399 x30.Q_N a_6845_2340# 0.0463f
C4400 a_10156_4112# comparator_out 5.5e-20
C4401 a_4681_4801# a_5845_4801# 6.38e-20
C4402 a_4855_4775# a_6011_4801# 1.83e-19
C4403 a_4368_4775# a_4367_3213# 0.00121f
C4404 VDD a_9237_2340# 0.784f
C4405 x5.X a_11076_5167# 0.00471f
C4406 x4.X a_2198_2732# 9.81e-19
C4407 a_6844_2640# a_7561_2366# 0.00105f
C4408 check[3] a_11289_4394# 1.21e-21
C4409 D[1] a_11856_3239# 3.54e-20
C4410 a_8237_4801# a_9465_4801# 0.0334f
C4411 a_8403_4801# a_9639_4775# 0.0264f
C4412 a_8858_4775# a_9152_4775# 0.199f
C4413 x36.Q_N a_12102_4296# 1.85e-19
C4414 VDD a_4368_4775# 0.453f
C4415 a_6846_4086# a_6465_3213# 5.04e-19
C4416 a_7050_4086# a_6010_3239# 2.9e-19
C4417 a_6305_4112# a_7246_3213# 9.49e-19
C4418 a_6547_4086# a_6759_3213# 2.12e-19
C4419 comparator_out a_2777_2732# 8.11e-19
C4420 a_12031_4775# a_11966_4801# 4.2e-20
C4421 a_11857_4801# a_12147_4801# 0.0282f
C4422 a_5844_3239# a_6010_3239# 0.782f
C4423 a_5372_4112# a_5170_4112# 3.67e-19
C4424 a_9442_4086# a_8696_2366# 7.14e-22
C4425 a_9237_4386# a_9236_2640# 1.32e-20
C4426 a_9238_4086# a_8938_2340# 3.47e-21
C4427 VDD a_11544_4775# 0.449f
C4428 x77.Y a_4452_2640# 4.61e-20
C4429 check[4] D[1] 0.435f
C4430 a_9755_4801# a_9151_3213# 1.05e-20
C4431 check[6] comparator_out 0.0236f
C4432 VDD a_12547_2366# 0.109f
C4433 x48.Q a_4008_4801# 3.94e-19
C4434 x27.Q_N a_5561_3239# 0.00748f
C4435 a_2389_5648# sel_bit[0] 0.137f
C4436 check[3] comparator_out 0.0244f
C4437 D[1] a_11629_2340# 1.09e-20
C4438 a_9237_2340# x60.Q_N 1.07e-19
C4439 a_9441_2340# a_9709_2550# 0.205f
C4440 a_6845_4386# a_6304_2366# 1.93e-22
C4441 a_2883_5674# a_2463_4775# 6.31e-19
C4442 sel_bit[1] a_1508_5167# 5.1e-20
C4443 a_12548_4112# a_12030_3213# 2.07e-19
C4444 a_12031_4775# a_12737_3239# 4.94e-20
C4445 a_3453_4801# a_4318_5083# 0.00276f
C4446 a_3900_5167# a_3984_5167# 0.00972f
C4447 a_4855_4775# a_4681_4801# 0.197f
C4448 a_11331_4086# x39.Q_N 0.029f
C4449 x5.X a_8768_5167# 4.18e-19
C4450 a_11630_4086# a_11834_4086# 0.117f
C4451 a_11629_4386# a_12102_4296# 0.155f
C4452 x20.Q_N a_2579_4801# 0.00429f
C4453 a_2060_2640# D[6] 0.00655f
C4454 a_2265_2340# a_2777_2732# 6.69e-20
C4455 a_2061_2340# a_2979_2366# 0.0708f
C4456 D[2] a_12547_2366# 6.35e-19
C4457 a_7247_4775# a_9465_4801# 1.86e-21
C4458 D[3] a_12101_2550# 1.91e-20
C4459 x4.X a_11159_3605# 9.07e-19
C4460 VDD a_8897_4394# 0.00506f
C4461 check[1] a_6845_4386# 0.163f
C4462 a_3373_5674# a_3600_4086# 2.25e-20
C4463 a_11544_4775# a_10983_4801# 3.29e-21
C4464 a_11076_5167# a_11160_5167# 0.00972f
C4465 a_12031_4775# a_11857_4801# 0.197f
C4466 comparator_out a_8896_2648# 1.53e-19
C4467 a_10629_4801# a_11494_5083# 0.00276f
C4468 VDD a_7363_4801# 0.0101f
C4469 a_4658_4086# a_5372_4112# 6.99e-20
C4470 a_4155_4086# a_4593_4112# 0.00276f
C4471 a_4926_4296# a_5170_4478# 0.00972f
C4472 a_3913_4112# a_4794_4112# 0.00943f
C4473 a_4454_4086# a_5897_4086# 3.23e-19
C4474 check[2] a_5562_4801# 4.53e-20
C4475 a_8697_4112# a_9173_4478# 0.00133f
C4476 x33.Q_N a_8236_3239# 2.78e-19
C4477 a_8998_4801# a_9151_3213# 1.61e-20
C4478 a_9639_4775# a_9710_4296# 2.97e-21
C4479 a_9465_4801# a_9442_4086# 2.59e-19
C4480 a_9152_4775# x42.Q_N 9.8e-21
C4481 a_4214_4801# x77.Y 1.91e-20
C4482 sel_bit[0] a_3619_4801# 8.15e-19
C4483 a_3599_2340# a_4453_2340# 0.0492f
C4484 a_3912_2366# a_4452_2640# 0.139f
C4485 a_3258_5648# x4.X 3.57e-21
C4486 a_6010_3239# x72.Q_N 5.46e-21
C4487 a_4970_3239# a_4789_3239# 4.11e-20
C4488 a_7072_3239# a_7158_3605# 0.00976f
C4489 x4.X a_12101_2550# 0.00146f
C4490 sel_bit[1] x4.X 2.49e-19
C4491 x5.X D[0] 0.00133f
C4492 x4.X a_4794_4112# 0.00375f
C4493 a_4680_3239# a_4925_2550# 1.85e-20
C4494 a_4213_3239# a_3599_2340# 4.6e-20
C4495 a_6845_4386# a_7050_4086# 0.153f
C4496 a_6305_4112# x45.Q_N 0.093f
C4497 a_6845_4386# a_5844_3239# 6.5e-20
C4498 x5.X a_7159_5167# 1.05e-19
C4499 a_10629_4801# a_10681_4086# 6.04e-19
C4500 a_5371_2366# a_5991_2340# 8.26e-21
C4501 a_6011_4801# a_6400_4801# 0.0019f
C4502 a_6760_4775# a_6931_5083# 0.00652f
C4503 a_6466_4775# a_6606_4801# 0.07f
C4504 a_5845_4801# a_6978_4801# 2.56e-19
C4505 a_4452_2640# a_6410_2366# 2.44e-20
C4506 a_4367_3213# x75.Q_N 0.00553f
C4507 a_4854_3213# a_5088_3521# 0.00945f
C4508 a_3806_3239# a_4007_3239# 3.67e-19
C4509 a_4680_3239# a_4585_3239# 0.00276f
C4510 check[0] a_4767_5167# 1.92e-19
C4511 eob a_3600_4086# 4.72e-22
C4512 D[0] a_7181_3239# 9.28e-21
C4513 a_1511_4112# a_1520_2366# 7.01e-19
C4514 a_9465_4801# a_9574_4801# 0.00707f
C4515 VDD x75.Q_N 0.0719f
C4516 x20.Q_N a_2479_2648# 0.00136f
C4517 VDD a_6606_4801# 0.0332f
C4518 x39.Q_N x66.Q_N 3.91e-19
C4519 a_3619_4801# check[6] 5.82e-21
C4520 x39.Q_N a_11195_4112# 0.0451f
C4521 VDD a_12030_3213# 0.568f
C4522 a_11834_4086# a_12346_4478# 6.69e-20
C4523 a_11331_4086# a_11769_4112# 0.00276f
C4524 a_11630_4086# a_12548_4112# 0.0708f
C4525 a_11089_4112# a_11970_4112# 0.00943f
C4526 check[1] a_8236_3239# 0.0444f
C4527 eob a_1682_4775# 0.0484f
C4528 check[5] a_8403_4801# 0.162f
C4529 a_6546_2340# a_6780_2366# 0.00707f
C4530 a_6304_2366# a_6984_2366# 3.73e-19
C4531 a_6844_2640# a_8288_2340# 6.58e-19
C4532 check[1] a_7264_4394# 6.91e-21
C4533 a_9151_3213# a_9573_3239# 2.87e-21
C4534 a_9638_3213# a_9754_3239# 0.0397f
C4535 a_2389_5648# a_2788_5674# 2.97e-20
C4536 a_8997_3239# a_9369_3239# 3.34e-19
C4537 check[4] a_11966_4801# 9.01e-21
C4538 a_10795_4801# check[3] 8.42e-19
C4539 comparator_out a_1520_2366# 0.00311f
C4540 x42.Q_N a_10628_3239# 1.47e-19
C4541 a_1682_4775# x4.A 0.00205f
C4542 VDD a_10346_4801# 0.192f
C4543 x5.X a_5372_4112# 9.6e-19
C4544 x42.Q_N a_9369_3239# 0.00401f
C4545 check[2] a_6305_4112# 1.74e-20
C4546 x4.X x39.Q_N 0.253f
C4547 x30.Q_N a_9236_2640# 1.21e-20
C4548 x48.Q a_3505_4086# 0.0868f
C4549 a_5372_4112# a_4854_3213# 2.07e-19
C4550 check[3] a_11194_2366# 1.29e-19
C4551 a_2463_4775# a_2289_4801# 0.197f
C4552 a_1508_5167# a_1592_5167# 0.00972f
C4553 x5.X x27.Q_N 0.00103f
C4554 VDD a_11628_2640# 0.269f
C4555 x27.Q_N a_4854_3213# 0.0125f
C4556 x27.Q_N a_6292_5167# 5.48e-20
C4557 VDD a_2784_5996# 0.00533f
C4558 check[4] a_8697_4112# 3.77e-22
C4559 x4.X a_4388_2732# 4.32e-19
C4560 a_8383_2340# a_9172_2732# 7.71e-20
C4561 a_8696_2366# a_8896_2648# 0.00185f
C4562 VDD a_5897_4086# 0.189f
C4563 x5.X x36.Q_N 0.00489f
C4564 a_10628_3239# a_10680_2340# 4.5e-19
C4565 a_12030_3213# D[2] 0.00376f
C4566 x4.X a_6930_3521# 9.99e-19
C4567 a_9754_3239# a_9236_2640# 5.05e-21
C4568 a_9152_4775# a_9873_5083# 0.00185f
C4569 a_8684_5167# x33.Q_N 1.74e-20
C4570 x4.X a_6505_4394# 1.75e-19
C4571 a_5844_3239# a_8236_3239# 0.00176f
C4572 comparator_out a_4871_2648# 6.94e-19
C4573 x27.Q_N a_5169_2366# 0.00224f
C4574 x45.Q_N a_6605_3239# 0.031f
C4575 a_5844_3239# a_6977_3239# 2.56e-19
C4576 x48.Q a_1227_4801# 5.44e-21
C4577 x4.X x75.Q 8.71e-19
C4578 a_6845_4386# a_7764_4112# 0.162f
C4579 a_6305_4112# a_6781_4112# 2.87e-21
C4580 a_7050_4086# a_7264_4394# 0.0104f
C4581 a_6846_4086# a_7562_4478# 0.0018f
C4582 check[0] a_6291_3605# 7.4e-20
C4583 check[4] a_9709_2550# 0.00101f
C4584 a_7073_4801# check[5] 6.72e-20
C4585 a_1207_2340# a_2533_2550# 4.7e-22
C4586 a_1520_2366# a_2265_2340# 0.199f
C4587 a_1762_2340# a_2061_2340# 0.0334f
C4588 D[2] a_11628_2640# 0.00729f
C4589 a_12737_3239# a_11629_2340# 4.83e-19
C4590 a_12030_3213# a_11969_2366# 1.2e-20
C4591 a_9236_2640# x63.Q_N 1.48e-19
C4592 eob a_3452_3239# 3.51e-19
C4593 check[4] a_11857_4801# 4.17e-20
C4594 a_1227_4801# a_2147_5083# 1.09e-19
C4595 a_1682_4775# a_1926_5083# 0.0104f
C4596 a_4155_4086# a_4658_4086# 0.00187f
C4597 a_3600_4086# x48.Q_N 0.124f
C4598 a_4453_4386# a_4454_4086# 0.75f
C4599 a_3913_4112# a_4926_4296# 0.0633f
C4600 check[0] a_6304_2366# 0.00297f
C4601 x5.X a_11629_4386# 0.00326f
C4602 a_12346_4478# a_12548_4112# 8.94e-19
C4603 a_2979_2366# a_4453_2340# 3.65e-21
C4604 D[6] a_4452_2640# 1.85e-19
C4605 a_11629_2340# a_11768_2366# 2.56e-19
C4606 a_12101_2550# a_12547_2366# 0.0367f
C4607 a_11628_2640# a_11969_2366# 0.00118f
C4608 a_12147_4801# a_12102_4296# 1.9e-20
C4609 VDD a_11630_4086# 0.809f
C4610 x4.X a_4926_4296# 0.0211f
C4611 check[6] a_4657_2340# 6.83e-20
C4612 check[1] check[0] 0.0116f
C4613 a_4367_3213# a_4970_3239# 0.0552f
C4614 a_7073_4801# a_7246_3213# 4.82e-21
C4615 a_7247_4775# a_7072_3239# 1.33e-23
C4616 x4.X a_11769_4112# 6.71e-19
C4617 check[2] x48.Q 0.0879f
C4618 x33.Q_N a_8791_3239# 6.75e-20
C4619 x42.Q_N a_9578_4112# 0.00172f
C4620 a_9238_4086# a_11331_4086# 1.67e-21
C4621 a_9710_4296# a_10776_4086# 7.98e-21
C4622 x36.Q_N a_12345_2366# 0.00224f
C4623 a_1976_4775# a_3170_4801# 6.04e-19
C4624 a_1508_5167# x27.D 4.66e-22
C4625 x77.Y comparator_out 0.00119f
C4626 VDD a_4970_3239# 0.00144f
C4627 check[6] a_6710_5083# 2.57e-21
C4628 a_8236_3239# a_8857_3213# 0.117f
C4629 a_4453_2340# a_4793_2366# 6.04e-20
C4630 a_4657_2340# a_4592_2366# 9.75e-19
C4631 a_4452_2640# a_5991_2340# 3.67e-19
C4632 x72.Q_N a_8236_3239# 2.94e-19
C4633 x5.X a_10345_3239# 0.00125f
C4634 x42.Q_N a_6759_3213# 3.3e-20
C4635 a_11630_4086# D[2] 3.53e-19
C4636 x20.Q_N a_1207_2340# 0.144f
C4637 x30.Q_N D[0] 3.29e-19
C4638 x33.Q_N a_9172_2366# 9.42e-19
C4639 check[0] a_3877_5674# 0.00787f
C4640 x5.X a_1976_4775# 0.00314f
C4641 VDD D[1] 0.3f
C4642 VDD x57.Q_N 0.0716f
C4643 check[0] a_7050_4086# 1.2e-19
C4644 check[0] a_5844_3239# 0.051f
C4645 D[5] a_6984_2366# 8.02e-20
C4646 a_6844_2640# a_6982_2732# 1.09e-19
C4647 a_6304_2366# a_7263_2648# 1.21e-20
C4648 a_6546_2340# a_6410_2366# 0.0282f
C4649 a_8236_3239# a_8383_2340# 8.35e-19
C4650 D[0] a_9754_3239# 1.61e-20
C4651 D[7] a_1996_2366# 1.53e-19
C4652 a_11544_4775# x39.Q_N 9.93e-21
C4653 a_12031_4775# a_12102_4296# 2.97e-21
C4654 a_11857_4801# a_11834_4086# 2.59e-19
C4655 a_3505_4086# a_3599_2340# 1.57e-20
C4656 VDD a_2463_4775# 0.704f
C4657 x20.Q_N a_4018_2366# 1.31e-20
C4658 x4.X x27.D 0.00252f
C4659 x5.X a_4155_4086# 7.39e-20
C4660 x5.X a_12048_4394# 1.32e-19
C4661 x48.Q a_4074_4775# 0.00395f
C4662 a_3913_4112# a_4680_3239# 2.16e-19
C4663 a_4453_4386# a_4367_3213# 5.72e-19
C4664 a_3600_4086# a_3806_3239# 2.44e-19
C4665 check[3] a_10775_2340# 2.56e-20
C4666 a_4855_4775# a_5561_3239# 4.94e-20
C4667 x48.Q x20.Q_N 0.0441f
C4668 a_10794_3239# a_11714_3521# 1.09e-19
C4669 a_11249_3213# a_11493_3521# 0.0104f
C4670 VDD a_4453_4386# 0.593f
C4671 check[5] a_9370_4801# 7.95e-20
C4672 VDD a_12346_4478# 0.0042f
C4673 a_9238_4086# D[3] 1.26e-20
C4674 comparator_out a_3912_2366# 0.00684f
C4675 a_11762_4801# check[3] 7.79e-21
C4676 x27.Q_N a_5896_2340# 1.79e-19
C4677 check[5] a_6010_3239# 2.24e-21
C4678 x4.X a_4680_3239# 0.0059f
C4679 x4.X a_6760_4775# 0.104f
C4680 check[2] a_8403_4801# 4.08e-19
C4681 a_2463_4775# a_3807_4801# 8.26e-21
C4682 a_10681_4086# a_10776_4086# 0.0968f
C4683 a_9173_4112# a_9578_4112# 2.46e-21
C4684 a_6199_4801# comparator_out 1.97e-20
C4685 check[1] a_9172_2366# 1.35e-19
C4686 a_1822_4801# a_2194_4801# 3.34e-19
C4687 x4.X a_6504_2648# 0.00102f
C4688 a_8802_2366# a_9172_2366# 4.11e-20
C4689 x27.Q_N x30.Q_N 2.3e-20
C4690 x4.X a_9101_3521# 2.91e-19
C4691 a_11856_3239# a_11833_2340# 1.03e-19
C4692 a_12030_3213# a_12101_2550# 1.66e-21
C4693 x4.X a_9238_4086# 0.0468f
C4694 a_8403_4801# a_9151_3213# 2.05e-21
C4695 a_8684_5167# a_8857_3213# 3.52e-21
C4696 a_8858_4775# a_8683_3605# 1.33e-23
C4697 check[0] D[5] 0.228f
C4698 a_7318_4296# x42.Q_N 8.46e-20
C4699 a_4855_4775# a_4658_4086# 4.44e-19
C4700 a_4368_4775# a_4926_4296# 2.85e-19
C4701 x42.Q_N comparator_out 0.00133f
C4702 a_3619_4801# x77.Y 5.26e-21
C4703 a_6010_3239# a_7246_3213# 0.0264f
C4704 a_6465_3213# a_6759_3213# 0.199f
C4705 a_2533_2550# a_3599_2340# 7.98e-21
C4706 a_2061_2340# a_4154_2340# 6.38e-20
C4707 a_2265_2340# a_3912_2366# 9.6e-21
C4708 check[3] a_11089_4112# 0.0033f
C4709 a_11330_2340# x63.Q_N 9.58e-21
C4710 a_11628_2640# a_12101_2550# 0.145f
C4711 a_11629_2340# a_11833_2340# 0.117f
C4712 a_2883_5674# a_2969_6040# 0.0136f
C4713 comparator_out a_10680_2340# 7.8e-19
C4714 a_5372_4112# a_5992_4086# 8.26e-21
C4715 x4.X a_2579_4801# 0.0171f
C4716 check[2] a_7073_4801# 4.32e-20
C4717 x5.X a_5845_4801# 0.27f
C4718 x4.X a_9755_4801# 0.00557f
C4719 x36.Q_N x63.Q_N 4.08e-19
C4720 a_3452_3239# a_3806_3239# 0.0662f
C4721 a_3618_3239# a_4680_3239# 0.137f
C4722 a_5845_4801# a_6292_5167# 0.15f
C4723 a_6011_4801# a_6466_4775# 0.153f
C4724 a_3899_3605# a_4367_3213# 0.0632f
C4725 sel_bit[0] a_3600_4086# 3.59e-19
C4726 check[0] a_3453_4801# 0.00279f
C4727 a_4452_2640# a_5371_2366# 0.159f
C4728 a_4657_2340# a_4871_2648# 0.0104f
C4729 a_4453_2340# a_5169_2732# 0.0018f
C4730 a_6010_3239# a_6844_2640# 4.04e-20
C4731 a_6759_3213# a_5991_2340# 9.06e-19
C4732 a_6465_3213# a_6546_2340# 4.18e-20
C4733 a_6291_3605# a_6304_2366# 1.71e-19
C4734 x5.X a_12147_4801# 2.09e-19
C4735 VDD a_3899_3605# 0.182f
C4736 VDD a_6011_4801# 0.593f
C4737 check[1] a_9377_4112# 3.4e-20
C4738 check[6] a_6845_2340# 3.11e-22
C4739 a_12102_4296# a_11856_3239# 2.37e-20
C4740 x39.Q_N a_12030_3213# 0.144f
C4741 check[1] x33.Q_N 0.0011f
C4742 VDD a_11966_4801# 7.87e-19
C4743 x5.X a_8384_4086# 0.0202f
C4744 x33.Q_N a_8802_2366# 0.0102f
C4745 check[2] a_9710_4296# 0.00118f
C4746 sel_bit[0] a_1682_4775# 7.55e-20
C4747 a_7954_4801# a_6846_4086# 6.67e-19
C4748 check[5] a_6845_4386# 0.0306f
C4749 x27.D a_4368_4775# 0.00307f
C4750 VDD a_8767_3605# 0.0042f
C4751 D[7] a_1626_2366# 0.00202f
C4752 x75.Q_N x75.Q 2.81e-20
C4753 a_8236_3239# a_10794_3239# 2.9e-21
C4754 a_8402_3239# a_10628_3239# 4e-20
C4755 a_5991_2340# a_6546_2340# 0.197f
C4756 a_9151_3213# a_9550_3605# 0.00133f
C4757 a_8236_3239# a_9872_3521# 1.25e-19
C4758 a_8402_3239# a_9369_3239# 0.00126f
C4759 a_8683_3605# a_8997_3239# 0.0258f
C4760 VDD a_8697_4112# 0.448f
C4761 x42.Q_N a_8683_3605# 0.152f
C4762 a_9442_4086# a_9638_3213# 2.47e-19
C4763 a_9710_4296# a_9151_3213# 1.71e-19
C4764 x20.Q_N a_3599_2340# 3.36e-19
C4765 x4.X a_9954_4478# 9.15e-19
C4766 a_12102_4296# a_11629_2340# 6.08e-21
C4767 x39.Q_N a_11628_2640# 4.61e-20
C4768 x30.Q_N a_7317_2550# 0.181f
C4769 a_8289_4086# x42.Q_N 0.18f
C4770 a_8384_4086# a_9237_4386# 0.0264f
C4771 a_8697_4112# a_8939_4086# 0.124f
C4772 x5.X a_4855_4775# 0.00928f
C4773 x4.X a_8998_4801# 7.25e-19
C4774 a_4855_4775# a_6292_5167# 7.98e-21
C4775 a_4855_4775# a_4854_3213# 0.00237f
C4776 VDD a_12737_3239# 0.189f
C4777 VDD a_9709_2550# 0.172f
C4778 check[1] a_6304_2366# 1.25e-21
C4779 x5.X a_12031_4775# 0.00483f
C4780 x4.X a_2479_2648# 2.86e-19
C4781 a_6845_2340# a_8896_2648# 4.06e-20
C4782 a_8858_4775# a_9465_4801# 0.00187f
C4783 a_8237_4801# a_8768_5167# 0.0018f
C4784 a_8403_4801# a_8591_4801# 0.162f
C4785 a_8684_5167# a_9639_4775# 4.7e-22
C4786 VDD a_4681_4801# 0.346f
C4787 a_6846_4086# a_6759_3213# 1.61e-19
C4788 x45.Q_N a_6010_3239# 0.346f
C4789 a_6845_4386# a_7246_3213# 3.78e-19
C4790 comparator_out D[6] 0.00566f
C4791 comparator_out a_6465_3213# 4.84e-19
C4792 a_5844_3239# a_6291_3605# 0.15f
C4793 x42.Q_N a_8696_2366# 6.41e-20
C4794 a_9238_4086# a_9237_2340# 1.55e-19
C4795 a_9237_4386# a_9441_2340# 1.26e-21
C4796 x4.X a_5562_4801# 0.00612f
C4797 x77.Y a_4657_2340# 1.11e-19
C4798 VDD a_11857_4801# 0.343f
C4799 x48.Q a_5170_4478# 5.12e-20
C4800 a_5897_4086# x75.Q 0.00123f
C4801 x4.X a_12738_4801# 0.00262f
C4802 VDD a_11768_2366# 6.2e-19
C4803 check[1] a_8802_2366# 0.00244f
C4804 x48.Q a_5089_5083# 1.17e-19
C4805 a_12737_3239# D[2] 0.0747f
C4806 a_8696_2366# a_10680_2340# 7.33e-21
C4807 a_8383_2340# a_9172_2366# 4.2e-20
C4808 a_2853_5648# a_1511_4112# 6.37e-19
C4809 a_6846_4086# a_6546_2340# 3.47e-21
C4810 a_7050_4086# a_6304_2366# 7.14e-22
C4811 a_6845_4386# a_6844_2640# 1.32e-20
C4812 check[1] a_9954_4112# 5.77e-22
C4813 comparator_out a_5991_2340# 0.00445f
C4814 a_5844_3239# a_6304_2366# 1.89e-19
C4815 a_8237_4801# D[0] 1.99e-20
C4816 check[5] a_8236_3239# 0.00639f
C4817 sel_bit[1] a_2463_4775# 5.3e-20
C4818 x5.X a_9173_4478# 3.15e-19
C4819 check[2] a_10681_4086# 0.126f
C4820 check[0] a_4453_2340# 0.00712f
C4821 a_3619_4801# a_4539_5083# 1.09e-19
C4822 a_4074_4775# a_4318_5083# 0.0104f
C4823 a_11834_4086# a_12102_4296# 0.205f
C4824 a_11630_4086# x39.Q_N 0.00117f
C4825 x5.X a_7182_4801# 5.34e-20
C4826 a_2265_2340# D[6] 1.59e-19
C4827 a_2533_2550# a_2979_2366# 0.0367f
C4828 a_6760_4775# a_7363_4801# 0.0552f
C4829 VDD a_9375_4478# 0.0163f
C4830 x4.X a_9573_3239# 1.05e-19
C4831 check[1] a_7050_4086# 7.72e-19
C4832 check[1] a_5844_3239# 2.07e-22
C4833 comparator_out a_9374_2732# 9.52e-19
C4834 a_11250_4775# a_11494_5083# 0.0104f
C4835 a_10795_4801# a_11715_5083# 1.09e-19
C4836 a_10156_4112# a_9638_3213# 2.07e-19
C4837 VDD a_9102_5083# 0.00984f
C4838 a_4454_4086# a_4593_4112# 2.56e-19
C4839 a_4453_4386# a_4794_4112# 0.00118f
C4840 a_4155_4086# a_5992_4086# 1.86e-21
C4841 check[5] a_6984_2366# 9.43e-20
C4842 a_8697_4112# a_8803_4112# 0.051f
C4843 a_8939_4086# a_9375_4478# 0.00412f
C4844 a_9237_4386# a_9173_4478# 2.13e-19
C4845 a_9238_4086# a_8897_4394# 1.25e-19
C4846 x33.Q_N a_8857_3213# 5.46e-19
C4847 VDD a_1996_2732# 0.00483f
C4848 check[6] a_3452_3239# 1.79e-20
C4849 a_3599_2340# a_4925_2550# 4.7e-22
C4850 sel_bit[0] a_3900_5167# 2.68e-19
C4851 a_7246_3213# a_8236_3239# 0.00116f
C4852 a_6759_3213# a_8402_3239# 1.98e-19
C4853 a_4154_2340# a_4453_2340# 0.0334f
C4854 a_3912_2366# a_4657_2340# 0.199f
C4855 a_11768_2366# a_11969_2366# 3.34e-19
C4856 a_6759_3213# a_7480_3521# 0.00185f
C4857 a_621_4112# x3.A 0.129f
C4858 reset a_897_4112# 0.00119f
C4859 eob a_1976_4775# 0.0525f
C4860 VDD a_897_4112# 0.414f
C4861 x4.X a_6305_4112# 0.11f
C4862 x39.Q_N D[1] 3.4e-19
C4863 a_6846_4086# a_7318_4296# 0.15f
C4864 a_6845_4386# x45.Q_N 0.00117f
C4865 a_6846_4086# comparator_out 3.21e-20
C4866 a_7050_4086# a_5844_3239# 0.00195f
C4867 x33.Q_N a_8383_2340# 0.142f
C4868 check[0] a_4019_4112# 1.03e-20
C4869 x5.X a_6400_4801# 2.84e-19
C4870 eob D[7] 2.52e-20
C4871 D[5] a_6304_2366# 8.64e-19
C4872 a_1112_2340# a_1207_2340# 0.0968f
C4873 a_5845_4801# x30.Q_N 2.24e-19
C4874 a_6760_4775# a_6606_4801# 0.00943f
C4875 a_6292_5167# a_6400_4801# 0.00812f
C4876 a_7073_4801# a_6931_5083# 0.00412f
C4877 a_6466_4775# a_6978_4801# 9.75e-19
C4878 a_7247_4775# a_7159_5167# 7.71e-20
C4879 a_4680_3239# x75.Q_N 9.58e-21
C4880 a_2389_5648# a_2853_5648# 0.202f
C4881 a_1511_4112# a_2060_2640# 0.00164f
C4882 x33.Q_N a_10629_4801# 7.17e-19
C4883 VDD a_6978_4801# 0.00445f
C4884 x20.Q_N a_2979_2366# 0.00156f
C4885 a_4368_4775# a_5562_4801# 6.04e-19
C4886 a_3900_5167# check[6] 1.4e-21
C4887 VDD a_10982_3239# 0.109f
C4888 a_11630_4086# a_11769_4112# 2.56e-19
C4889 a_12102_4296# a_12548_4112# 0.0367f
C4890 a_11629_4386# a_11970_4112# 0.00118f
C4891 x5.X check[4] 0.167f
C4892 a_8857_3213# a_8802_2366# 5.71e-21
C4893 check[1] x72.Q_N 4.68e-20
C4894 a_6546_2340# a_7185_2366# 0.00316f
C4895 a_6844_2640# a_6984_2366# 0.00126f
C4896 a_6304_2366# a_8383_2340# 7.3e-21
C4897 check[5] a_8684_5167# 0.00124f
C4898 x4.X a_1207_2340# 0.117f
C4899 a_9464_3239# a_9573_3239# 0.00707f
C4900 check[1] a_7764_4112# 0.165f
C4901 check[2] a_2993_5674# 0.0021f
C4902 comparator_out a_2060_2640# 0.113f
C4903 a_11076_5167# check[3] 5.35e-19
C4904 a_11544_4775# a_12738_4801# 6.04e-19
C4905 x5.X a_11629_2340# 4.23e-20
C4906 check[2] a_6845_4386# 1.41e-20
C4907 x42.Q_N x69.Q_N 3.92e-19
C4908 x30.Q_N a_9441_2340# 9.31e-21
C4909 x48.Q a_3913_4112# 8.72e-19
C4910 a_4454_4086# a_5561_3239# 4.72e-19
C4911 a_5845_4801# a_5992_4086# 0.00159f
C4912 a_1976_4775# a_1926_5083# 1.21e-20
C4913 VDD a_3648_5972# 0.0123f
C4914 VDD a_11833_2340# 0.304f
C4915 check[1] a_8383_2340# 0.0126f
C4916 VDD a_2969_6040# 0.00654f
C4917 a_8938_2340# a_9172_2732# 0.00976f
C4918 a_8383_2340# a_8802_2366# 0.0397f
C4919 a_8696_2366# a_9374_2732# 0.00652f
C4920 a_10346_4801# a_9238_4086# 6.67e-19
C4921 check[4] a_9237_4386# 0.028f
C4922 x4.X a_4018_2366# 3.78e-20
C4923 VDD a_4593_4112# 0.00494f
C4924 a_9754_3239# a_9441_2340# 3.49e-20
C4925 x4.X a_6605_3239# 0.00267f
C4926 a_2853_5648# a_3619_4801# 3.82e-19
C4927 a_9639_4775# x33.Q_N 0.126f
C4928 check[1] a_3453_4801# 9.29e-20
C4929 a_5844_3239# D[5] 5.19e-19
C4930 x45.Q_N a_8236_3239# 1.49e-19
C4931 comparator_out a_5371_2366# 0.155f
C4932 x4.X a_6983_4478# 0.00114f
C4933 comparator_out a_8402_3239# 0.147f
C4934 x45.Q_N a_6977_3239# 0.00399f
C4935 x48.Q x4.X 0.188f
C4936 a_5844_3239# x72.Q_N 1.07e-19
C4937 a_6305_4112# a_7186_4112# 0.00943f
C4938 a_6547_4086# a_6985_4112# 0.00276f
C4939 a_6846_4086# a_8289_4086# 3.23e-19
C4940 a_7318_4296# a_7562_4478# 0.00972f
C4941 a_7050_4086# a_7764_4112# 6.99e-20
C4942 a_10155_2366# a_9953_2366# 3.67e-19
C4943 a_1520_2366# x51.Q_N 0.00553f
C4944 a_2060_2640# a_2265_2340# 0.153f
C4945 a_10680_2340# a_10775_2340# 0.0968f
C4946 a_9172_2366# a_9577_2366# 2.46e-21
C4947 D[2] a_11833_2340# 4.68e-20
C4948 x4.X a_8288_2340# 0.00317f
C4949 a_1227_4801# a_1822_4801# 0.00118f
C4950 a_4155_4086# x48.Q_N 9.58e-21
C4951 a_4454_4086# a_4658_4086# 0.117f
C4952 a_4453_4386# a_4926_4296# 0.155f
C4953 check[0] a_6844_2640# 2.7e-19
C4954 x5.X a_11834_4086# 3.65e-19
C4955 a_3600_4086# x77.Y 1.36e-19
C4956 a_6010_3239# a_7953_3239# 1e-20
C4957 D[6] a_4657_2340# 2.71e-19
C4958 a_11833_2340# a_11969_2366# 0.07f
C4959 x30.Q_N a_7182_4801# 7.02e-20
C4960 check[2] a_8236_3239# 6.24e-22
C4961 VDD a_12102_4296# 0.317f
C4962 comparator_out a_11564_2732# 1.8e-19
C4963 a_4680_3239# a_4970_3239# 0.0282f
C4964 a_4854_3213# a_4789_3239# 4.2e-20
C4965 x4.X a_12346_4112# 6.38e-19
C4966 x33.Q_N a_7763_2366# 1.34e-20
C4967 x33.Q_N a_10794_3239# 3.79e-20
C4968 VDD a_4112_2648# 0.00555f
C4969 a_2463_4775# x27.D 0.00431f
C4970 a_9238_4086# a_11630_4086# 1.37e-19
C4971 x48.Q a_3618_3239# 2.51e-19
C4972 a_8697_4112# x39.Q_N 1.05e-20
C4973 a_4367_3213# a_5561_3239# 6.04e-19
C4974 VDD a_6709_3521# 0.00984f
C4975 a_4452_2640# a_6546_2340# 4.11e-20
C4976 a_4925_2550# a_4793_2366# 0.0258f
C4977 a_4453_2340# a_6304_2366# 3.16e-19
C4978 a_8236_3239# a_9151_3213# 0.126f
C4979 a_8402_3239# a_8683_3605# 0.155f
C4980 VDD a_5170_4112# 1.14e-19
C4981 VDD a_5561_3239# 0.19f
C4982 x20.Q_N a_1762_2340# 0.162f
C4983 x39.Q_N a_12737_3239# 3.23e-19
C4984 x4.X a_8403_4801# 0.005f
C4985 x33.Q_N a_9577_2366# 0.0403f
C4986 x5.X a_2289_4801# 0.00166f
C4987 a_12738_4801# a_12030_3213# 3.19e-20
C4988 check[3] a_11543_3213# 1.04e-19
C4989 check[0] x45.Q_N 0.0173f
C4990 a_6844_2640# a_7263_2648# 2.46e-19
C4991 a_6304_2366# a_7763_2366# 5.76e-21
C4992 a_7049_2340# a_6982_2732# 9.46e-19
C4993 x57.Q_N a_6504_2648# 2.02e-20
C4994 D[7] a_2401_2366# 4.38e-19
C4995 a_8402_3239# a_8696_2366# 5.94e-19
C4996 a_8857_3213# a_8383_2340# 2.5e-19
C4997 a_6400_4801# x30.Q_N 3.71e-20
C4998 VDD a_1415_4801# 0.12f
C4999 a_3913_4112# a_3599_2340# 5.05e-21
C5000 a_9238_4086# D[1] 3.36e-19
C5001 x33.Q_N a_11184_4801# 3.99e-20
C5002 x5.X a_4454_4086# 0.258f
C5003 sel_bit[1] a_897_4112# 1.46e-20
C5004 check[6] a_5372_4112# 0.00256f
C5005 x5.X a_12548_4112# 5.39e-19
C5006 x48.Q a_4368_4775# 0.0017f
C5007 a_4454_4086# a_4854_3213# 7.94e-19
C5008 a_4658_4086# a_4367_3213# 0.0014f
C5009 check[3] a_11330_2340# 1.32e-19
C5010 x27.Q_N check[6] 0.934f
C5011 x77.Y a_3452_3239# 0.51f
C5012 clk_sar a_621_4112# 9.27e-21
C5013 a_8288_2340# a_9237_2340# 1.03e-19
C5014 x4.X a_3599_2340# 0.117f
C5015 VDD a_4658_4086# 0.489f
C5016 a_10794_3239# a_11389_3239# 0.00118f
C5017 a_10982_3239# a_11159_3605# 8.94e-19
C5018 a_11543_3213# a_11493_3521# 1.21e-20
C5019 VDD a_1062_5674# 0.23f
C5020 check[5] x33.Q_N 3.66e-21
C5021 VDD a_11565_4112# 3.47e-19
C5022 comparator_out a_4452_2640# 0.109f
C5023 x36.Q_N check[3] 1.17f
C5024 x27.Q_N a_4592_2366# 0.00474f
C5025 x4.X a_7073_4801# 0.00316f
C5026 x4.X a_3983_3605# 0.00103f
C5027 check[2] a_8684_5167# 1.92e-19
C5028 a_2463_4775# a_2579_4801# 0.0397f
C5029 a_1976_4775# a_2398_4801# 2.87e-21
C5030 check[2] check[0] 0.872f
C5031 check[1] a_9577_2366# 4.4e-19
C5032 a_1822_4801# x20.Q_N 1.36e-19
C5033 a_9236_2640# a_9953_2366# 0.00105f
C5034 a_5845_4801# a_8237_4801# 0.00176f
C5035 x4.X a_6982_2732# 9.81e-19
C5036 x4.X a_9550_3605# 4.4e-19
C5037 a_6846_4086# D[4] 1.26e-20
C5038 comparator_out a_7561_2732# 8.23e-19
C5039 comparator_out a_10628_3239# 0.148f
C5040 a_3600_4086# a_4113_4394# 0.00945f
C5041 x4.X a_9710_4296# 0.021f
C5042 check[5] a_6304_2366# 1.15e-20
C5043 a_9465_4801# a_8402_3239# 6.75e-21
C5044 a_4681_4801# a_4926_4296# 3.59e-20
C5045 a_8237_4801# a_8384_4086# 0.00159f
C5046 a_3900_5167# x77.Y 7.98e-21
C5047 check[0] a_6781_4112# 9.63e-22
C5048 a_1520_2366# x54.Q_N 5.89e-21
C5049 a_2061_2340# a_4453_2340# 0.00176f
C5050 a_3648_5972# a_3258_5648# 8.72e-19
C5051 sel_bit[0] a_1976_4775# 1.72e-19
C5052 a_6291_3605# a_7246_3213# 4.7e-22
C5053 a_6010_3239# a_6198_3239# 0.163f
C5054 a_6465_3213# a_7072_3239# 0.00187f
C5055 a_11629_2340# x63.Q_N 1.07e-19
C5056 a_11833_2340# a_12101_2550# 0.205f
C5057 check[3] a_11629_4386# 0.138f
C5058 a_12738_4801# a_11630_4086# 6.67e-19
C5059 a_2883_5674# a_3373_5674# 4.47e-19
C5060 a_12031_4775# a_11970_4112# 1.79e-20
C5061 VDD a_3170_4801# 0.212f
C5062 a_3452_3239# a_3912_2366# 1.89e-19
C5063 a_3618_3239# a_3599_2340# 3.73e-19
C5064 check[1] check[5] 0.343f
C5065 a_5897_4086# a_6305_4112# 4.37e-19
C5066 a_4593_4112# a_4794_4112# 3.34e-19
C5067 x33.Q_N a_6844_2640# 0.00104f
C5068 x5.X a_6466_4775# 0.00314f
C5069 VDD a_1996_2366# 4.24e-19
C5070 a_5845_4801# a_7247_4775# 0.0492f
C5071 a_6011_4801# a_6760_4775# 0.139f
C5072 a_6466_4775# a_6292_5167# 0.205f
C5073 a_4073_3213# a_3806_3239# 6.99e-20
C5074 a_4367_3213# a_4854_3213# 0.273f
C5075 a_3618_3239# a_3983_3605# 4.45e-20
C5076 a_3452_3239# a_4317_3521# 0.00276f
C5077 a_7953_3239# a_8236_3239# 8.18e-19
C5078 check[0] a_4074_4775# 5.86e-19
C5079 a_4453_2340# D[5] 0.338f
C5080 a_4925_2550# a_5169_2732# 0.00972f
C5081 a_4657_2340# a_5371_2366# 6.99e-20
C5082 a_7246_3213# a_6304_2366# 8.4e-19
C5083 a_6010_3239# a_7049_2340# 0.00154f
C5084 a_6465_3213# a_6845_2340# 0.00199f
C5085 a_6759_3213# a_6546_2340# 2.17e-19
C5086 VDD x5.X 2.74f
C5087 a_9152_4775# a_10795_4801# 8.44e-20
C5088 a_9639_4775# a_10629_4801# 0.00116f
C5089 VDD a_4854_3213# 0.572f
C5090 VDD a_6292_5167# 0.317f
C5091 a_10776_4086# a_11389_3239# 1.16e-20
C5092 x39.Q_N a_10982_3239# 7.52e-20
C5093 x5.X a_8939_4086# 0.00115f
C5094 VDD a_5169_2366# 4e-20
C5095 x27.D a_4681_4801# 2.31e-21
C5096 check[5] a_5844_3239# 1.81e-20
C5097 check[1] a_7246_3213# 0.00245f
C5098 eob a_2883_5674# 6.72e-19
C5099 a_6304_2366# a_6844_2640# 0.139f
C5100 a_5991_2340# a_6845_2340# 0.0492f
C5101 a_9464_3239# a_9550_3605# 0.00976f
C5102 a_7362_3239# a_7181_3239# 4.11e-20
C5103 a_8402_3239# x69.Q_N 4.5e-21
C5104 VDD a_9237_4386# 0.59f
C5105 x5.X D[2] 0.0046f
C5106 x42.Q_N a_9638_3213# 0.144f
C5107 a_9710_4296# a_9464_3239# 2.37e-20
C5108 x4.X a_10681_4086# 0.0036f
C5109 x20.Q_N a_4154_2340# 2.93e-20
C5110 x39.Q_N a_11833_2340# 1.11e-19
C5111 x5.X a_3807_4801# 5.48e-19
C5112 a_6985_4112# x42.Q_N 1.96e-20
C5113 a_8939_4086# a_9237_4386# 0.137f
C5114 a_8697_4112# a_9238_4086# 0.125f
C5115 x4.X a_9370_4801# 5.55e-19
C5116 x5.A a_897_4112# 5.71e-20
C5117 check[1] a_6844_2640# 7.55e-20
C5118 a_7763_2366# a_8383_2340# 8.26e-21
C5119 x5.X a_10983_4801# 0.00551f
C5120 a_6844_2640# a_8802_2366# 1.71e-20
C5121 x4.X a_2979_2366# 4.09e-19
C5122 x4.X a_6010_3239# 0.0446f
C5123 D[1] a_9573_3239# 9.28e-21
C5124 a_8403_4801# a_7363_4801# 4.14e-20
C5125 a_8858_4775# a_8768_5167# 6.69e-20
C5126 a_8684_5167# a_8591_4801# 0.0367f
C5127 a_9152_4775# a_9465_4801# 0.124f
C5128 check[3] a_12048_4394# 5.14e-21
C5129 VDD a_3984_5167# 0.0046f
C5130 x45.Q_N a_6291_3605# 0.152f
C5131 a_7050_4086# a_7246_3213# 2.47e-19
C5132 a_7318_4296# a_6759_3213# 1.71e-19
C5133 a_5844_3239# a_7246_3213# 0.0492f
C5134 comparator_out a_6759_3213# 7.49e-19
C5135 a_9710_4296# a_9237_2340# 6.08e-21
C5136 x42.Q_N a_9236_2640# 4.61e-20
C5137 VDD a_11160_5167# 0.0042f
C5138 a_10795_4801# a_10628_3239# 9.04e-19
C5139 a_10629_4801# a_10794_3239# 8.16e-19
C5140 x77.Y a_5088_3521# 8.16e-21
C5141 a_9236_2640# a_10680_2340# 6.83e-19
C5142 a_8696_2366# a_9376_2366# 3.73e-19
C5143 a_8938_2340# a_9172_2366# 0.00707f
C5144 a_2853_5648# a_3600_4086# 2.47e-19
C5145 a_11389_3239# a_11761_3239# 3.34e-19
C5146 a_6845_4386# a_7049_2340# 1.26e-21
C5147 x45.Q_N a_6304_2366# 6.37e-20
C5148 a_6846_4086# a_6845_2340# 1.55e-19
C5149 a_5844_3239# a_6844_2640# 6.01e-20
C5150 comparator_out a_6546_2340# 0.00104f
C5151 x27.Q_N a_6780_2366# 9.28e-21
C5152 x20.Q_N a_4389_4478# 3.31e-21
C5153 check[2] a_9377_4112# 6.45e-20
C5154 check[5] x72.Q_N 0.00322f
C5155 a_4368_4775# a_4318_5083# 1.21e-20
C5156 a_3807_4801# a_3984_5167# 8.94e-19
C5157 a_3619_4801# a_4214_4801# 0.00118f
C5158 check[5] a_7764_4112# 0.00263f
C5159 check[2] x33.Q_N 0.0366f
C5160 a_12102_4296# x39.Q_N 0.00244f
C5161 x5.X a_9323_5083# 5.14e-19
C5162 a_10775_2340# a_11564_2732# 7.71e-20
C5163 a_11088_2366# a_11288_2648# 0.00185f
C5164 x4.X a_9172_2732# 4.32e-19
C5165 a_7073_4801# a_7363_4801# 0.0282f
C5166 a_7247_4775# a_7182_4801# 4.2e-20
C5167 x4.X a_11714_3521# 9.99e-19
C5168 check[1] x45.Q_N 0.00102f
C5169 VDD a_9656_4394# 0.00984f
C5170 a_1061_4801# a_1511_4112# 0.00351f
C5171 comparator_out a_9655_2648# 7e-19
C5172 a_10795_4801# a_11390_4801# 0.00118f
C5173 a_3452_3239# D[6] 2.82e-19
C5174 a_10983_4801# a_11160_5167# 8.94e-19
C5175 a_11544_4775# a_11494_5083# 1.21e-20
C5176 a_1062_5674# sel_bit[1] 0.039f
C5177 VDD a_9551_5167# 0.00371f
C5178 check[5] a_8383_2340# 3.32e-21
C5179 a_4454_4086# a_5992_4086# 2.98e-19
C5180 a_4658_4086# a_4794_4112# 0.07f
C5181 a_4453_4386# a_6305_4112# 8.96e-20
C5182 a_1511_4112# comparator_out 8.67e-19
C5183 a_9238_4086# a_9375_4478# 0.00907f
C5184 x42.Q_N a_7562_4112# 2.85e-21
C5185 x33.Q_N a_9151_3213# 0.00498f
C5186 VDD a_1626_2366# 0.00785f
C5187 check[6] a_5845_4801# 0.416f
C5188 a_5562_4801# a_6011_4801# 4.06e-19
C5189 x27.Q_N x77.Y 0.00357f
C5190 a_6759_3213# a_8683_3605# 4.38e-20
C5191 a_7072_3239# a_8402_3239# 3.9e-20
C5192 a_4452_2640# a_4657_2340# 0.153f
C5193 a_3912_2366# x54.Q_N 0.00553f
C5194 a_8403_4801# a_10346_4801# 9.65e-21
C5195 a_8237_4801# check[4] 8.28e-20
C5196 a_7246_3213# x72.Q_N 0.124f
C5197 eob a_2289_4801# 0.0076f
C5198 a_7764_4112# a_7246_3213# 2.07e-19
C5199 x4.X a_6845_4386# 0.048f
C5200 check[3] a_12147_4801# 2.59e-19
C5201 a_9578_4112# a_8696_2366# 1.26e-20
C5202 a_7050_4086# x45.Q_N 0.00116f
C5203 x45.Q_N a_5844_3239# 0.0434f
C5204 x33.Q_N a_8938_2340# 0.16f
C5205 a_5561_3239# x75.Q 0.0955f
C5206 VDD a_5896_2340# 0.189f
C5207 D[5] a_6844_2640# 4.09e-20
C5208 a_5371_2366# a_6845_2340# 3.65e-21
C5209 D[7] a_1520_2366# 0.00164f
C5210 a_10629_4801# a_10776_4086# 0.00159f
C5211 a_6760_4775# a_6978_4801# 3.73e-19
C5212 a_7073_4801# a_6606_4801# 0.00316f
C5213 a_6466_4775# x30.Q_N 1.17e-19
C5214 check[0] a_5089_5083# 4.43e-19
C5215 check[2] check[1] 2.29f
C5216 D[0] a_8997_3239# 1.6e-19
C5217 a_1511_4112# a_2265_2340# 0.00119f
C5218 x33.Q_N a_11250_4775# 4.4e-20
C5219 x42.Q_N D[0] 3.91e-19
C5220 VDD x30.Q_N 0.444f
C5221 a_3258_5648# a_3170_4801# 0.00133f
C5222 a_2389_5648# a_1511_4112# 0.00132f
C5223 sel_bit[1] a_3170_4801# 1.85e-19
C5224 x30.Q_N a_7362_3239# 0.00342f
C5225 check[2] a_9954_4112# 1.28e-19
C5226 a_12738_4801# a_12737_3239# 9.85e-20
C5227 x48.Q a_2463_4775# 9e-19
C5228 a_4855_4775# check[6] 0.0103f
C5229 check[1] a_9151_3213# 1.78e-20
C5230 a_11834_4086# a_11970_4112# 0.07f
C5231 VDD a_9754_3239# 4.88e-19
C5232 x39.Q_N a_11565_4112# 0.0014f
C5233 a_6844_2640# a_8383_2340# 3.42e-19
C5234 a_7049_2340# a_6984_2366# 9.75e-19
C5235 a_6845_2340# a_7185_2366# 6.04e-20
C5236 a_10628_3239# a_11249_3213# 0.117f
C5237 check[5] a_9639_4775# 2.58e-20
C5238 x4.X a_1762_2340# 0.00671f
C5239 x69.Q_N a_10628_3239# 2.94e-19
C5240 check[1] a_6781_4112# 1.37e-20
C5241 a_12345_2366# VSS 8.87e-19
C5242 a_11969_2366# VSS 0.182f
C5243 a_11768_2366# VSS 0.00989f
C5244 a_11564_2366# VSS 0.00207f
C5245 a_12547_2366# VSS 0.0962f
C5246 a_12345_2732# VSS 3.33e-19
C5247 a_12047_2648# VSS 4.04e-19
C5248 a_11194_2366# VSS 0.158f
C5249 a_11766_2732# VSS 0.0011f
C5250 a_11564_2732# VSS 1.58e-19
C5251 a_11288_2648# VSS 1.45e-19
C5252 a_9953_2366# VSS 6.96e-19
C5253 x63.Q_N VSS 0.1f
C5254 a_12101_2550# VSS 0.262f
C5255 a_11833_2340# VSS 0.29f
C5256 a_11629_2340# VSS 0.606f
C5257 a_11628_2640# VSS 0.419f
C5258 a_11330_2340# VSS 0.251f
C5259 a_11088_2366# VSS 0.387f
C5260 a_10775_2340# VSS 0.458f
C5261 a_9577_2366# VSS 0.18f
C5262 a_9376_2366# VSS 0.00923f
C5263 a_9172_2366# VSS 0.00192f
C5264 a_10680_2340# VSS 0.225f
C5265 D[3] VSS 0.365f
C5266 a_10155_2366# VSS 0.0926f
C5267 a_8802_2366# VSS 0.157f
C5268 a_9374_2732# VSS 3.84e-19
C5269 a_7561_2366# VSS 6.96e-19
C5270 x60.Q_N VSS 0.1f
C5271 a_9709_2550# VSS 0.256f
C5272 a_9441_2340# VSS 0.286f
C5273 a_9237_2340# VSS 0.512f
C5274 a_9236_2640# VSS 0.4f
C5275 a_8938_2340# VSS 0.249f
C5276 a_8696_2366# VSS 0.385f
C5277 a_8383_2340# VSS 0.456f
C5278 a_7185_2366# VSS 0.18f
C5279 a_6984_2366# VSS 0.00923f
C5280 a_6780_2366# VSS 0.00192f
C5281 a_8288_2340# VSS 0.225f
C5282 D[4] VSS 0.365f
C5283 a_7763_2366# VSS 0.0926f
C5284 a_6410_2366# VSS 0.157f
C5285 a_6982_2732# VSS 3.84e-19
C5286 a_5169_2366# VSS 6.96e-19
C5287 x57.Q_N VSS 0.1f
C5288 a_7317_2550# VSS 0.256f
C5289 a_7049_2340# VSS 0.286f
C5290 a_6845_2340# VSS 0.513f
C5291 a_6844_2640# VSS 0.4f
C5292 a_6546_2340# VSS 0.249f
C5293 a_6304_2366# VSS 0.385f
C5294 a_5991_2340# VSS 0.456f
C5295 a_4793_2366# VSS 0.18f
C5296 a_4592_2366# VSS 0.00923f
C5297 a_4388_2366# VSS 0.00192f
C5298 a_5896_2340# VSS 0.225f
C5299 D[5] VSS 0.393f
C5300 a_5371_2366# VSS 0.0926f
C5301 a_4018_2366# VSS 0.157f
C5302 a_4590_2732# VSS 3.84e-19
C5303 a_2777_2366# VSS 0.00168f
C5304 x54.Q_N VSS 0.1f
C5305 a_4925_2550# VSS 0.256f
C5306 a_4657_2340# VSS 0.286f
C5307 a_4453_2340# VSS 0.513f
C5308 a_4452_2640# VSS 0.4f
C5309 a_4154_2340# VSS 0.249f
C5310 a_3912_2366# VSS 0.385f
C5311 a_3599_2340# VSS 0.458f
C5312 a_2401_2366# VSS 0.18f
C5313 a_2200_2366# VSS 0.00923f
C5314 a_1996_2366# VSS 0.00192f
C5315 a_3504_2340# VSS 0.226f
C5316 D[6] VSS 0.604f
C5317 a_2979_2366# VSS 0.0988f
C5318 a_1626_2366# VSS 0.157f
C5319 a_2198_2732# VSS 3.84e-19
C5320 x51.Q_N VSS 0.1f
C5321 a_2533_2550# VSS 0.263f
C5322 a_2265_2340# VSS 0.289f
C5323 a_2061_2340# VSS 0.517f
C5324 a_2060_2640# VSS 0.527f
C5325 a_1762_2340# VSS 0.25f
C5326 a_1520_2366# VSS 0.387f
C5327 a_1207_2340# VSS 0.469f
C5328 D[7] VSS 0.536f
C5329 a_1112_2340# VSS 0.247f
C5330 a_11965_3239# VSS 0.00208f
C5331 a_12146_3239# VSS 0.159f
C5332 D[2] VSS 1.11f
C5333 a_12737_3239# VSS 0.252f
C5334 x66.Q_N VSS 0.102f
C5335 a_12264_3521# VSS 3.9e-19
C5336 a_11761_3239# VSS 0.00967f
C5337 a_11183_3239# VSS 0.00168f
C5338 a_11389_3239# VSS 0.181f
C5339 a_11942_3605# VSS 2.25e-19
C5340 a_11714_3521# VSS 0.00103f
C5341 a_11493_3521# VSS 2.34e-19
C5342 a_9573_3239# VSS 0.00192f
C5343 a_9754_3239# VSS 0.157f
C5344 a_10982_3239# VSS 0.0988f
C5345 a_11856_3239# VSS 0.25f
C5346 a_12030_3213# VSS 0.463f
C5347 a_11543_3213# VSS 0.389f
C5348 a_11075_3605# VSS 0.259f
C5349 a_11249_3213# VSS 0.281f
C5350 a_10794_3239# VSS 0.519f
C5351 a_10628_3239# VSS 0.509f
C5352 D[1] VSS 0.467f
C5353 a_10345_3239# VSS 0.222f
C5354 x69.Q_N VSS 0.1f
C5355 a_9369_3239# VSS 0.00923f
C5356 a_8791_3239# VSS 0.00168f
C5357 a_8997_3239# VSS 0.18f
C5358 a_9322_3521# VSS 3.84e-19
C5359 a_7181_3239# VSS 0.00192f
C5360 a_7362_3239# VSS 0.157f
C5361 a_8590_3239# VSS 0.0988f
C5362 a_9464_3239# VSS 0.246f
C5363 a_9638_3213# VSS 0.446f
C5364 a_9151_3213# VSS 0.38f
C5365 a_8683_3605# VSS 0.258f
C5366 a_8857_3213# VSS 0.28f
C5367 a_8402_3239# VSS 0.519f
C5368 a_8236_3239# VSS 0.506f
C5369 D[0] VSS 0.471f
C5370 a_7953_3239# VSS 0.222f
C5371 x72.Q_N VSS 0.1f
C5372 a_6977_3239# VSS 0.00923f
C5373 a_6399_3239# VSS 0.00168f
C5374 a_6605_3239# VSS 0.18f
C5375 a_6930_3521# VSS 3.84e-19
C5376 a_4789_3239# VSS 0.00196f
C5377 a_4970_3239# VSS 0.157f
C5378 a_6198_3239# VSS 0.0988f
C5379 a_7072_3239# VSS 0.246f
C5380 a_7246_3213# VSS 0.446f
C5381 a_6759_3213# VSS 0.38f
C5382 a_6291_3605# VSS 0.258f
C5383 a_6465_3213# VSS 0.28f
C5384 a_6010_3239# VSS 0.519f
C5385 comparator_out VSS 11.6f
C5386 a_5844_3239# VSS 0.506f
C5387 x75.Q VSS 0.239f
C5388 a_5561_3239# VSS 0.222f
C5389 x75.Q_N VSS 0.1f
C5390 a_4585_3239# VSS 0.00943f
C5391 a_4007_3239# VSS 0.00202f
C5392 a_4213_3239# VSS 0.181f
C5393 a_4538_3521# VSS 3.84e-19
C5394 a_3806_3239# VSS 0.263f
C5395 a_4680_3239# VSS 0.246f
C5396 a_4854_3213# VSS 0.446f
C5397 a_4367_3213# VSS 0.379f
C5398 a_3899_3605# VSS 0.261f
C5399 a_4073_3213# VSS 0.28f
C5400 a_3618_3239# VSS 0.751f
C5401 a_3452_3239# VSS 0.888f
C5402 x77.Y VSS 1.02f
C5403 a_12346_4112# VSS 0.00226f
C5404 a_11970_4112# VSS 0.183f
C5405 a_11769_4112# VSS 0.00991f
C5406 a_11565_4112# VSS 0.00168f
C5407 a_12548_4112# VSS 0.102f
C5408 a_12346_4478# VSS 3.33e-19
C5409 a_12048_4394# VSS 3.91e-19
C5410 a_11195_4112# VSS 0.148f
C5411 a_11767_4478# VSS 0.00107f
C5412 a_11565_4478# VSS 1.58e-19
C5413 a_11289_4394# VSS 1.48e-19
C5414 a_9954_4112# VSS 0.00168f
C5415 x39.Q_N VSS 1.23f
C5416 a_12102_4296# VSS 0.261f
C5417 a_11834_4086# VSS 0.279f
C5418 a_11630_4086# VSS 0.588f
C5419 a_11629_4386# VSS 0.537f
C5420 a_11331_4086# VSS 0.238f
C5421 a_11089_4112# VSS 0.318f
C5422 a_10776_4086# VSS 0.425f
C5423 a_9578_4112# VSS 0.18f
C5424 a_9377_4112# VSS 0.00923f
C5425 a_9173_4112# VSS 0.00155f
C5426 a_10681_4086# VSS 0.207f
C5427 a_10156_4112# VSS 0.0984f
C5428 a_8803_4112# VSS 0.147f
C5429 a_9375_4478# VSS 3.84e-19
C5430 a_7562_4112# VSS 0.00168f
C5431 x42.Q_N VSS 1.22f
C5432 a_9710_4296# VSS 0.255f
C5433 a_9442_4086# VSS 0.275f
C5434 a_9238_4086# VSS 0.484f
C5435 a_9237_4386# VSS 0.515f
C5436 a_8939_4086# VSS 0.236f
C5437 a_8697_4112# VSS 0.316f
C5438 a_8384_4086# VSS 0.423f
C5439 a_7186_4112# VSS 0.18f
C5440 a_6985_4112# VSS 0.00923f
C5441 a_6781_4112# VSS 0.00157f
C5442 a_8289_4086# VSS 0.205f
C5443 a_7764_4112# VSS 0.0984f
C5444 a_6411_4112# VSS 0.147f
C5445 a_6983_4478# VSS 3.84e-19
C5446 a_5170_4112# VSS 0.00168f
C5447 x45.Q_N VSS 1.22f
C5448 a_7318_4296# VSS 0.255f
C5449 a_7050_4086# VSS 0.275f
C5450 a_6846_4086# VSS 0.484f
C5451 a_6845_4386# VSS 0.515f
C5452 a_6547_4086# VSS 0.236f
C5453 a_6305_4112# VSS 0.316f
C5454 a_5992_4086# VSS 0.423f
C5455 a_4794_4112# VSS 0.18f
C5456 a_4593_4112# VSS 0.00923f
C5457 a_4389_4112# VSS 0.00192f
C5458 a_5897_4086# VSS 0.211f
C5459 a_5372_4112# VSS 0.0984f
C5460 a_4019_4112# VSS 0.157f
C5461 a_4591_4478# VSS 3.84e-19
C5462 x48.Q_N VSS 0.1f
C5463 a_4926_4296# VSS 0.255f
C5464 a_4658_4086# VSS 0.275f
C5465 a_4454_4086# VSS 0.486f
C5466 a_4453_4386# VSS 0.515f
C5467 a_4155_4086# VSS 0.243f
C5468 a_3913_4112# VSS 0.373f
C5469 a_3600_4086# VSS 0.443f
C5470 a_3505_4086# VSS 0.225f
C5471 a_1511_4112# VSS 2.05f
C5472 x4.A VSS 0.932f
C5473 a_897_4112# VSS 0.522f
C5474 x3.A VSS 0.206f
C5475 a_621_4112# VSS 0.284f
C5476 reset VSS 0.247f
C5477 a_11966_4801# VSS 0.00215f
C5478 a_12147_4801# VSS 0.161f
C5479 check[3] VSS 1.3f
C5480 a_12738_4801# VSS 0.255f
C5481 x36.Q_N VSS 1.28f
C5482 a_12265_5083# VSS 5.88e-19
C5483 a_11762_4801# VSS 0.00989f
C5484 a_11184_4801# VSS 0.00168f
C5485 a_11390_4801# VSS 0.181f
C5486 a_11943_5167# VSS 2.29e-19
C5487 a_11715_5083# VSS 0.00114f
C5488 a_11494_5083# VSS 2.58e-19
C5489 a_9574_4801# VSS 0.00192f
C5490 a_9755_4801# VSS 0.157f
C5491 a_10983_4801# VSS 0.0987f
C5492 a_11857_4801# VSS 0.25f
C5493 a_12031_4775# VSS 0.46f
C5494 a_11544_4775# VSS 0.386f
C5495 a_11076_5167# VSS 0.257f
C5496 a_11250_4775# VSS 0.279f
C5497 a_10795_4801# VSS 0.517f
C5498 a_10629_4801# VSS 0.488f
C5499 check[4] VSS 0.823f
C5500 a_10346_4801# VSS 0.21f
C5501 x33.Q_N VSS 1.25f
C5502 a_9370_4801# VSS 0.00923f
C5503 a_8792_4801# VSS 0.00168f
C5504 a_8998_4801# VSS 0.18f
C5505 a_9323_5083# VSS 3.84e-19
C5506 a_7182_4801# VSS 0.00192f
C5507 a_7363_4801# VSS 0.157f
C5508 a_8591_4801# VSS 0.0987f
C5509 a_9465_4801# VSS 0.244f
C5510 a_9639_4775# VSS 0.435f
C5511 a_9152_4775# VSS 0.373f
C5512 a_8684_5167# VSS 0.257f
C5513 a_8858_4775# VSS 0.276f
C5514 a_8403_4801# VSS 0.515f
C5515 a_8237_4801# VSS 0.484f
C5516 check[5] VSS 0.83f
C5517 a_7954_4801# VSS 0.207f
C5518 x30.Q_N VSS 1.26f
C5519 a_6978_4801# VSS 0.00923f
C5520 a_6400_4801# VSS 0.00168f
C5521 a_6606_4801# VSS 0.18f
C5522 a_6931_5083# VSS 3.84e-19
C5523 a_4790_4801# VSS 0.00192f
C5524 a_4971_4801# VSS 0.157f
C5525 a_6199_4801# VSS 0.0987f
C5526 a_7073_4801# VSS 0.244f
C5527 a_7247_4775# VSS 0.435f
C5528 a_6760_4775# VSS 0.373f
C5529 a_6292_5167# VSS 0.257f
C5530 a_6466_4775# VSS 0.276f
C5531 a_6011_4801# VSS 0.515f
C5532 a_5845_4801# VSS 0.484f
C5533 check[6] VSS 0.845f
C5534 a_5562_4801# VSS 0.207f
C5535 x27.Q_N VSS 1.25f
C5536 a_4586_4801# VSS 0.00923f
C5537 a_4008_4801# VSS 0.00168f
C5538 a_4214_4801# VSS 0.18f
C5539 a_4539_5083# VSS 3.84e-19
C5540 a_2398_4801# VSS 0.00192f
C5541 a_2579_4801# VSS 0.157f
C5542 a_3807_4801# VSS 0.0987f
C5543 a_4681_4801# VSS 0.244f
C5544 a_4855_4775# VSS 0.435f
C5545 a_4368_4775# VSS 0.373f
C5546 a_3900_5167# VSS 0.257f
C5547 a_4074_4775# VSS 0.275f
C5548 a_3619_4801# VSS 0.513f
C5549 a_3453_4801# VSS 0.481f
C5550 x27.D VSS 0.243f
C5551 a_3170_4801# VSS 0.22f
C5552 x20.Q_N VSS 1.25f
C5553 a_2194_4801# VSS 0.00923f
C5554 a_1616_4801# VSS 0.00168f
C5555 a_1822_4801# VSS 0.18f
C5556 a_2147_5083# VSS 3.84e-19
C5557 a_1415_4801# VSS 0.0987f
C5558 a_2289_4801# VSS 0.242f
C5559 a_2463_4775# VSS 0.429f
C5560 a_1976_4775# VSS 0.37f
C5561 a_1508_5167# VSS 0.256f
C5562 x4.X VSS 16.6f
C5563 a_1682_4775# VSS 0.275f
C5564 a_1227_4801# VSS 0.516f
C5565 a_1061_4801# VSS 0.541f
C5566 a_3877_5674# VSS 0.00437f
C5567 a_3671_5674# VSS 0.00563f
C5568 a_2993_5674# VSS 0.00182f
C5569 a_2788_5674# VSS 0.00372f
C5570 a_3373_5674# VSS 0.115f
C5571 a_3258_5648# VSS 0.229f
C5572 check[0] VSS 2.45f
C5573 x48.Q VSS 0.615f
C5574 sel_bit[1] VSS 1.15f
C5575 a_2883_5674# VSS 0.185f
C5576 a_2784_5996# VSS 2.03e-19
C5577 eob VSS 2.1f
C5578 x5.X VSS 12.6f
C5579 check[1] VSS 2.3f
C5580 a_2853_5648# VSS 0.373f
C5581 sel_bit[0] VSS 0.54f
C5582 check[2] VSS 4.17f
C5583 a_2389_5648# VSS 0.48f
C5584 a_1338_5674# VSS 0.322f
C5585 x5.A VSS 0.226f
C5586 a_1062_5674# VSS 0.274f
C5587 clk_sar VSS 0.214f
C5588 VDD VSS 0.105p
.ends

