* NGSPICE file created from hgu_sw_cap.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_L7T3GD a_n33_n130# a_15_n42# a_n73_n42# VSUBS
X0 a_15_n42# a_n33_n130# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt hgu_sw_cap SW CTOP delay_signal
XXM14 SW delay_signal x2/CBOT VSUBS sky130_fd_pr__nfet_01v8_L7T3GD
.ends

