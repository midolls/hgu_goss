* NGSPICE file created from hgu_cdac_cap_64.ext - technology: sky130A

.subckt hgu_cdac_cap_64 CTOP CBOT SUB
C0 CTOP CBOT 0.323p
C1 CTOP SUB 27.6f
C2 CBOT SUB 16.8f
.ends

