magic
tech sky130A
magscale 1 2
timestamp 1699184817
<< nwell >>
rect 6688 3774 7508 3812
rect 6688 3772 7592 3774
rect 6602 3168 7592 3772
rect 6602 3138 7254 3168
rect 6690 2894 7004 3138
rect 6690 2842 7010 2894
rect 6693 2840 7010 2842
rect 6693 2591 6754 2840
rect 6713 -1799 6992 -1241
rect 6221 -1860 6992 -1799
rect 6188 -2464 6992 -1860
rect 6221 -2467 6992 -2464
<< pwell >>
rect 24 -606 13310 1820
<< psubdiff >>
rect 76 1702 194 1722
rect 76 1645 103 1702
rect 169 1645 194 1702
rect 76 1623 194 1645
<< nsubdiff >>
rect 7015 3666 7101 3692
rect 7015 3632 7041 3666
rect 7075 3632 7101 3666
rect 7015 3606 7101 3632
rect 7004 3494 7090 3520
rect 7004 3460 7030 3494
rect 7064 3460 7090 3494
rect 7004 3434 7090 3460
rect 7004 3302 7090 3328
rect 7004 3268 7030 3302
rect 7064 3268 7090 3302
rect 7004 3242 7090 3268
rect 6412 -1914 6498 -1888
rect 6412 -1948 6438 -1914
rect 6472 -1948 6498 -1914
rect 6412 -1974 6498 -1948
rect 6412 -2110 6498 -2084
rect 6412 -2144 6438 -2110
rect 6472 -2144 6498 -2110
rect 6412 -2170 6498 -2144
rect 6412 -2285 6498 -2259
rect 6412 -2319 6438 -2285
rect 6472 -2319 6498 -2285
rect 6412 -2345 6498 -2319
<< psubdiffcont >>
rect 103 1645 169 1702
<< nsubdiffcont >>
rect 7041 3632 7075 3666
rect 7030 3460 7064 3494
rect 7030 3268 7064 3302
rect 6438 -1948 6472 -1914
rect 6438 -2144 6472 -2110
rect 6438 -2319 6472 -2285
<< locali >>
rect 7015 3666 7101 3692
rect 7015 3632 7041 3666
rect 7075 3632 7101 3666
rect 7015 3606 7101 3632
rect 7004 3494 7090 3520
rect 7004 3460 7030 3494
rect 7064 3460 7090 3494
rect 7004 3434 7090 3460
rect 7004 3302 7090 3328
rect 7004 3268 7030 3302
rect 7064 3268 7090 3302
rect 7004 3242 7090 3268
rect 77 1702 195 1721
rect 77 1645 103 1702
rect 169 1645 195 1702
rect 77 1622 195 1645
rect 6412 -1914 6498 -1888
rect 6412 -1948 6438 -1914
rect 6472 -1948 6498 -1914
rect 6412 -1974 6498 -1948
rect 6412 -2110 6498 -2084
rect 6412 -2144 6438 -2110
rect 6472 -2144 6498 -2110
rect 6412 -2170 6498 -2144
rect 6412 -2285 6498 -2259
rect 6412 -2319 6438 -2285
rect 6472 -2319 6498 -2285
rect 6412 -2345 6498 -2319
<< viali >>
rect 7041 3632 7075 3666
rect 7030 3460 7064 3494
rect 7030 3268 7064 3302
rect 105 1649 163 1700
rect 6438 -1948 6472 -1914
rect 6438 -2144 6472 -2110
rect 6438 -2319 6472 -2285
<< metal1 >>
rect 7011 3673 7101 3689
rect 7011 3621 7030 3673
rect 7082 3621 7101 3673
rect 7011 3605 7101 3621
rect 7000 3501 7090 3517
rect 7000 3449 7019 3501
rect 7071 3449 7090 3501
rect 7000 3433 7090 3449
rect 7000 3309 7090 3325
rect 7000 3257 7019 3309
rect 7071 3257 7090 3309
rect 7000 3241 7090 3257
rect 0 2774 138 2808
rect 6709 2774 6847 2808
rect 37 2391 705 2438
rect 6685 2386 6755 2438
rect 13382 2389 13492 2435
rect 88 1700 186 1715
rect 88 1644 105 1700
rect 165 1644 186 1700
rect 88 1625 186 1644
rect 2489 1047 2547 1072
rect 283 1019 2547 1047
rect 4915 991 4973 1070
rect 283 963 4973 991
rect 5771 935 5829 1072
rect 283 907 5829 935
rect 9198 879 9256 1070
rect 283 851 9256 879
rect 11624 823 11682 1072
rect 283 795 11682 823
rect 12480 767 12538 1064
rect 283 739 12538 767
rect 283 685 12574 711
rect 283 684 12504 685
rect 283 632 900 684
rect 952 677 12504 684
rect 952 674 7609 677
rect 952 632 5800 674
rect 283 622 5800 632
rect 5853 624 7609 674
rect 7661 624 12504 677
rect 5853 622 12504 624
rect 283 621 12504 622
rect 12568 621 12574 685
rect 283 599 12574 621
rect 283 543 10975 571
rect 283 487 8549 515
rect 283 431 7693 459
rect 283 375 4266 403
rect 283 319 1840 347
rect 283 263 984 291
rect 925 258 984 263
rect 1782 254 1840 319
rect 4208 251 4266 375
rect 7635 249 7693 431
rect 8491 245 8549 487
rect 10917 254 10975 543
rect 24 -1114 78 -1068
rect 6708 -1117 6770 -1068
rect 13446 -1070 13492 2389
rect 13419 -1117 13492 -1070
rect 6617 -1487 6755 -1453
rect 13326 -1487 13464 -1453
rect 6412 -1903 6502 -1887
rect 6412 -1955 6431 -1903
rect 6483 -1955 6502 -1903
rect 6412 -1971 6502 -1955
rect 6412 -2099 6502 -2083
rect 6412 -2151 6431 -2099
rect 6483 -2151 6502 -2099
rect 6412 -2167 6502 -2151
rect 6412 -2274 6502 -2258
rect 6412 -2326 6431 -2274
rect 6483 -2326 6502 -2274
rect 6412 -2342 6502 -2326
<< via1 >>
rect 7030 3666 7082 3673
rect 7030 3632 7041 3666
rect 7041 3632 7075 3666
rect 7075 3632 7082 3666
rect 7030 3621 7082 3632
rect 7019 3494 7071 3501
rect 7019 3460 7030 3494
rect 7030 3460 7064 3494
rect 7064 3460 7071 3494
rect 7019 3449 7071 3460
rect 7019 3302 7071 3309
rect 7019 3268 7030 3302
rect 7030 3268 7064 3302
rect 7064 3268 7071 3302
rect 7019 3257 7071 3268
rect 105 1649 163 1700
rect 163 1649 165 1700
rect 105 1644 165 1649
rect 900 632 952 684
rect 5800 622 5853 674
rect 7609 624 7661 677
rect 12504 621 12568 685
rect 6431 -1914 6483 -1903
rect 6431 -1948 6438 -1914
rect 6438 -1948 6472 -1914
rect 6472 -1948 6483 -1914
rect 6431 -1955 6483 -1948
rect 6431 -2110 6483 -2099
rect 6431 -2144 6438 -2110
rect 6438 -2144 6472 -2110
rect 6472 -2144 6483 -2110
rect 6431 -2151 6483 -2144
rect 6431 -2285 6483 -2274
rect 6431 -2319 6438 -2285
rect 6438 -2319 6472 -2285
rect 6472 -2319 6483 -2285
rect 6431 -2326 6483 -2319
<< metal2 >>
rect 7019 3675 7093 3679
rect 7019 3619 7028 3675
rect 7084 3619 7093 3675
rect 7019 3615 7093 3619
rect 7008 3503 7082 3507
rect 7008 3447 7017 3503
rect 7073 3447 7082 3503
rect 7008 3443 7082 3447
rect 7008 3311 7082 3315
rect 7008 3255 7017 3311
rect 7073 3255 7082 3311
rect 7008 3251 7082 3255
rect 72 1701 199 1716
rect 72 1643 102 1701
rect 169 1643 199 1701
rect 72 1625 199 1643
rect 900 687 952 2218
rect 891 684 961 687
rect 891 632 900 684
rect 952 632 961 684
rect 7609 681 7661 2222
rect 12498 685 12574 686
rect 891 624 961 632
rect 5791 674 5861 681
rect 5791 622 5800 674
rect 5853 622 5861 674
rect 7602 677 7670 681
rect 7602 624 7609 677
rect 7661 624 7670 677
rect 5791 614 5861 622
rect 12498 621 12504 685
rect 12568 621 12574 685
rect 5799 -913 5851 614
rect 12511 -900 12563 621
rect 6420 -1901 6494 -1897
rect 6420 -1957 6429 -1901
rect 6485 -1957 6494 -1901
rect 6420 -1961 6494 -1957
rect 6420 -2097 6494 -2093
rect 6420 -2153 6429 -2097
rect 6485 -2153 6494 -2097
rect 6420 -2157 6494 -2153
rect 6420 -2272 6494 -2268
rect 6420 -2328 6429 -2272
rect 6485 -2328 6494 -2272
rect 6420 -2332 6494 -2328
<< via2 >>
rect 7028 3673 7084 3675
rect 7028 3621 7030 3673
rect 7030 3621 7082 3673
rect 7082 3621 7084 3673
rect 7028 3619 7084 3621
rect 7017 3501 7073 3503
rect 7017 3449 7019 3501
rect 7019 3449 7071 3501
rect 7071 3449 7073 3501
rect 7017 3447 7073 3449
rect 7017 3309 7073 3311
rect 7017 3257 7019 3309
rect 7019 3257 7071 3309
rect 7071 3257 7073 3309
rect 7017 3255 7073 3257
rect 102 1700 169 1701
rect 102 1644 105 1700
rect 105 1644 165 1700
rect 165 1644 169 1700
rect 102 1643 169 1644
rect 6429 -1903 6485 -1901
rect 6429 -1955 6431 -1903
rect 6431 -1955 6483 -1903
rect 6483 -1955 6485 -1903
rect 6429 -1957 6485 -1955
rect 6429 -2099 6485 -2097
rect 6429 -2151 6431 -2099
rect 6431 -2151 6483 -2099
rect 6483 -2151 6485 -2099
rect 6429 -2153 6485 -2151
rect 6429 -2274 6485 -2272
rect 6429 -2326 6431 -2274
rect 6431 -2326 6483 -2274
rect 6483 -2326 6485 -2274
rect 6429 -2328 6485 -2326
<< metal3 >>
rect 6993 3679 7119 3689
rect 6993 3615 7024 3679
rect 7088 3615 7119 3679
rect 6993 3605 7119 3615
rect 6982 3507 7108 3517
rect 6982 3443 7013 3507
rect 7077 3443 7108 3507
rect 6982 3433 7108 3443
rect 6982 3315 7108 3325
rect 6982 3251 7013 3315
rect 7077 3251 7108 3315
rect 6982 3241 7108 3251
rect 49 1707 213 1734
rect 49 1701 106 1707
rect 49 1643 102 1701
rect 171 1643 213 1707
rect 49 1612 213 1643
rect 6394 -1897 6520 -1887
rect 6394 -1961 6425 -1897
rect 6489 -1961 6520 -1897
rect 6394 -1971 6520 -1961
rect 6394 -2093 6520 -2083
rect 6394 -2157 6425 -2093
rect 6489 -2157 6520 -2093
rect 6394 -2167 6520 -2157
rect 6394 -2268 6520 -2258
rect 6394 -2332 6425 -2268
rect 6489 -2332 6520 -2268
rect 6394 -2342 6520 -2332
<< via3 >>
rect 7024 3675 7088 3679
rect 7024 3619 7028 3675
rect 7028 3619 7084 3675
rect 7084 3619 7088 3675
rect 7024 3615 7088 3619
rect 7013 3503 7077 3507
rect 7013 3447 7017 3503
rect 7017 3447 7073 3503
rect 7073 3447 7077 3503
rect 7013 3443 7077 3447
rect 7013 3311 7077 3315
rect 7013 3255 7017 3311
rect 7017 3255 7073 3311
rect 7073 3255 7077 3311
rect 7013 3251 7077 3255
rect 106 1701 171 1707
rect 106 1643 169 1701
rect 169 1643 171 1701
rect 6425 -1901 6489 -1897
rect 6425 -1957 6429 -1901
rect 6429 -1957 6485 -1901
rect 6485 -1957 6489 -1901
rect 6425 -1961 6489 -1957
rect 6425 -2097 6489 -2093
rect 6425 -2153 6429 -2097
rect 6429 -2153 6485 -2097
rect 6485 -2153 6489 -2097
rect 6425 -2157 6489 -2153
rect 6425 -2272 6489 -2268
rect 6425 -2328 6429 -2272
rect 6429 -2328 6485 -2272
rect 6485 -2328 6489 -2272
rect 6425 -2332 6489 -2328
<< metal4 >>
rect 106 3854 13893 3855
rect 106 3732 13943 3854
rect 13459 3731 13943 3732
rect 6960 3679 7162 3708
rect 6960 3615 7024 3679
rect 7088 3615 7162 3679
rect 6960 3581 7162 3615
rect 6949 3507 7151 3536
rect 6949 3443 7013 3507
rect 7077 3443 7151 3507
rect 6949 3409 7151 3443
rect 6949 3315 7151 3344
rect 6949 3251 7013 3315
rect 7077 3251 7151 3315
rect 6949 3217 7151 3251
rect 3 1707 267 2547
rect 3 1643 106 1707
rect 171 1643 267 1707
rect 3 1150 267 1643
rect 13200 1150 13464 1222
rect 3 1047 13464 1150
rect 4 867 13464 1047
rect 4 483 933 867
rect 2237 483 2772 867
rect 3884 483 4284 867
rect 5779 866 13464 867
rect 5779 503 7001 866
rect 8138 503 8727 866
rect 9605 503 10116 866
rect 11111 503 11641 866
rect 12555 503 13464 866
rect 5779 483 13464 503
rect 4 256 13464 483
rect 3 217 13464 256
rect 3 120 267 217
rect 13200 -1205 13464 217
rect 6354 -1897 6573 -1868
rect 6354 -1961 6425 -1897
rect 6489 -1961 6573 -1897
rect 6354 -2002 6573 -1961
rect 6354 -2093 6573 -2064
rect 6354 -2157 6425 -2093
rect 6489 -2157 6573 -2093
rect 6354 -2198 6573 -2157
rect 6354 -2268 6573 -2239
rect 6354 -2332 6425 -2268
rect 6489 -2332 6573 -2268
rect 6354 -2373 6573 -2332
rect 13544 -2392 13943 3731
rect -2 -2536 13943 -2392
use hgu_delay_no_code  x1
timestamp 1699184232
transform 1 0 -2529 0 1 795
box 9238 267 15997 2986
use hgu_delay_no_code  x2
timestamp 1699184232
transform -1 0 22702 0 -1 526
box 9238 267 15997 2986
use hgu_delay_no_code  x3
timestamp 1699184232
transform -1 0 15993 0 -1 526
box 9238 267 15997 2986
use hgu_delay_no_code  x4
timestamp 1699184232
transform 1 0 -9238 0 1 795
box 9238 267 15997 2986
<< labels >>
flabel metal1 24 -1114 78 -1068 0 FreeSans 320 0 0 0 out
port 1 nsew
flabel metal4 106 3732 13465 3796 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel metal1 283 599 900 711 0 FreeSans 320 0 0 0 sample_delay_offset
port 4 nsew
flabel metal1 37 2391 705 2438 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel metal1 0 2774 138 2808 0 FreeSans 320 0 0 0 sample_code0[3]
port 6 nsew
flabel metal1 6709 2774 6847 2808 0 FreeSans 320 0 0 0 sample_code1[3]
port 7 nsew
flabel metal1 13326 -1487 13464 -1453 0 FreeSans 320 0 0 0 sample_code2[3]
port 8 nsew
flabel metal1 6617 -1487 6755 -1453 0 FreeSans 320 0 0 0 sample_code3[3]
port 9 nsew
flabel metal1 283 795 11682 823 0 FreeSans 320 0 0 0 sample_code1[1]
port 14 nsew
flabel metal1 283 739 12538 767 0 FreeSans 320 0 0 0 sample_code1[0]
port 15 nsew
flabel metal1 283 263 984 291 0 FreeSans 320 0 0 0 sample_code3[0]
port 16 nsew
flabel metal1 283 319 1840 347 0 FreeSans 320 0 0 0 sample_code3[1]
port 17 nsew
flabel metal1 283 375 4266 403 0 FreeSans 320 0 0 0 sample_code3[2]
port 18 nsew
flabel metal1 283 431 7693 459 0 FreeSans 320 0 0 0 sample_code2[0]
port 19 nsew
flabel metal1 283 487 8549 515 0 FreeSans 320 0 0 0 sample_code2[1]
port 20 nsew
flabel metal1 283 543 10975 571 0 FreeSans 320 0 0 0 sample_code2[2]
port 22 nsew
flabel metal1 283 851 9256 879 0 FreeSans 320 0 0 0 sample_code1[2]
port 28 nsew
flabel metal4 12555 217 13464 1150 0 FreeSans 320 0 0 0 VSS
port 30 nsew
flabel metal1 283 1019 2547 1047 0 FreeSans 320 0 0 0 sample_code0[2]
port 31 nsew
flabel metal1 283 963 4973 991 0 FreeSans 320 0 0 0 sample_code0[1]
port 32 nsew
flabel metal1 283 907 5829 935 0 FreeSans 320 0 0 0 sample_code0[0]
port 34 nsew
<< end >>
