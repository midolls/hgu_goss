* NGSPICE file created from hgu_cdac_cap_4.ext - technology: sky130A

.subckt hgu_cdac_cap_4 SUB
C0 x1[3].CTOP x1[2].CTOP 10.1f
C1 x1[3].CBOT x1[3].CTOP 10.1f
.ends

