magic
tech sky130A
magscale 1 2
timestamp 1699343576
<< nwell >>
rect -164 -122 164 262
<< pmoslvt >>
rect -35 -84 35 84
<< pdiff >>
rect -93 72 -35 84
rect -93 -72 -81 72
rect -47 -72 -35 72
rect -93 -84 -35 -72
rect 35 72 93 84
rect 35 -72 47 72
rect 81 -72 93 72
rect 35 -84 93 -72
<< pdiffc >>
rect -81 -72 -47 72
rect 47 -72 81 72
<< poly >>
rect -35 84 35 115
rect -35 -111 35 -84
<< locali >>
rect -81 72 -47 88
rect -81 -88 -47 -72
rect 47 72 81 88
rect 47 -88 81 -72
<< viali >>
rect -81 -72 -47 72
rect 47 -72 81 72
<< metal1 >>
rect -87 72 -41 84
rect -87 -72 -81 72
rect -47 -72 -41 72
rect -87 -84 -41 -72
rect 41 72 87 84
rect 41 -72 47 72
rect 81 -72 87 72
rect 41 -84 87 -72
<< properties >>
string FIXED_BBOX -178 -250 178 250
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 0.84 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
