** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic.sch
.subckt hgu_sarlogic VDD VSS COMP_RESULT READY EXT_CLK sar_clk sar_result[0] sar_result[1]
+ sar_result[2] sar_result[3] sar_result[4] sar_result[5] sar_result[6] sar_result[7] sample_clk sel_bit[0]
+ sel_bit[1] sample_delay_cap_ctrl_code[0] sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[2]
+ sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[4] sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[6]
+ sample_delay_cap_ctrl_code[7] sample_delay_cap_ctrl_code[8] sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[10]
+ sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[12] sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[14]
+ sample_delay_cap_ctrl_code[15] sample_clk_b vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6] vdd_sw[7] vdd_sw_b[1]
+ vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] vss_sw[1] vss_sw[2] vss_sw[3] vss_sw[4]
+ vss_sw[5] vss_sw[6] vss_sw[7] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4] vss_sw_b[5] vss_sw_b[6]
+ vss_sw_b[7] async_resetb_delay_cap_ctrl_code[0] async_resetb_delay_cap_ctrl_code[1]
+ async_resetb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[3] async_setb_delay_cap_ctrl_code[0]
+ async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[2] async_setb_delay_cap_ctrl_code[3] async_delay_offset
+ sample_delay_offset retimer_delay_code[0] retimer_delay_code[1] retimer_delay_code[2] retimer_delay_code[3]
+ retimer_eob_delay_offset
*.PININFO VDD:I VSS:I COMP_RESULT:I READY:I EXT_CLK:I sar_clk:O sar_result[0:7]:O sample_clk:O
*+ sel_bit[0:1]:I sample_delay_cap_ctrl_code[0:15]:I sample_clk_b:O vdd_sw[1:7]:O vdd_sw_b[1:7]:O vss_sw[1:7]:O
*+ vss_sw_b[1:7]:O async_resetb_delay_cap_ctrl_code[0:3]:I async_setb_delay_cap_ctrl_code[0:3]:I async_delay_offset:I
*+ sample_delay_offset:I retimer_delay_code[0:3]:I retimer_eob_delay_offset:I
x1 sar_clk VDD VSS sample_clk EOB READY async_delay_offset async_resetb_delay_cap_ctrl_code[0]
+ async_resetb_delay_cap_ctrl_code[1] async_resetb_delay_cap_ctrl_code[2] async_resetb_delay_cap_ctrl_code[3]
+ async_setb_delay_cap_ctrl_code[0] async_setb_delay_cap_ctrl_code[1] async_setb_delay_cap_ctrl_code[2]
+ async_setb_delay_cap_ctrl_code[3] hgu_clk_async
x2 sample_clk_b VDD VSS EXT_CLK VSS VSS sample_clk sample_delay_cap_ctrl_code[0]
+ sample_delay_cap_ctrl_code[1] sample_delay_cap_ctrl_code[2] sample_delay_cap_ctrl_code[3] sample_delay_cap_ctrl_code[4]
+ sample_delay_cap_ctrl_code[5] sample_delay_cap_ctrl_code[6] sample_delay_cap_ctrl_code[7] sample_delay_cap_ctrl_code[8]
+ sample_delay_cap_ctrl_code[9] sample_delay_cap_ctrl_code[10] sample_delay_cap_ctrl_code[11] sample_delay_cap_ctrl_code[12]
+ sample_delay_cap_ctrl_code[13] sample_delay_cap_ctrl_code[14] sample_delay_cap_ctrl_code[15] sample_delay_offset hgu_clk_sample
x3 sel_bit[0] sel_bit[1] EOB sar_clk sar_result_temp[0] sar_result_temp[1] sar_result_temp[2]
+ sar_result_temp[3] sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] COMP_RESULT check[0]
+ check[1] check[2] check[3] check[4] check[5] check[6] sample_clk_b VDD VSS hgu_sarlogic_8bit_logic
x4 VDD VSS vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6] vdd_sw[7] vdd_sw_b[1]
+ vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] sar_result_temp[1] sar_result_temp[2]
+ sar_result_temp[3] sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] vss_sw[1] vss_sw[2]
+ vss_sw[3] vss_sw[4] vss_sw[5] vss_sw[6] vss_sw[7] check[0] check[1] check[2] check[3] check[4] check[5]
+ check[6] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4] vss_sw_b[5] vss_sw_b[6] vss_sw_b[7] sar_clk
+ sample_clk_b hgu_sarlogic_sw_ctrl
x5 VDD VSS sar_result_temp[0] sar_result_temp[1] sar_result_temp[2] sar_result_temp[3]
+ sar_result_temp[4] sar_result_temp[5] sar_result_temp[6] sar_result_temp[7] EOB retimer_delay_code[0]
+ retimer_delay_code[1] retimer_delay_code[2] retimer_delay_code[3] retimer_eob_delay_offset sar_result[0] sar_result[1]
+ sar_result[2] sar_result[3] sar_result[4] sar_result[5] sar_result[6] sar_result[7] hgu_sarlogic_retimer
**** begin user architecture code


.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include /foss/designs/hgu_goss/hgu/mag/hgu_cdac_unit.spice



**** end user architecture code
.ends

* expanding   symbol:  ../xschem/hgu_clk_async.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_async.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_async.sch
.subckt hgu_clk_async ASYNC_CLK_SAR VDD VSS sample_clk EOB READY delay_offset
+ async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1] async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[3]
+ async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[1] async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[3]
*.PININFO VDD:I ASYNC_CLK_SAR:O VSS:I sample_clk:I EOB:I READY:I async_resetb_delay_ctrl_code[0:3]:I
*+ async_setb_delay_ctrl_code[0:3]:I delay_offset:I
x3 net1 VSS sample_clk VSS VSS vDD VDD net4 sky130_fd_sc_hd__mux2_1
x8 net4 VSS EOB VSS VSS vDD VDD ASYNC_CLK_SAR sky130_fd_sc_hd__mux2_1
x27 sample_clk VDD net5 net6 VSS VSS vDD VDD net1 net7 sky130_fd_sc_hd__dfbbp_1
x9 net2 VSS VSS vDD VDD net6 sky130_fd_sc_hd__inv_1
x10 net3 VSS VSS vDD VDD net5 sky130_fd_sc_hd__inv_1
x2 VDD READY net2 VSS async_setb_delay_ctrl_code[0] async_setb_delay_ctrl_code[1]
+ async_setb_delay_ctrl_code[2] async_setb_delay_ctrl_code[3] delay_offset hgu_delay_no_code
x4 VDD ASYNC_CLK_SAR net3 VSS async_resetb_delay_ctrl_code[0] async_resetb_delay_ctrl_code[1]
+ async_resetb_delay_ctrl_code[2] async_resetb_delay_ctrl_code[3] delay_offset hgu_delay_no_code

.ends


* expanding   symbol:  ../xschem/hgu_clk_sample.sym # of pins=12
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_sample.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_sample.sch
.subckt hgu_clk_sample SAMPLE_CLK_b VDD VSS CLK RESET SET SAMPLE_CLK CAP_CTRL_CODE0[0]
+ CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[3] CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[2]
+ CAP_CTRL_CODE1[3] CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[1] CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[3] CAP_CTRL_CODE3[0]
+ CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[3] sample_delay_offset
*.PININFO VDD:I VSS:I SET:I RESET:I CLK:I SAMPLE_CLK:O SAMPLE_CLK_b:O CAP_CTRL_CODE1[0:3]:I
*+ CAP_CTRL_CODE2[0:3]:I CAP_CTRL_CODE3[0:3]:I CAP_CTRL_CODE0[0:3]:I sample_delay_offset:I
x1 VDD VSS CLK net2 RESET SET hgu_clk_div
x2 net8 net2 VDD VSS CAP_CTRL_CODE0[0] CAP_CTRL_CODE0[1] CAP_CTRL_CODE0[2] CAP_CTRL_CODE0[3]
+ CAP_CTRL_CODE1[0] CAP_CTRL_CODE1[1] CAP_CTRL_CODE1[2] CAP_CTRL_CODE1[3] CAP_CTRL_CODE2[0] CAP_CTRL_CODE2[1]
+ CAP_CTRL_CODE2[2] CAP_CTRL_CODE2[3] CAP_CTRL_CODE3[0] CAP_CTRL_CODE3[1] CAP_CTRL_CODE3[2] CAP_CTRL_CODE3[3]
+ sample_delay_offset hgu_delay
x7 net8 VSS VSS vDD VDD net1 sky130_fd_sc_hd__inv_1

x3 net2 net1 VSS VSS vDD VDD net4 sky130_fd_sc_hd__nand2_1
XM7 net7 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 net7 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.26 nf=1 m=1
XM9 net5 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net5 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=1 m=1
XM11 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 net6 net5 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.26 nf=1 m=1
XM13 net4 VSS net3 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.9 nf=1 m=1
XM14 net4 VDD net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM18 SAMPLE_CLK_b net7 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=3 m=1
XM17 SAMPLE_CLK_b net7 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.78 nf=3 m=1
XM15 SAMPLE_CLK net6 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=3 m=1
XM16 SAMPLE_CLK net6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.78 nf=3 m=1
.ends


* expanding   symbol:  ../xschem/hgu_sarlogic_8bit_logic.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_8bit_logic.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_8bit_logic.sch
.subckt hgu_sarlogic_8bit_logic sel_bit[0] sel_bit[1] EOB clk_sar D[0] D[1] D[2] D[3] D[4] D[5] D[6]
+ D[7] comparator_out check[0] check[1] check[2] check[3] check[4] check[5] check[6] reset VDD VSS
*.PININFO clk_sar:I VDD:I VSS:I comparator_out:I reset:I EOB:O D[0:7]:O check[0:6]:O sel_bit[0:1]:I
x20 clk_sar_buff EOB VDD resetb VSS VSS VDD VDD net1 net4 sky130_fd_sc_hd__dfbbp_1
x27 clk_sar_buff net1 resetb VDD VSS VSS VDD VDD check[6] net5 sky130_fd_sc_hd__dfbbp_1
x30 clk_sar_buff check[6] resetb VDD VSS VSS VDD VDD check[5] net6 sky130_fd_sc_hd__dfbbp_1
x33 clk_sar_buff check[5] resetb VDD VSS VSS VDD VDD check[4] net7 sky130_fd_sc_hd__dfbbp_1
x36 clk_sar_buff check[4] resetb VDD VSS VSS VDD VDD check[3] net8 sky130_fd_sc_hd__dfbbp_1
x39 clk_sar_buff check[3] resetb VDD VSS VSS VDD VDD check[2] net9 sky130_fd_sc_hd__dfbbp_1
x42 clk_sar_buff check[2] resetb VDD VSS VSS VDD VDD check[1] net10 sky130_fd_sc_hd__dfbbp_1
x45 clk_sar_buff check[1] resetb VDD VSS VSS VDD VDD check[0] net11 sky130_fd_sc_hd__dfbbp_1
x48 clk_sar_buff check[0] resetb VDD VSS VSS VDD VDD net3 net12 sky130_fd_sc_hd__dfbbp_1
x51 D[6] comparator_out_buff resetb net4 VSS VSS VDD VDD D[7] net13 sky130_fd_sc_hd__dfbbp_1
x54 D[5] comparator_out_buff resetb net5 VSS VSS VDD VDD D[6] net14 sky130_fd_sc_hd__dfbbp_1
x57 D[4] comparator_out_buff resetb net6 VSS VSS VDD VDD D[5] net15 sky130_fd_sc_hd__dfbbp_1
x60 D[3] comparator_out_buff resetb net7 VSS VSS VDD VDD D[4] net16 sky130_fd_sc_hd__dfbbp_1
x63 D[2] comparator_out_buff resetb net8 VSS VSS VDD VDD D[3] net17 sky130_fd_sc_hd__dfbbp_1
x66 D[1] comparator_out_buff resetb net9 VSS VSS VDD VDD D[2] net18 sky130_fd_sc_hd__dfbbp_1
x69 D[0] comparator_out_buff resetb net10 VSS VSS VDD VDD D[1] net19 sky130_fd_sc_hd__dfbbp_1
x72 net2 comparator_out_buff resetb net11 VSS VSS VDD VDD D[0] net20 sky130_fd_sc_hd__dfbbp_1
x75 VSS VSS resetb net21 VSS VSS VDD VDD net2 net22 sky130_fd_sc_hd__dfbbp_1
x77 EOB VSS VSS VDD VDD net21 sky130_fd_sc_hd__inv_1
x78 check[2] check[1] check[0] net3 sel_bit[0] sel_bit[1] VSS VSS VDD VDD EOB
+ sky130_fd_sc_hd__mux4_4

x1 reset VSS VSS VDD VDD net23 sky130_fd_sc_hd__buf_1
x2 clk_sar VSS VSS VDD VDD net24 sky130_fd_sc_hd__buf_1
x3 net23 VSS VSS VDD VDD net25 sky130_fd_sc_hd__buf_4
x4 net25 VSS VSS VDD VDD resetb sky130_fd_sc_hd__buf_16
x5 net24 VSS VSS VDD VDD clk_sar_buff sky130_fd_sc_hd__buf_4
x6 comparator_out VSS VSS VDD VDD net26 sky130_fd_sc_hd__buf_1
x7 net26 VSS VSS VDD VDD comparator_out_buff sky130_fd_sc_hd__buf_4
.ends


* expanding   symbol:  ../xschem/hgu_sarlogic_sw_ctrl.sym # of pins=10
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_sw_ctrl.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_sw_ctrl.sch
.subckt hgu_sarlogic_sw_ctrl VDD VSS vdd_sw[1] vdd_sw[2] vdd_sw[3] vdd_sw[4] vdd_sw[5] vdd_sw[6]
+ vdd_sw[7] vdd_sw_b[1] vdd_sw_b[2] vdd_sw_b[3] vdd_sw_b[4] vdd_sw_b[5] vdd_sw_b[6] vdd_sw_b[7] D[1] D[2] D[3]
+ D[4] D[5] D[6] D[7] vss_sw[1] vss_sw[2] vss_sw[3] vss_sw[4] vss_sw[5] vss_sw[6] vss_sw[7] check[0]
+ check[1] check[2] check[3] check[4] check[5] check[6] vss_sw_b[1] vss_sw_b[2] vss_sw_b[3] vss_sw_b[4]
+ vss_sw_b[5] vss_sw_b[6] vss_sw_b[7] READY reset
*.PININFO vdd_sw[1:7]:O vdd_sw_b[1:7]:O vss_sw[1:7]:O vss_sw_b[1:7]:O VDD:I VSS:I READY:I D[1:7]:I
*+ check[0:6]:I reset:I
x4 net1 D[7] VDD resetb VSS VSS VDD VDD vdd_sw[7] vdd_sw_b[7] sky130_fd_sc_hd__dfbbn_1
x5 net2 D[7] resetb VDD VSS VSS VDD VDD vss_sw[7] vss_sw_b[7] sky130_fd_sc_hd__dfbbn_1
x19 net3 D[6] VDD resetb VSS VSS VDD VDD vdd_sw[6] vdd_sw_b[6] sky130_fd_sc_hd__dfbbn_1
x21 net4 D[6] resetb VDD VSS VSS VDD VDD vss_sw[6] vss_sw_b[6] sky130_fd_sc_hd__dfbbn_1
x23 net5 D[5] VDD resetb VSS VSS VDD VDD vdd_sw[5] vdd_sw_b[5] sky130_fd_sc_hd__dfbbn_1
x24 net6 D[5] resetb VDD VSS VSS VDD VDD vss_sw[5] vss_sw_b[5] sky130_fd_sc_hd__dfbbn_1
x25 net7 D[4] VDD resetb VSS VSS VDD VDD vdd_sw[4] vdd_sw_b[4] sky130_fd_sc_hd__dfbbn_1
x26 net8 D[4] resetb VDD VSS VSS VDD VDD vss_sw[4] vss_sw_b[4] sky130_fd_sc_hd__dfbbn_1
x28 net9 D[3] VDD resetb VSS VSS VDD VDD vdd_sw[3] vdd_sw_b[3] sky130_fd_sc_hd__dfbbn_1
x29 net10 D[3] resetb VDD VSS VSS VDD VDD vss_sw[3] vss_sw_b[3] sky130_fd_sc_hd__dfbbn_1
x31 net11 D[2] VDD resetb VSS VSS VDD VDD vdd_sw[2] vdd_sw_b[2] sky130_fd_sc_hd__dfbbn_1
x32 net12 D[2] resetb VDD VSS VSS VDD VDD vss_sw[2] vss_sw_b[2] sky130_fd_sc_hd__dfbbn_1
x34 net13 D[1] VDD resetb VSS VSS VDD VDD vdd_sw[1] vdd_sw_b[1] sky130_fd_sc_hd__dfbbn_1
x35 net14 D[1] resetb VDD VSS VSS VDD VDD vss_sw[1] vss_sw_b[1] sky130_fd_sc_hd__dfbbn_1
x6 VSS READY_buff check[6] VSS VSS VDD VDD net1 sky130_fd_sc_hd__mux2_1
x7 VSS READY_buff check[6] VSS VSS VDD VDD net2 sky130_fd_sc_hd__mux2_1
x8 VSS READY_buff check[5] VSS VSS VDD VDD net3 sky130_fd_sc_hd__mux2_1
x9 VSS READY_buff check[5] VSS VSS VDD VDD net4 sky130_fd_sc_hd__mux2_1
x10 VSS READY_buff check[4] VSS VSS VDD VDD net5 sky130_fd_sc_hd__mux2_1
x11 VSS READY_buff check[4] VSS VSS VDD VDD net6 sky130_fd_sc_hd__mux2_1
x12 VSS READY_buff check[3] VSS VSS VDD VDD net7 sky130_fd_sc_hd__mux2_1
x13 VSS READY_buff check[3] VSS VSS VDD VDD net8 sky130_fd_sc_hd__mux2_1
x14 VSS READY_buff check[2] VSS VSS VDD VDD net9 sky130_fd_sc_hd__mux2_1
x15 VSS READY_buff check[2] VSS VSS VDD VDD net10 sky130_fd_sc_hd__mux2_1
x16 VSS READY_buff check[1] VSS VSS VDD VDD net11 sky130_fd_sc_hd__mux2_1
x17 VSS READY_buff check[1] VSS VSS VDD VDD net12 sky130_fd_sc_hd__mux2_1
x18 VSS READY_buff check[0] VSS VSS VDD VDD net13 sky130_fd_sc_hd__mux2_1
x20 VSS READY_buff check[0] VSS VSS VDD VDD net14 sky130_fd_sc_hd__mux2_1
x1 reset VSS VSS VDD VDD net15 sky130_fd_sc_hd__buf_1
x3 net15 VSS VSS VDD VDD net16 sky130_fd_sc_hd__buf_4
x2 net16 VSS VSS VDD VDD resetb sky130_fd_sc_hd__buf_16
x22 READY VSS VSS VDD VDD net17 sky130_fd_sc_hd__buf_1
x27 net17 VSS VSS VDD VDD net18 sky130_fd_sc_hd__buf_4
x30 net18 VSS VSS VDD VDD READY_buff sky130_fd_sc_hd__buf_16
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sym # of pins=7
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sarlogic_retimer.sch
.subckt hgu_sarlogic_retimer VDD VSS sar_logic[0] sar_logic[1] sar_logic[2] sar_logic[3]
+ sar_logic[4] sar_logic[5] sar_logic[6] sar_logic[7] eob delay_code[0] delay_code[1] delay_code[2] delay_code[3]
+ delay_offset sar_retimer[0] sar_retimer[1] sar_retimer[2] sar_retimer[3] sar_retimer[4] sar_retimer[5]
+ sar_retimer[6] sar_retimer[7]
*.PININFO sar_logic[0:7]:I sar_retimer[0:7]:O eob:I VDD:I VSS:I delay_code[0:3]:I delay_offset:I
x1[0] eob_delay sar_logic[0] VDD VDD VSS VSS VDD VDD sar_retimer[0] net2[7] sky130_fd_sc_hd__dfbbp_1
x1[1] eob_delay sar_logic[1] VDD VDD VSS VSS VDD VDD sar_retimer[1] net2[6] sky130_fd_sc_hd__dfbbp_1
x1[2] eob_delay sar_logic[2] VDD VDD VSS VSS VDD VDD sar_retimer[2] net2[5] sky130_fd_sc_hd__dfbbp_1
x1[3] eob_delay sar_logic[3] VDD VDD VSS VSS VDD VDD sar_retimer[3] net2[4] sky130_fd_sc_hd__dfbbp_1
x1[4] eob_delay sar_logic[4] VDD VDD VSS VSS VDD VDD sar_retimer[4] net2[3] sky130_fd_sc_hd__dfbbp_1
x1[5] eob_delay sar_logic[5] VDD VDD VSS VSS VDD VDD sar_retimer[5] net2[2] sky130_fd_sc_hd__dfbbp_1
x1[6] eob_delay sar_logic[6] VDD VDD VSS VSS VDD VDD sar_retimer[6] net2[1] sky130_fd_sc_hd__dfbbp_1
x1[7] eob_delay sar_logic[7] VDD VDD VSS VSS VDD VDD sar_retimer[7] net2[0] sky130_fd_sc_hd__dfbbp_1
x2 VDD eob net1 VSS delay_code[0] delay_code[1] delay_code[2] delay_code[3] delay_offset
+ hgu_delay_no_code
x3 net1 VSS VSS VDD VDD eob_delay sky130_fd_sc_hd__buf_2
.ends


* expanding   symbol:  ../xschem/hgu_delay_no_code.sym # of pins=6
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sch
.subckt hgu_delay_no_code VDD IN OUT VSS code[0] code[1] code[2] code[3] code_offset
*.PININFO IN:I VDD:I VSS:I OUT:O code[0:3]:I code_offset:I
XM13 OUT net1 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM15 net3 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM46 OUT net1 net2 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM47 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
x2 code[0] VSS net1 net6 hgu_sw_cap
x3[1] code[1] VSS net1 net7 hgu_sw_cap
x3[0] code[1] VSS net1 net7 hgu_sw_cap
x4[3] code[2] VSS net1 net8 hgu_sw_cap
x4[2] code[2] VSS net1 net8 hgu_sw_cap
x4[1] code[2] VSS net1 net8 hgu_sw_cap
x4[0] code[2] VSS net1 net8 hgu_sw_cap
x5[7] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[6] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[5] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[4] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[3] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[2] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[1] net4 net1 VDD net9 hgu_sw_cap_pmos
x5[0] net4 net1 VDD net9 hgu_sw_cap_pmos
x10 code[3] VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x7 code_offset VSS net1 net10 hgu_sw_cap
x6 net5 net1 VDD net11 hgu_sw_cap_pmos
x11 code_offset VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x8 VDD IN net1 hgu_pfet_hvt_stack_in_delay
x9 IN net1 VSS hgu_nfet_hvt_stack_in_delay
XM48 VSS OUT net2 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.84 nf=2 m=1
XM1 VDD OUT net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 m=1
.ends


* expanding   symbol:  ../xschem/hgu_clk_div.sym # of pins=6
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_div.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_div.sch
.subckt hgu_clk_div VDD VSS CLK DIV_CLK RESET SET
*.PININFO DIV_CLK:O SET:I RESET:I CLK:I VDD:I VSS:I
x2 CLK D_loop net1 net2 VSS VSS vDD VDD DIV_CLK D_loop sky130_fd_sc_hd__dfbbp_1
x3 SET VSS VSS vDD VDD net2 sky130_fd_sc_hd__inv_1
x4 RESET VSS VSS vDD VDD net1 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  ../xschem/hgu_delay.sym # of pins=9
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay.sch
.subckt hgu_delay OUT IN VDD VSS SAMPLE_CODE0[0] SAMPLE_CODE0[1] SAMPLE_CODE0[2] SAMPLE_CODE0[3]
+ SAMPLE_CODE1[0] SAMPLE_CODE1[1] SAMPLE_CODE1[2] SAMPLE_CODE1[3] SAMPLE_CODE2[0] SAMPLE_CODE2[1] SAMPLE_CODE2[2]
+ SAMPLE_CODE2[3] SAMPLE_CODE3[0] SAMPLE_CODE3[1] SAMPLE_CODE3[2] SAMPLE_CODE3[3] sample_delay_offset
*.PININFO IN:I VDD:I VSS:I OUT:O SAMPLE_CODE1[0:3]:I SAMPLE_CODE2[0:3]:I SAMPLE_CODE3[0:3]:I
*+ SAMPLE_CODE0[0:3]:I sample_delay_offset:I
x4 VDD IN net1 VSS SAMPLE_CODE0[0] SAMPLE_CODE0[1] SAMPLE_CODE0[2] SAMPLE_CODE0[3]
+ sample_delay_offset hgu_delay_no_code
x1 VDD net1 net2 VSS SAMPLE_CODE1[0] SAMPLE_CODE1[1] SAMPLE_CODE1[2] SAMPLE_CODE1[3]
+ sample_delay_offset hgu_delay_no_code
x2 VDD net2 net3 VSS SAMPLE_CODE2[0] SAMPLE_CODE2[1] SAMPLE_CODE2[2] SAMPLE_CODE2[3]
+ sample_delay_offset hgu_delay_no_code
x3 VDD net3 OUT VSS SAMPLE_CODE3[0] SAMPLE_CODE3[1] SAMPLE_CODE3[2] SAMPLE_CODE3[3]
+ sample_delay_offset hgu_delay_no_code
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sym # of pins=4
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap.sch
.subckt hgu_sw_cap SW VSS DELAY_SIGNAL floating
*.PININFO SW:I VSS:I DELAY_SIGNAL:B floating:B
XM14 DELAY_SIGNAL SW floating VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
*x2 floating VSS VSS hgu_cdac_unit
.ends


* expanding   symbol:  /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sym # of pins=4
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_sw_cap_pmos.sch
.subckt hgu_sw_cap_pmos SW DELAY_SIGNAL VDD floating
*.PININFO SW:I VDD:I DELAY_SIGNAL:B floating:B
XM16 floating SW DELAY_SIGNAL VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
*x1 VDD floating VDD hgu_cdac_unit
.ends


* expanding   symbol:
*+  /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sym # of pins=3
** sym_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sym
** sch_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_pfet_hvt_stack_in_delay.sch
.subckt hgu_pfet_hvt_stack_in_delay VDD input_stack output_stack
*.PININFO VDD:I input_stack:I output_stack:B
XM1 output_stack input_stack net1 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM2 net1 input_stack net2 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM3 net2 input_stack net3 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM4 net3 input_stack net4 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM5 net4 input_stack net5 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
XM6 net5 input_stack VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.42 nf=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sym # of pins=3
** sym_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sym
** sch_path:
*+ /foss/designs/hgu_goss/hgu/xschem/../../../hgu_goss/hgu/xschem/hgu_nfet_hvt_stack_in_delay.sch
.subckt hgu_nfet_hvt_stack_in_delay input_stack output_stack VSS
*.PININFO VSS:I input_stack:I output_stack:B
XM1 output_stack input_stack net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 net1 input_stack net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM3 net2 input_stack net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net3 input_stack net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 net4 input_stack net5 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 net5 input_stack net6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM7 net6 input_stack net7 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 net7 input_stack net8 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM9 net8 input_stack net9 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net9 input_stack net10 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 net10 input_stack net11 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 net11 input_stack net12 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM13 net12 input_stack net13 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM14 net13 input_stack net14 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM15 net14 input_stack net15 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM16 net15 input_stack VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends

.end
