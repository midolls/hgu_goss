* NGSPICE file created from hgu_sarlogic_8bit_logic_flat.ext - technology: sky130A

.subckt hgu_sarlogic_8bit_logic_flat sel_bit[0] sel_bit[1] reset eob comparator_out
+ D[7] D[6] check[6] D[5] check[0] check[5] check[1] check[4] check[2] check[3] D[2]
+ D[3] D[1] D[4] D[0] clk_sar VSS VDD
X0 VDD.t61 a_10680_2340# D[3].t1 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1 VDD.t86 a_8289_4086# check[1].t1 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 VDD.t549 D[0].t2 a_8236_3239# VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3 VDD.t418 a_2389_5648# eob.t4 VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X4 a_12030_3213# a_11856_3239# a_12146_3239# VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X5 VDD.t198 a_1338_5674# x5.X.t3 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_4971_4801# VDD.t743 VSS.t174 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 a_2147_5083# a_1682_4775# VDD.t395 VDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X8 a_1822_4801# x4.X.t32 VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X9 a_11330_2340# a_11628_2640# a_11564_2732# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X10 VSS.t252 a_12030_3213# a_12737_3239# VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_4213_3239# a_4367_3213# a_4073_3213# VSS.t601 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X12 a_8591_4801# check[5].t2 VSS.t423 VSS.t422 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X13 a_9710_4296# a_9238_4086# a_9954_4478# VDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X14 VSS.t593 x30.Q_N a_7185_2366# VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X15 VDD.t543 a_11250_4775# a_11160_5167# VDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X16 VSS.t413 a_5992_4086# x45.Q_N VSS.t412 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_3599_2340# a_3912_2366# a_4018_2366# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X18 x72.Q_N a_7246_3213# VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X19 VSS.t360 x27.Q_N a_4018_2366# VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X20 a_4854_3213# x77.Y VDD.t670 VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 a_7072_3239# a_5844_3239# a_6930_3521# VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X22 a_9442_4086# a_8697_4112# a_9578_4112# VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X23 VSS.t268 x4.X.t33 a_9151_3213# VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X24 VDD.t132 a_7246_3213# a_7158_3605# VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X25 VDD.t39 a_5897_4086# check[0].t0 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X26 a_11089_4112# x4.X.t34 VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X27 a_4793_2366# a_4925_2550# a_4657_2340# VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 VDD.t10 x75.Q a_5844_3239# VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_6978_4801# a_6466_4775# VSS.t302 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X30 a_4388_2732# a_3599_2340# VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X31 a_2788_5674# check[2].t2 VSS.t577 VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.107 ps=1 w=0.42 l=0.15
X32 a_10794_3239# a_10628_3239# VDD.t255 VDD.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 VSS.t673 D[0].t3 a_8236_3239# VSS.t672 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X34 VDD.t112 x4.X.t35 a_4368_4775# VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X35 a_9465_4801# a_8403_4801# a_9370_4801# VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X36 VSS.t356 a_1511_4112# x4.X.t31 VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_12048_4394# a_11089_4112# VDD.t280 VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X38 a_9101_3521# a_8683_3605# a_8857_3213# VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X39 a_7247_4775# VDD.t187 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X40 VDD.t682 a_6846_4086# a_6845_4386# VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X41 VSS.t116 x20.Q_N a_1626_2366# VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X42 D[2].t1 a_12737_3239# VSS.t603 VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X43 a_11250_4775# a_11076_5167# a_11390_4801# VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X44 a_4680_3239# a_3452_3239# a_4538_3521# VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X45 a_2479_2648# a_1520_2366# VDD.t488 VDD.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X46 VDD.t48 a_4854_3213# a_4766_3605# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X47 a_11184_4801# a_10795_4801# a_11076_5167# VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X48 a_2784_5996# check[2].t3 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.154 ps=1.34 w=0.64 l=0.15
X49 a_4593_4112# a_4453_4386# a_4155_4086# VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X50 a_1996_2732# a_1207_2340# VDD.t591 VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X51 a_7181_3239# a_5844_3239# a_7072_3239# VSS.t574 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X52 a_6198_3239# x7.X VSS.t619 VSS.t618 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X53 x4.X.t15 a_1511_4112# VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X54 a_2265_2340# a_1520_2366# a_2401_2366# VSS.t461 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X55 a_12031_4775# a_11857_4801# a_12147_4801# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X56 VSS.t12 x75.Q a_5844_3239# VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 VDD.t186 VDD.t184 a_1976_4775# VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X58 VSS.t651 a_7050_4086# a_6985_4112# VSS.t650 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X59 a_1762_2340# a_2060_2640# a_1996_2732# VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X60 VDD.t539 check[1].t2 a_2969_6040# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.138 ps=1.16 w=0.64 l=0.15
X61 a_2883_5674# a_2853_5648# a_2788_5674# VSS.t645 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.066 ps=0.745 w=0.36 l=0.15
X62 a_7562_4478# a_7050_4086# VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X63 a_10775_2340# a_11088_2366# a_11194_2366# VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X64 a_6504_2648# a_6304_2366# VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X65 a_4214_4801# a_4368_4775# a_4074_4775# VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X66 VSS.t683 x36.Q_N a_11194_2366# VSS.t682 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X67 a_10794_3239# a_10628_3239# VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 a_1511_4112# x4.A VSS.t540 VSS.t539 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X69 a_4855_4775# VDD.t181 VDD.t183 VDD.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X70 a_7073_4801# a_5845_4801# a_6931_5083# VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X71 VDD.t67 a_4454_4086# a_4453_4386# VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X72 VDD.t320 a_7247_4775# a_7159_5167# VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X73 x4.A a_897_4112# VDD.t603 VDD.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 VDD.t196 a_1338_5674# x5.X.t2 VDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X75 x30.Q_N a_7247_4775# VSS.t293 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X76 x4.X.t14 a_1511_4112# VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 a_12345_2732# a_11833_2340# VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X78 VSS.t407 check[0].t2 a_5372_4112# VSS.t406 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X79 a_8803_4112# a_8939_4086# a_8384_4086# VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X80 VSS.t118 x4.X.t36 a_9152_4775# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X81 a_3806_3239# VSS.t544 VSS.t546 VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X82 VDD.t108 x20.Q_N a_1207_2340# VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X83 VSS.t230 check[1].t3 a_2993_5674# VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0786 ps=0.805 w=0.42 l=0.15
X84 VSS.t172 VDD.t744 a_8803_4112# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X85 VSS.t443 a_10776_4086# x39.Q_N VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X86 a_6291_3605# a_5844_3239# a_6198_3239# VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X87 x75.Q_N a_4854_3213# VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X88 VSS.t415 x5.X.t8 a_8237_4801# VSS.t414 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X89 VSS.t473 a_6465_3213# a_6399_3239# VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X90 a_1822_4801# a_1976_4775# a_1682_4775# VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X91 VDD.t496 a_10775_2340# x63.Q_N VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X92 a_9102_5083# a_8684_5167# a_8858_4775# VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X93 a_11856_3239# a_10628_3239# a_11714_3521# VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X94 a_4681_4801# a_3453_4801# a_4539_5083# VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X95 VDD.t104 a_4855_4775# a_4767_5167# VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X96 a_9953_2366# a_9441_2340# VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X97 check[3].t1 a_12738_4801# VSS.t437 VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X98 a_11769_4112# a_11629_4386# a_11331_4086# VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X99 a_1112_2340# a_1207_2340# VSS.t556 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X100 x7.X a_929_3238# VSS.t663 VSS.t662 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X101 a_2579_4801# x4.X.t37 VSS.t435 VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X102 a_4155_4086# a_4453_4386# a_4389_4478# VDD.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X103 a_7480_3521# a_7072_3239# a_7246_3213# VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X104 VSS.t170 VDD.t745 a_9578_4112# VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X105 a_5992_4086# a_6305_4112# a_6411_4112# VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X106 VDD.t658 x7.X a_12547_2366# VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X107 a_6199_4801# check[6].t2 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X108 a_7182_4801# a_5845_4801# a_7073_4801# VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X109 VSS.t168 VDD.t746 a_6411_4112# VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X110 VDD.t456 x4.X.t38 a_6759_3213# VDD.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X111 x33.Q_N a_9639_4775# VSS.t311 VSS.t310 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X112 VSS.t358 x27.Q_N a_4793_2366# VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X113 a_3899_3605# a_3452_3239# a_3806_3239# VSS.t378 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X114 VSS.t417 x5.X.t9 a_5845_4801# VSS.t416 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X115 D[1].t0 a_10345_3239# VDD.t665 VDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X116 a_6710_5083# a_6292_5167# a_6466_4775# VDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X117 a_11195_4112# a_11331_4086# a_10776_4086# VSS.t240 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X118 a_6375_3605# a_5844_3239# a_6291_3605# VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 a_2969_6040# a_2853_5648# a_2883_5674# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.0567 ps=0.69 w=0.42 l=0.15
X120 a_8288_2340# a_8383_2340# VDD.t730 VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X121 a_10795_4801# a_10629_4801# VSS.t266 VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X122 a_7050_4086# a_6305_4112# a_7186_4112# VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X123 a_11965_3239# a_10628_3239# a_11856_3239# VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X124 a_12102_4296# a_11629_4386# a_12346_4112# VSS.t475 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X125 VSS.t209 a_2463_4775# a_3170_4801# VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X126 a_11970_4112# a_12102_4296# a_11834_4086# VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X127 VDD.t126 a_3505_4086# x48.Q VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X128 a_8590_3239# x7.X VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X129 VDD.t579 VSS.t692 a_3452_3239# VDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X130 x4.X.t13 a_1511_4112# VDD.t379 VDD.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X131 a_4113_4394# a_3913_4112# VDD.t240 VDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X132 VSS.t364 a_11834_4086# a_11769_4112# VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X133 a_3807_4801# x27.D VSS.t579 VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X134 a_4790_4801# a_3453_4801# a_4681_4801# VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X135 VSS.t114 x20.Q_N a_2401_2366# VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X136 VDD.t716 a_929_3238# x7.X VDD.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X137 a_1511_4112# x4.A VSS.t538 VSS.t537 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X138 a_11564_2366# a_10775_2340# VSS.t469 VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X139 a_7763_2366# a_6844_2640# a_7317_2550# VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 a_11714_3521# a_11249_3213# VDD.t344 VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X141 a_11857_4801# a_10629_4801# a_11715_5083# VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X142 x4.A a_897_4112# VDD.t601 VDD.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X143 a_6292_5167# a_5845_4801# a_6199_4801# VSS.t686 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X144 VDD.t589 a_1207_2340# x51.Q_N VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X145 a_3983_3605# a_3452_3239# a_3899_3605# VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 a_2389_5648# a_3258_5648# a_2883_5674# VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X147 a_5896_2340# a_5991_2340# VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X148 VSS.t300 a_6466_4775# a_6400_4801# VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X149 a_4658_4086# a_3913_4112# a_4794_4112# VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X150 VDD.t228 a_2463_4775# a_3170_4801# VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X151 a_7481_5083# a_7073_4801# a_7247_4775# VDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X152 a_9237_2340# D[3].t2 VDD.t214 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X153 VDD.t236 reset.t0 a_621_4112# VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X154 a_9173_4112# a_8384_4086# VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X155 VDD.t654 x7.X a_2979_2366# VDD.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X156 VDD.t474 a_11833_2340# a_11766_2732# VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X157 VSS.t543 VSS.t541 a_3452_3239# VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X158 VDD.t276 a_9442_4086# a_9375_4478# VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X159 VDD.t630 x30.Q_N a_7049_2340# VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X160 a_4317_3521# a_3899_3605# a_4073_3213# VDD.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X161 a_6376_5167# a_5845_4801# a_6292_5167# VDD.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X162 a_3900_5167# a_3453_4801# a_3807_4801# VSS.t277 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X163 VSS.t679 a_8383_2340# x60.Q_N VSS.t678 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X164 a_11249_3213# x39.Q_N VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X165 x7.X a_929_3238# VSS.t661 VSS.t660 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X166 a_1227_4801# a_1061_4801# VSS.t482 VSS.t481 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 a_4074_4775# VDD.t178 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X168 a_8997_3239# x42.Q_N VSS.t490 VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X169 a_8591_4801# check[5].t3 VDD.t674 VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X170 a_11289_4394# a_11089_4112# VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X171 a_1511_4112# x4.A VDD.t577 VDD.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X172 x4.X.t30 a_1511_4112# VSS.t354 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X173 x75.Q a_5561_3239# VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X174 a_11966_4801# a_10629_4801# a_11857_4801# VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X175 a_9376_2366# a_9236_2640# a_8938_2340# VSS.t304 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X176 eob.t5 a_2389_5648# VSS.t395 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X177 a_6781_4112# a_5992_4086# VSS.t411 VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X178 x77.Y eob.t8 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X179 x5.X.t7 a_1338_5674# VSS.t183 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 a_9237_2340# D[3].t3 VSS.t195 VSS.t194 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X181 a_11715_5083# a_11250_4775# VDD.t541 VDD.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X182 x27.Q_N a_4855_4775# VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X183 a_3984_5167# a_3453_4801# a_3900_5167# VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X184 a_8791_3239# a_8402_3239# a_8683_3605# VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X185 a_11089_4112# x4.X.t39 VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X186 a_5991_2340# a_6546_2340# a_6504_2648# VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X187 a_11075_3605# a_10794_3239# a_10982_3239# VDD.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X188 VDD.t428 check[0].t3 a_5372_4112# VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X189 VDD.t307 a_11629_2340# a_11628_2640# VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X190 a_9638_3213# a_9464_3239# a_9754_3239# VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X191 a_5088_3521# a_4680_3239# a_4854_3213# VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X192 x4.X.t12 a_1511_4112# VDD.t377 VDD.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X193 VDD.t177 VDD.t175 a_9442_4086# VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X194 a_6984_2366# a_6844_2640# a_6546_2340# VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X195 VDD.t450 x4.X.t40 a_4367_3213# VDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X196 VDD.t714 a_929_3238# x7.X VDD.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 a_7318_4296# a_6846_4086# a_7562_4478# VDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X198 VSS.t37 a_9441_2340# a_9376_2366# VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X199 a_4318_5083# a_3900_5167# a_4074_4775# VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X200 check[4].t0 a_10346_4801# VDD.t242 VDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X201 VDD.t375 a_1511_4112# x4.X.t11 VDD.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X202 a_12548_4112# a_11629_4386# a_12102_4296# VDD.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_12101_2550# a_11629_2340# a_12345_2732# VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X204 VSS.t64 x5.X.t10 a_3453_4801# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X205 a_11250_4775# VDD.t172 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X206 a_4453_2340# D[5].t2 VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X207 a_3373_5674# a_3258_5648# a_2389_5648# VDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X208 VSS.t17 x4.X.t41 a_6759_3213# VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X209 VSS.t217 reset.t1 a_621_4112# VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X210 a_1762_2340# a_2061_2340# a_1996_2366# VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X211 a_9550_3605# a_8402_3239# a_9464_3239# VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X212 a_8998_4801# VDD.t747 VSS.t166 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X213 x4.X.t29 a_1511_4112# VSS.t352 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 a_7049_2340# a_7317_2550# a_7263_2648# VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X215 a_6198_3239# x7.X VDD.t652 VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X216 VSS.t617 x7.X a_7763_2366# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X217 a_2398_4801# a_1061_4801# a_2289_4801# VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X218 VSS.t282 a_11629_2340# a_11628_2640# VSS.t281 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X219 VDD.t622 a_6759_3213# a_7480_3521# VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X220 a_3877_5674# a_2853_5648# a_3373_5674# VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X221 a_9656_4394# a_8697_4112# VDD.t440 VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X222 a_7185_2366# a_7317_2550# a_7049_2340# VSS.t287 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X223 a_10155_2366# a_9237_2340# a_9709_2550# VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X224 a_1926_5083# a_1508_5167# a_1682_4775# VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X225 a_9370_4801# a_8858_4775# VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X226 VDD.t171 VDD.t169 a_11834_4086# VDD.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X227 a_3504_2340# a_3599_2340# VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X228 a_11076_5167# a_10795_4801# a_10983_4801# VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X229 a_8792_4801# a_8403_4801# a_8684_5167# VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X230 a_5089_5083# a_4681_4801# a_4855_4775# VDD.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X231 x4.X.t28 a_1511_4112# VSS.t350 VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X232 VDD.t532 a_2061_2340# a_2060_2640# VDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X233 a_3671_5674# x48.Q VSS.t284 VSS.t283 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0819 ps=0.81 w=0.42 l=0.15
X234 a_4453_2340# D[5].t3 VSS.t387 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X235 a_4657_2340# a_4925_2550# a_4871_2648# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X236 a_3806_3239# VSS.t693 VDD.t581 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X237 x5.X.t6 a_1338_5674# VSS.t181 VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X238 a_9639_4775# a_9465_4801# a_9755_4801# VSS.t599 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X239 VDD.t269 a_12030_3213# a_12737_3239# VDD.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X240 a_4970_3239# a_4367_3213# a_4854_3213# VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X241 a_8857_3213# a_8683_3605# a_8997_3239# VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X242 a_3600_4086# a_4155_4086# a_4113_4394# VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X243 a_8383_2340# a_8696_2366# a_8802_2366# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X244 VDD.t500 a_6465_3213# a_6375_3605# VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X245 VSS.t492 check[0].t4 a_3877_5674# VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.066 ps=0.745 w=0.42 l=0.15
X246 VSS.t207 a_2463_4775# a_2398_4801# VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X247 VSS.t96 a_8289_4086# check[1].t0 VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X248 x5.A a_1062_5674# VDD.t563 VDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X249 VDD.t519 check[0].t5 a_3876_6040# VDD.t518 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0974 ps=0.97 w=0.64 l=0.15
X250 a_11390_4801# VDD.t748 VSS.t164 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X251 VSS.t215 a_5991_2340# x57.Q_N VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X252 a_4590_2732# a_4453_2340# a_4154_2340# VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X253 VDD.t222 a_8288_2340# D[4].t0 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X254 VSS.t615 x7.X a_10155_2366# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X255 a_9953_2732# a_9441_2340# VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X256 a_8289_4086# a_8384_4086# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X257 a_2697_5083# a_2289_4801# a_2463_4775# VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X258 a_9551_5167# a_8403_4801# a_9465_4801# VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X259 a_9441_2340# a_8696_2366# a_9577_2366# VSS.t521 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X260 a_6199_4801# check[6].t3 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X261 a_11630_4086# x5.X.t11 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X262 VSS.t19 x4.X.t42 a_6760_4775# VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X263 a_5170_4112# a_4658_4086# VSS.t486 VSS.t485 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X264 a_10680_2340# a_10775_2340# VSS.t467 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X265 VSS.t7 sel_bit[1].t0 a_3258_5648# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.113 ps=1.38 w=0.42 l=0.15
X266 a_9173_4478# a_8384_4086# VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X267 VDD.t5 sel_bit[1].t1 a_3258_5648# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X268 check[6].t0 a_5562_4801# VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X269 VDD.t547 a_6760_4775# a_7481_5083# VDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X270 a_4389_4112# a_3600_4086# VSS.t520 VSS.t519 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X271 a_5372_4112# a_4454_4086# a_4926_4296# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X272 a_9375_4478# a_9238_4086# a_8939_4086# VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X273 VSS.t504 a_2061_2340# a_2060_2640# VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_6465_3213# a_6291_3605# a_6605_3239# VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X275 VSS.t49 a_5897_4086# check[0].t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X276 a_6399_3239# a_6010_3239# a_6291_3605# VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X277 VSS.t46 a_3599_2340# x54.Q_N VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X278 eob.t3 a_2389_5648# VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X279 VDD.t694 x5.X.t12 a_1061_4801# VDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X280 VDD.t340 a_5896_2340# D[5].t0 VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X281 VDD.t387 x27.Q_N a_3599_2340# VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X282 a_11389_3239# a_11543_3213# a_11249_3213# VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X283 VDD.t513 a_4658_4086# a_4591_4478# VDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X284 VDD.t528 a_9237_2340# a_9236_2640# VDD.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X285 a_5897_4086# a_5992_4086# VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X286 a_8289_4086# a_8384_4086# VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X287 a_6304_2366# x4.X.t43 VSS.t405 VSS.t404 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X288 a_3807_4801# x27.D VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X289 a_12146_3239# x39.Q_N VSS.t94 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X290 VSS.t246 a_12031_4775# a_12738_4801# VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X291 a_6781_4478# a_5992_4086# VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X292 VSS.t637 a_1112_2340# D[7].t1 VSS.t636 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X293 a_12146_3239# a_11543_3213# a_12030_3213# VSS.t557 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X294 a_6983_4478# a_6846_4086# a_6547_4086# VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X295 VDD.t168 VDD.t166 a_8384_4086# VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X296 a_9238_4086# x5.X.t13 VDD.t696 VDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X297 a_12047_2648# a_11088_2366# VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X298 a_6546_2340# a_6844_2640# a_6780_2732# VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X299 a_1520_2366# x4.X.t44 VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X300 a_4585_3239# a_4073_3213# VSS.t86 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X301 VDD.t329 a_6466_4775# a_6376_5167# VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X302 VSS.t104 a_7049_2340# a_6984_2366# VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X303 a_11564_2732# a_10775_2340# VDD.t494 VDD.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X304 x4.X.t10 a_1511_4112# VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X305 a_11766_2732# a_11629_2340# a_11330_2340# VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 a_11833_2340# a_11088_2366# a_11969_2366# VSS.t188 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X307 a_4971_4801# a_4368_4775# a_4855_4775# VSS.t400 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X308 a_4155_4086# a_4454_4086# a_4389_4112# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X309 a_10156_4112# a_9237_4386# a_9710_4296# VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X310 a_7072_3239# a_6010_3239# a_6977_3239# VSS.t254 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X311 a_4007_3239# a_3618_3239# a_3899_3605# VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X312 a_8858_4775# a_8684_5167# a_8998_4801# VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X313 x4.X.t27 a_1511_4112# VSS.t348 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X314 VDD.t293 x4.X.t45 a_11544_4775# VDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X315 a_6305_4112# x4.X.t46 VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X316 a_4018_2366# a_4154_2340# a_3599_2340# VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X317 a_5897_4086# a_5992_4086# VSS.t409 VSS.t408 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X318 VDD.t263 a_12031_4775# a_12738_4801# VDD.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X319 a_3912_2366# x4.X.t47 VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X320 a_7158_3605# a_6010_3239# a_7072_3239# VDD.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X321 a_12346_4112# a_11834_4086# VSS.t362 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X322 a_9578_4112# a_9710_4296# a_9442_4086# VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X323 a_12548_4112# a_11630_4086# a_12102_4296# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X324 VDD.t15 a_8384_4086# x42.Q_N VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X325 VSS.t500 a_9237_2340# a_9236_2640# VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X326 a_4925_2550# a_4452_2640# a_5169_2366# VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X327 VDD.t165 VDD.t163 a_5992_4086# VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X328 x4.A a_897_4112# VSS.t566 VSS.t565 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 VSS.t124 a_4657_2340# a_4592_2366# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X330 x5.A a_1062_5674# VSS.t526 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X331 x4.X.t26 a_1511_4112# VSS.t346 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X332 a_2579_4801# a_1976_4775# a_2463_4775# VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X333 VDD.t734 x36.Q_N a_10775_2340# VDD.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X334 a_4680_3239# a_3618_3239# a_4585_3239# VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X335 a_6466_4775# a_6292_5167# a_6606_4801# VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X336 VDD.t575 x4.A a_1511_4112# VDD.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X337 a_3913_4112# x4.X.t48 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X338 a_1626_2366# a_1762_2340# a_1207_2340# VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X339 VSS.t35 a_9638_3213# a_10345_3239# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X340 VDD.t313 a_9151_3213# a_9101_3521# VDD.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X341 a_1112_2340# a_1207_2340# VDD.t587 VDD.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X342 a_11390_4801# a_11544_4775# a_11250_4775# VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X343 VSS.t641 a_6846_4086# a_6845_4386# VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X344 a_4766_3605# a_3618_3239# a_4680_3239# VDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X345 VDD.t3 a_11630_4086# a_11629_4386# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X346 x75.Q_N a_4854_3213# VSS.t58 VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X347 a_2533_2550# a_2060_2640# a_2777_2366# VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X348 a_2401_2366# a_2533_2550# a_2265_2340# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X349 a_12147_4801# VDD.t749 VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X350 VSS.t82 check[3].t2 a_12548_4112# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X351 a_12147_4801# a_11544_4775# a_12031_4775# VSS.t446 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X352 a_10982_3239# x7.X VSS.t613 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X353 a_4586_4801# a_4074_4775# VSS.t550 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X354 a_2198_2732# a_2061_2340# a_1762_2340# VDD.t530 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X355 a_8857_3213# x42.Q_N VDD.t517 VDD.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X356 a_8403_4801# a_8237_4801# VDD.t708 VDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X357 a_4008_4801# a_3619_4801# a_3900_5167# VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X358 a_7073_4801# a_6011_4801# a_6978_4801# VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X359 x66.Q_N a_12030_3213# VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X360 VDD.t620 a_6759_3213# a_6709_3521# VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X361 a_7159_5167# a_6011_4801# a_7073_4801# VDD.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X362 a_4454_4086# x5.X.t14 VDD.t688 VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X363 VSS.t73 a_4454_4086# a_4453_4386# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X364 a_8897_4394# a_8697_4112# VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X365 a_12030_3213# x39.Q_N VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X366 D[1].t1 a_10345_3239# VSS.t626 VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X367 VDD.t561 x5.A a_1338_5674# VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X368 a_3373_5674# a_2853_5648# a_3648_5972# VDD.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.164 ps=1.33 w=0.42 l=0.15
X369 a_11331_4086# a_11629_4386# a_11565_4478# VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X370 a_11856_3239# a_10794_3239# a_11761_3239# VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X371 a_8697_4112# x4.X.t49 VSS.t633 VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X372 a_8683_3605# a_8402_3239# a_8590_3239# VDD.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X373 D[0].t1 a_7953_3239# VDD.t468 VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X374 a_6011_4801# a_5845_4801# VDD.t736 VDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X375 VSS.t681 x36.Q_N a_11969_2366# VSS.t680 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X376 a_4681_4801# a_3619_4801# a_4586_4801# VSS.t477 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X377 VDD.t136 a_9152_4775# a_9102_5083# VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X378 VSS.t128 a_3505_4086# x48.Q VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X379 a_4767_5167# a_3619_4801# a_4681_4801# VDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X380 x4.X.t25 a_1511_4112# VSS.t344 VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X381 VSS.t160 VDD.t750 a_1976_4775# VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X382 a_5170_4478# a_4658_4086# VDD.t511 VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X383 a_4112_2648# a_3912_2366# VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X384 VDD.t742 a_3504_2340# D[6].t0 VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X385 VSS.t309 a_9639_4775# a_10346_4801# VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X386 a_2463_4775# x4.X.t50 VDD.t672 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X387 a_3505_4086# a_3600_4086# VDD.t555 VDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X388 a_4389_4478# a_3600_4086# VDD.t553 VDD.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X389 VDD.t650 x7.X a_7763_2366# VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X390 VSS.t659 a_929_3238# x7.X VSS.t658 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X391 VSS.t393 a_2389_5648# eob.t0 VSS.t392 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X392 VDD.t536 a_1976_4775# a_2697_5083# VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X393 x4.A a_897_4112# VSS.t564 VSS.t563 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X394 x27.Q_N a_4855_4775# VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X395 a_6411_4112# a_6547_4086# a_5992_4086# VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X396 VDD.t573 x4.A a_1511_4112# VDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X397 a_8858_4775# VDD.t160 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X398 a_10983_4801# check[4].t2 VSS.t669 VSS.t668 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X399 VDD.t545 a_6760_4775# a_6710_5083# VDD.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X400 a_7318_4296# a_6845_4386# a_7562_4112# VSS.t457 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X401 VDD.t338 a_9639_4775# a_10346_4801# VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X402 a_12031_4775# VDD.t157 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X403 a_1720_2648# a_1520_2366# VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X404 VSS.t84 a_4073_3213# a_4007_3239# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X405 a_3505_4086# a_3600_4086# VSS.t518 VSS.t517 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X406 VSS.t33 a_9638_3213# a_9573_3239# VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X407 a_2289_4801# a_1061_4801# a_2147_5083# VDD.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X408 a_6845_2340# D[4].t2 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X409 VDD.t226 a_2463_4775# a_2375_5167# VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X410 a_7561_2366# a_7049_2340# VSS.t102 VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X411 a_7763_2366# a_6845_2340# a_7317_2550# VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X412 check[4].t1 a_10346_4801# VSS.t221 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X413 VDD.t371 a_1511_4112# x4.X.t9 VDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 VDD.t27 a_9441_2340# a_9374_2732# VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X415 VSS.t158 VDD.t751 a_7186_4112# VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X416 a_8684_5167# a_8403_4801# a_8591_4801# VDD.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X417 a_11857_4801# a_10795_4801# a_11762_4801# VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X418 VDD.t648 x7.X a_10155_2366# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X419 a_8938_2340# a_9237_2340# a_9172_2366# VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X420 a_6930_3521# a_6465_3213# VDD.t498 VDD.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X421 VDD.t599 a_897_4112# x4.A VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X422 a_3600_4086# a_3913_4112# a_4019_4112# VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X423 a_1511_4112# x4.A VSS.t536 VSS.t535 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X424 VSS.t156 VDD.t752 a_4019_4112# VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X425 a_12346_4478# a_11834_4086# VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X426 a_11288_2648# a_11088_2366# VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X427 x75.Q a_5561_3239# VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X428 x77.Y eob.t9 VSS.t399 VSS.t398 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X429 VDD.t346 a_9238_4086# a_9237_4386# VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X430 a_11493_3521# a_11075_3605# a_11249_3213# VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X431 a_3373_5674# sel_bit[1].t2 a_2389_5648# VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X432 VDD.t551 a_3600_4086# x48.Q_N VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X433 a_9710_4296# a_9237_4386# a_9954_4112# VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X434 a_6845_2340# D[4].t3 VSS.t380 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X435 x4.X.t24 a_1511_4112# VSS.t342 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X436 a_6546_2340# a_6845_2340# a_6780_2366# VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X437 VSS.t250 a_12030_3213# a_11965_3239# VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X438 a_11075_3605# a_10628_3239# a_10982_3239# VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X439 x69.Q_N a_9638_3213# VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X440 a_1415_4801# eob.t10 VSS.t397 VSS.t396 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X441 VSS.t317 a_11249_3213# a_11183_3239# VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X442 VDD.t690 x5.X.t15 a_10629_4801# VDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X443 x36.Q_N a_12031_4775# VDD.t261 VDD.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X444 VSS.t657 a_929_3238# x7.X VSS.t656 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X445 a_5371_2366# a_4452_2640# a_4925_2550# VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 VSS.t548 a_4074_4775# a_4008_4801# VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X447 a_2993_5674# sel_bit[0].t0 a_2883_5674# VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.072 ps=0.76 w=0.36 l=0.15
X448 VDD.t74 check[3].t3 a_12548_4112# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X449 VSS.t71 a_10680_2340# D[3].t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X450 VDD.t571 x4.A a_1511_4112# VDD.t570 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X451 VSS.t340 a_1511_4112# x4.X.t23 VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X452 a_12264_3521# a_11856_3239# a_12030_3213# VDD.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X453 VSS.t307 a_9639_4775# a_9574_4801# VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X454 VSS.t391 a_2389_5648# eob.t7 VSS.t390 sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X455 VSS.t179 a_1338_5674# x5.X.t5 VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X456 a_6931_5083# a_6466_4775# VDD.t327 VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X457 a_10776_4086# a_11089_4112# a_11195_4112# VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X458 VDD.t50 x4.X.t51 a_11543_3213# VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X459 a_3619_4801# a_3453_4801# VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X460 VSS.t154 VDD.t753 a_11195_4112# VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X461 a_2289_4801# a_1227_4801# a_2194_4801# VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X462 check[5].t0 a_7954_4801# VDD.t452 VDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X463 a_11494_5083# a_11076_5167# a_11250_4775# VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X464 VDD.t385 x27.Q_N a_4657_2340# VDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X465 a_2979_2366# a_2060_2640# a_2533_2550# VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X466 a_11159_3605# a_10628_3239# a_11075_3605# VDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X467 check[6].t1 a_5562_4801# VSS.t667 VSS.t666 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X468 VDD.t702 a_7050_4086# a_6983_4478# VDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X469 a_9754_3239# x42.Q_N VSS.t488 VSS.t487 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X470 a_1508_5167# a_1061_4801# a_1415_4801# VSS.t479 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X471 a_9754_3239# a_9151_3213# a_9638_3213# VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X472 VSS.t368 a_1682_4775# a_1616_4801# VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X473 a_9655_2648# a_8696_2366# VDD.t559 VDD.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X474 VDD.t369 a_1511_4112# x4.X.t8 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X475 a_8384_4086# a_8939_4086# a_8897_4394# VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X476 x7.A a_653_3238# VSS.t570 VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X477 a_6605_3239# x45.Q_N VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X478 a_7764_4112# a_6845_4386# a_7318_4296# VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X479 a_3899_3605# a_3618_3239# a_3806_3239# VDD.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X480 a_8938_2340# a_9236_2640# a_9172_2732# VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X481 a_12547_2366# a_11628_2640# a_12101_2550# VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X482 a_9954_4112# a_9442_4086# VSS.t259 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X483 x20.Q_N a_2463_4775# VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X484 a_11076_5167# a_10629_4801# a_10983_4801# VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X485 VSS.t244 a_12031_4775# a_11966_4801# VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X486 VDD.t367 a_1511_4112# x4.X.t7 VDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X487 VDD.t106 x20.Q_N a_2265_2340# VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X488 a_1592_5167# a_1061_4801# a_1508_5167# VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X489 a_8696_2366# x4.X.t52 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X490 a_10680_2340# a_10775_2340# VDD.t492 VDD.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X491 a_5169_2366# a_4657_2340# VSS.t122 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X492 a_3599_2340# a_4154_2340# a_4112_2648# VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X493 a_12265_5083# a_11857_4801# a_12031_4775# VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X494 a_10982_3239# x7.X VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X495 a_7246_3213# a_7072_3239# a_7362_3239# VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X496 VDD.t661 x3.A a_897_4112# VDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X497 VDD.t156 VDD.t154 a_7050_4086# VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X498 VDD.t454 x7.A a_929_3238# VDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X499 a_4592_2366# a_4452_2640# a_4154_2340# VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X500 a_8402_3239# a_8236_3239# VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X501 a_4538_3521# a_4073_3213# VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X502 a_4926_4296# a_4454_4086# a_5170_4478# VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X503 a_10776_4086# a_11331_4086# a_11289_4394# VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X504 VDD.t732 x36.Q_N a_11833_2340# VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X505 a_9709_2550# a_9237_2340# a_9953_2732# VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X506 a_2061_2340# D[6].t2 VDD.t632 VDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X507 VSS.t643 x5.X.t16 a_1061_4801# VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X508 a_2777_2366# a_2265_2340# VSS.t225 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X509 a_1207_2340# a_1762_2340# a_1720_2648# VDD.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X510 a_9755_4801# VDD.t754 VSS.t152 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X511 a_2979_2366# a_2061_2340# a_2533_2550# VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X512 VSS.t528 x4.X.t53 a_4367_3213# VSS.t527 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X513 VSS.t177 a_1338_5674# x5.X.t4 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X514 a_9755_4801# a_9152_4775# a_9639_4775# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X515 a_6606_4801# VDD.t755 VSS.t150 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X516 a_11565_4112# a_10776_4086# VSS.t441 VSS.t440 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X517 a_8802_2366# a_8938_2340# a_8383_2340# VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X518 a_11088_2366# x4.X.t54 VDD.t565 VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X519 VSS.t611 x7.X a_5371_2366# VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X520 VDD.t122 a_4657_2340# a_4590_2732# VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X521 a_6010_3239# a_5844_3239# VDD.t609 VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X522 VDD.t640 a_4367_3213# a_5088_3521# VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X523 a_7264_4394# a_6305_4112# VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X524 a_8402_3239# a_8236_3239# VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 VSS.t583 x33.Q_N a_8802_2366# VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X526 a_9638_3213# x42.Q_N VDD.t515 VDD.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X527 VDD.t365 a_1511_4112# x4.X.t6 VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X528 VSS.t465 a_10775_2340# x63.Q_N VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X529 x4.X.t22 a_1511_4112# VSS.t338 VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X530 a_11834_4086# a_12102_4296# a_12048_4394# VDD.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X531 a_3648_5972# x48.Q VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0864 ps=0.91 w=0.64 l=0.15
X532 a_6400_4801# a_6011_4801# a_6292_5167# VSS.t384 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X533 a_10983_4801# check[4].t3 VDD.t722 VDD.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X534 a_6846_4086# x5.X.t17 VDD.t692 VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X535 a_11768_2366# a_11628_2640# a_11330_2340# VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X536 a_2061_2340# D[6].t3 VSS.t595 VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X537 a_4539_5083# a_4074_4775# VDD.t585 VDD.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X538 a_2265_2340# a_2533_2550# a_2479_2648# VDD.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X539 a_6605_3239# a_6759_3213# a_6465_3213# VSS.t585 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X540 a_7247_4775# a_7073_4801# a_7363_4801# VSS.t598 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X541 a_12102_4296# a_11630_4086# a_12346_4478# VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X542 a_11761_3239# a_11249_3213# VSS.t315 VSS.t314 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X543 VSS.t581 x33.Q_N a_9577_2366# VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X544 VDD.t23 a_9638_3213# a_10345_3239# VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X545 VDD.t363 a_1511_4112# x4.X.t5 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X546 a_4872_4394# a_3913_4112# VDD.t238 VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X547 VSS.t21 a_8384_4086# x42.Q_N VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X548 a_11331_4086# a_11630_4086# a_11565_4112# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X549 VDD.t728 a_8383_2340# x60.Q_N VDD.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X550 a_5991_2340# a_6304_2366# a_6410_2366# VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X551 a_6010_3239# a_5844_3239# VSS.t572 VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X552 VDD.t76 a_4073_3213# a_3983_3605# VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X553 VSS.t591 x30.Q_N a_6410_2366# VSS.t590 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.12 ps=1.08 w=0.42 l=0.15
X554 a_9464_3239# a_8236_3239# a_9322_3521# VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X555 VDD.t21 a_9638_3213# a_9550_3605# VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X556 VDD.t597 a_897_4112# x4.A VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 VSS.t270 x4.X.t55 a_11543_3213# VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X558 a_11194_2366# a_11330_2340# a_10775_2340# VSS.t458 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X559 a_7561_2732# a_7049_2340# VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X560 a_9377_4112# a_9237_4386# a_8939_4086# VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X561 VSS.t534 x4.A a_1511_4112# VSS.t533 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X562 a_7049_2340# a_6304_2366# a_7185_2366# VSS.t186 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X563 VSS.t272 x4.X.t56 a_4368_4775# VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X564 a_9238_4086# x5.X.t18 VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X565 a_12101_2550# a_11628_2640# a_12345_2366# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X566 x5.X.t1 a_1338_5674# VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X567 eob.t2 a_2389_5648# VDD.t414 VDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X568 VDD.t595 a_11543_3213# a_12264_3521# VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X569 x27.D a_3170_4801# VDD.t718 VDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X570 VDD.t422 a_4368_4775# a_5089_5083# VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X571 VDD.t361 a_1511_4112# x4.X.t4 VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X572 a_11969_2366# a_12101_2550# a_11833_2340# VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X573 VSS.t451 a_11833_2340# a_11768_2366# VSS.t450 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X574 a_4073_3213# a_3899_3605# a_4213_3239# VSS.t587 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X575 a_9639_4775# VDD.t151 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X576 VSS.t132 a_7246_3213# a_7953_3239# VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X577 VSS.t554 a_1207_2340# x51.Q_N VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X578 a_8403_4801# a_8237_4801# VSS.t655 VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X579 a_6985_4112# a_6845_4386# a_6547_4086# VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X580 a_9573_3239# a_8236_3239# a_9464_3239# VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X581 a_11942_3605# a_10794_3239# a_11856_3239# VDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X582 a_4854_3213# a_4680_3239# a_4970_3239# VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X583 a_4657_2340# a_3912_2366# a_4793_2366# VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X584 x66.Q_N a_12030_3213# VSS.t248 VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X585 a_1415_4801# eob.t11 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X586 VSS.t257 a_9442_4086# a_9377_4112# VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X587 VDD.t265 a_12030_3213# a_11942_3605# VDD.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X588 a_4591_4478# a_4454_4086# a_4155_4086# VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X589 a_4154_2340# a_4452_2640# a_4388_2732# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X590 VDD.t523 D[1].t2 a_10628_3239# VDD.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X591 a_9954_4478# a_9442_4086# VDD.t274 VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X592 VDD.t7 a_10681_4086# check[2].t0 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X593 a_8896_2648# a_8696_2366# VDD.t557 VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X594 VDD.t342 a_11249_3213# a_11159_3605# VDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X595 VDD.t583 a_4074_4775# a_3984_5167# VDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X596 a_11762_4801# a_11250_4775# VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X597 a_9322_3521# a_8857_3213# VDD.t448 VDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X598 a_9172_2366# a_8383_2340# VSS.t677 VSS.t676 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X599 a_9465_4801# a_8237_4801# a_9323_5083# VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X600 VSS.t56 a_4854_3213# a_5561_3239# VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X601 VDD.t336 a_9639_4775# a_9551_5167# VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X602 a_6011_4801# a_5845_4801# VSS.t685 VSS.t684 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X603 VDD.t13 x4.X.t57 a_9152_4775# VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X604 VSS.t228 check[1].t4 a_7764_4112# VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X605 D[0].t0 a_7953_3239# VSS.t445 VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X606 VSS.t15 x4.X.t58 a_11544_4775# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X607 VSS.t3 a_11630_4086# a_11629_4386# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X608 a_1520_2366# x4.X.t59 VSS.t27 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X609 VDD.t282 clk_sar.t0 a_1062_5674# VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X610 a_7186_4112# a_7318_4296# a_7050_4086# VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X611 a_10156_4112# a_9238_4086# a_9710_4296# VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X612 VDD.t472 a_11544_4775# a_12265_5083# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X613 a_3618_3239# a_3452_3239# VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X614 VDD.t430 a_5992_4086# x45.Q_N VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X615 a_8683_3605# a_8236_3239# a_8590_3239# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X616 VDD.t150 VDD.t148 a_3600_4086# VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X617 a_11249_3213# a_11075_3605# a_11389_3239# VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X618 x72.Q_N a_7246_3213# VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X619 VSS.t427 a_8857_3213# a_8791_3239# VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X620 VDD.t393 a_1682_4775# a_1592_5167# VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X621 x3.A a_621_4112# VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X622 a_6780_2366# a_5991_2340# VSS.t213 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X623 VSS.t223 a_2265_2340# a_2200_2366# VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X624 VSS.t568 comparator_out.t0 a_653_3238# VSS.t567 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X625 a_4074_4775# a_3900_5167# a_4214_4801# VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X626 VSS.t496 D[1].t3 a_10628_3239# VSS.t495 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X627 VSS.t532 x4.A a_1511_4112# VSS.t531 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X628 a_4454_4086# x5.X.t19 VSS.t140 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X629 VSS.t291 a_7247_4775# a_7954_4801# VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X630 a_6547_4086# a_6845_4386# a_6781_4478# VDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X631 a_10681_4086# a_10776_4086# VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X632 a_11943_5167# a_10795_4801# a_11857_4801# VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X633 a_11088_2366# x4.X.t60 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X634 a_9872_3521# a_9464_3239# a_9638_3213# VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X635 x5.X.t0 a_1338_5674# VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X636 a_3876_6040# sel_bit[0].t1 a_3373_5674# VDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.0974 pd=0.97 as=0.0567 ps=0.69 w=0.42 l=0.15
X637 a_11565_4478# a_10776_4086# VDD.t462 VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X638 VDD.t359 a_1511_4112# x4.X.t3 VDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X639 a_4794_4112# a_4926_4296# a_4658_4086# VSS.t262 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X640 a_4855_4775# a_4681_4801# a_4971_4801# VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X641 a_9574_4801# a_8237_4801# a_9465_4801# VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X642 a_8384_4086# a_8697_4112# a_8803_4112# VSS.t420 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X643 a_11767_4478# a_11630_4086# a_11331_4086# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X644 VDD.t259 a_12031_4775# a_11943_5167# VDD.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X645 x36.Q_N a_12031_4775# VSS.t242 VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X646 D[2].t0 a_12737_3239# VDD.t642 VDD.t641 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X647 a_9323_5083# a_8858_4775# VDD.t480 VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X648 VSS.t88 check[2].t4 a_10156_4112# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X649 VDD.t232 a_5991_2340# x57.Q_N VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X650 a_8767_3605# a_8236_3239# a_8683_3605# VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X651 a_3618_3239# a_3452_3239# VSS.t377 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X652 a_2194_4801# a_1682_4775# VSS.t366 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X653 a_1682_4775# a_1508_5167# a_1822_4801# VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X654 VDD.t318 a_7247_4775# a_7954_4801# VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X655 VSS.t336 a_1511_4112# x4.X.t21 VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X656 a_5169_2732# a_4657_2340# VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X657 a_6465_3213# x45.Q_N VDD.t251 VDD.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X658 VSS.t110 a_4855_4775# a_5562_4801# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X659 a_10681_4086# a_10776_4086# VSS.t439 VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X660 a_1616_4801# a_1227_4801# a_1508_5167# VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X661 VDD.t638 a_4367_3213# a_4317_3521# VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X662 VSS.t562 a_897_4112# x4.A VSS.t561 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X663 x7.A a_653_3238# VDD.t607 VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X664 a_6505_4394# a_6305_4112# VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.218 ps=2.2 w=0.84 l=0.15
X665 a_9709_2550# a_9236_2640# a_9953_2366# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X666 a_2463_4775# a_2289_4801# a_2579_4801# VSS.t624 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
X667 check[5].t1 a_7954_4801# VSS.t431 VSS.t430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X668 VDD.t147 VDD.t145 a_10776_4086# VDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X669 a_1511_4112# x4.A VDD.t569 VDD.t568 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X670 VSS.t516 a_3600_4086# x48.Q_N VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X671 VDD.t32 a_3599_2340# x54.Q_N VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X672 a_1207_2340# a_1520_2366# a_1626_2366# VSS.t460 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X673 a_8684_5167# a_8237_4801# a_8591_4801# VSS.t652 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X674 VSS.t453 a_8858_4775# a_8792_4801# VSS.t452 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X675 VDD.t100 a_4855_4775# a_5562_4801# VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X676 a_6305_4112# x4.X.t61 VSS.t372 VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X677 a_3373_5674# sel_bit[0].t2 a_3671_5674# VSS.t508 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0671 ps=0.75 w=0.36 l=0.15
X678 a_2777_2732# a_2265_2340# VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0798 ps=0.8 w=0.42 l=0.15
X679 a_6291_3605# a_6010_3239# a_6198_3239# VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X680 a_2883_5674# sel_bit[0].t3 a_2784_5996# VDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.105 ps=0.995 w=0.42 l=0.15
X681 a_9873_5083# a_9465_4801# a_9639_4775# VDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X682 VSS.t589 x5.X.t20 a_10629_4801# VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X683 a_11629_2340# D[2].t2 VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X684 VSS.t1 clk_sar.t1 a_1062_5674# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X685 a_2375_5167# a_1227_4801# a_2289_4801# VDD.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X686 VDD.t678 a_1112_2340# D[7].t0 VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X687 x69.Q_N a_9638_3213# VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X688 VDD.t460 a_10776_4086# x39.Q_N VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X689 a_11834_4086# a_11089_4112# a_11970_4112# VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X690 VDD.t644 x7.X a_5371_2366# VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X691 x20.Q_N a_2463_4775# VSS.t205 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X692 VDD.t626 x5.X.t21 a_8237_4801# VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X693 x3.A a_621_4112# VSS.t193 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X694 VDD.t618 x33.Q_N a_9441_2340# VDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X695 a_8768_5167# a_8237_4801# a_8684_5167# VDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X696 a_6709_3521# a_6291_3605# a_6465_3213# VDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X697 a_4019_4112# a_4155_4086# a_3600_4086# VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X698 x7.X a_929_3238# VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 VSS.t530 x4.A a_1511_4112# VSS.t529 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X700 a_7317_2550# a_6845_2340# a_7561_2732# VDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X701 a_6466_4775# VDD.t142 VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X702 a_3913_4112# x4.X.t62 VSS.t374 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X703 a_3619_4801# a_3453_4801# VSS.t276 VSS.t275 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X704 VSS.t203 a_8288_2340# D[4].t1 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X705 VDD.t593 a_11543_3213# a_11493_3521# VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X706 a_4926_4296# a_4453_4386# a_5170_4112# VSS.t418 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X707 VSS.t320 a_9238_4086# a_9237_4386# VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X708 a_4789_3239# a_3452_3239# a_4680_3239# VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X709 VDD.t420 a_4368_4775# a_4318_5083# VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X710 VSS.t510 a_11250_4775# a_11184_4801# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X711 VSS.t484 a_4658_4086# a_4593_4112# VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0935 ps=0.965 w=0.64 l=0.15
X712 a_11629_2340# D[2].t3 VSS.t274 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X713 VSS.t130 a_7246_3213# a_7181_3239# VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X714 VDD.t684 x5.X.t22 a_5845_4801# VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X715 x30.Q_N a_7247_4775# VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X716 VDD.t94 a_7049_2340# a_6982_2732# VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X717 a_5371_2366# a_4453_2340# a_4925_2550# VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X718 a_4388_2366# a_3599_2340# VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X719 VSS.t334 a_1511_4112# x4.X.t20 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X720 VSS.t148 VDD.t756 a_4794_4112# VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X721 a_8383_2340# a_8938_2340# a_8896_2648# VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X722 a_10795_4801# a_10629_4801# VDD.t286 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X723 VDD.t466 check[1].t5 a_7764_4112# VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X724 a_9442_4086# a_9710_4296# a_9656_4394# VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X725 a_6292_5167# a_6011_4801# a_6199_4801# VDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X726 VSS.t313 a_5896_2340# D[5].t1 VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X727 eob.t6 a_2389_5648# VSS.t389 VSS.t388 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.218 ps=1.97 w=0.65 l=0.15
X728 VDD.t534 a_1976_4775# a_1926_5083# VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X729 a_11160_5167# a_10629_4801# a_11076_5167# VDD.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X730 a_1511_4112# x4.A VDD.t567 VDD.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X731 a_8288_2340# a_8383_2340# VSS.t675 VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X732 VSS.t54 a_4854_3213# a_4789_3239# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X733 VSS.t332 a_1511_4112# x4.X.t19 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X734 a_1996_2366# a_1207_2340# VSS.t552 VSS.t551 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0588 ps=0.7 w=0.42 l=0.15
X735 check[3].t0 a_12738_4801# VDD.t458 VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X736 a_4073_3213# x77.Y VDD.t668 VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X737 a_8997_3239# a_9151_3213# a_8857_3213# VSS.t285 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X738 a_3900_5167# a_3619_4801# a_3807_4801# VDD.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X739 VDD.t470 a_11544_4775# a_11494_5083# VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X740 a_4154_2340# a_4453_2340# a_4388_2366# VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X741 VSS.t622 x3.A a_897_4112# VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X742 VDD.t324 a_6845_2340# a_6844_2640# VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X743 VSS.t433 x7.A a_929_3238# VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X744 x33.Q_N a_9639_4775# VDD.t334 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X745 a_9441_2340# a_9709_2550# a_9655_2648# VDD.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X746 VDD.t389 a_11834_4086# a_11767_4478# VDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X747 a_5896_2340# a_5991_2340# VSS.t211 VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X748 VDD.t311 a_9151_3213# a_9872_3521# VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X749 a_10775_2340# a_11330_2340# a_11288_2648# VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X750 a_12345_2366# a_11833_2340# VSS.t449 VSS.t448 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X751 VDD.t114 check[2].t5 a_10156_4112# VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X752 a_9577_2366# a_9709_2550# a_9441_2340# VSS.t688 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0864 ps=0.91 w=0.64 l=0.15
X753 a_12547_2366# a_11629_2340# a_12101_2550# VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X754 x7.X a_929_3238# VDD.t710 VDD.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X755 VSS.t289 a_7247_4775# a_7182_4801# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X756 a_9172_2732# a_8383_2340# VDD.t726 VDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X757 VSS.t146 VDD.t757 a_11970_4112# VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.101 ps=0.99 w=0.42 l=0.15
X758 a_9374_2732# a_9237_2340# a_8938_2340# VDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X759 VDD.t297 x4.X.t63 a_9151_3213# VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X760 a_1227_4801# a_1061_4801# VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X761 x4.X.t2 a_1511_4112# VDD.t357 VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X762 VDD.t219 a_4453_2340# a_4452_2640# VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X763 a_2389_5648# sel_bit[1].t3 a_2883_5674# VDD.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X764 VDD.t412 a_2389_5648# eob.t1 VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X765 x27.D a_3170_4801# VSS.t665 VSS.t664 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X766 VSS.t296 a_6845_2340# a_6844_2640# VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X767 a_7362_3239# x45.Q_N VSS.t232 VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X768 a_7263_2648# a_6304_2366# VDD.t202 VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X769 a_7362_3239# a_6759_3213# a_7246_3213# VSS.t584 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X770 VSS.t330 a_1511_4112# x4.X.t18 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X771 a_5992_4086# a_6547_4086# a_6505_4394# VDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0882 ps=1.05 w=0.84 l=0.15
X772 VDD.t446 a_8857_3213# a_8767_3605# VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X773 a_4213_3239# x77.Y VSS.t631 VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X774 VSS.t108 a_4855_4775# a_4790_4801# VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X775 a_6780_2732# a_5991_2340# VDD.t230 VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0819 ps=0.81 w=0.42 l=0.15
X776 a_5372_4112# a_4453_4386# a_4926_4296# VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X777 VDD.t616 x33.Q_N a_8383_2340# VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X778 a_11833_2340# a_12101_2550# a_12047_2648# VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X779 a_6982_2732# a_6845_2340# a_6546_2340# VDD.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X780 a_4925_2550# a_4453_2340# a_5169_2732# VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X781 a_11330_2340# a_11629_2340# a_11564_2366# VSS.t279 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X782 VSS.t609 x7.X a_12547_2366# VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X783 VDD.t299 x4.X.t64 a_6760_4775# VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X784 a_8998_4801# a_9152_4775# a_8858_4775# VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X785 a_10155_2366# a_9236_2640# a_9709_2550# VDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X786 a_7562_4112# a_7050_4086# VSS.t649 VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.084 ps=0.82 w=0.42 l=0.15
X787 VDD.t134 a_9152_4775# a_9873_5083# VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X788 VSS.t328 a_1511_4112# x4.X.t17 VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X789 a_7764_4112# a_6846_4086# a_7318_4296# VSS.t639 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X790 VSS.t199 a_4453_2340# a_4452_2640# VSS.t198 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X791 a_6304_2366# x4.X.t65 VDD.t442 VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X792 a_9369_3239# a_8857_3213# VSS.t425 VSS.t424 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X793 a_4970_3239# x77.Y VSS.t629 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X794 a_4871_2648# a_3912_2366# VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.225 ps=1.38 w=0.84 l=0.15
X795 VSS.t524 x5.A a_1338_5674# VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X796 VSS.t560 a_897_4112# x4.A VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X797 a_8939_4086# a_9238_4086# a_9173_4112# VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X798 a_8590_3239# x7.X VSS.t607 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X799 VDD.t128 a_7246_3213# a_7953_3239# VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X800 VDD.t628 x30.Q_N a_5991_2340# VDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.123 ps=1.17 w=0.42 l=0.15
X801 a_2533_2550# a_2061_2340# a_2777_2732# VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0945 ps=0.87 w=0.42 l=0.15
X802 a_1682_4775# x4.X.t66 VDD.t444 VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X803 VDD.t686 x5.X.t23 a_3453_4801# VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X804 VDD.t141 VDD.t139 a_4658_4086# VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.147 ps=1.23 w=0.42 l=0.15
X805 a_7050_4086# a_7318_4296# a_7264_4394# VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X806 VDD.t605 comparator_out.t1 a_653_3238# VDD.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X807 x4.X.t1 a_1511_4112# VDD.t355 VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X808 a_2200_2366# a_2060_2640# a_1762_2340# VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.0711 ps=0.755 w=0.36 l=0.15
X809 a_2853_5648# sel_bit[0].t4 VDD.t405 VDD.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X810 a_2853_5648# sel_bit[0].t5 VSS.t382 VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X811 a_8696_2366# x4.X.t67 VSS.t403 VSS.t402 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X812 a_6606_4801# a_6760_4775# a_6466_4775# VSS.t514 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X813 VSS.t326 a_1511_4112# x4.X.t16 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X814 VSS.t691 a_3504_2340# D[6].t1 VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X815 a_11630_4086# x5.X.t24 VDD.t634 VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X816 a_3912_2366# x4.X.t68 VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X817 a_6977_3239# a_6465_3213# VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X818 a_6846_4086# x5.X.t25 VSS.t597 VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X819 a_11389_3239# x39.Q_N VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X820 VDD.t478 a_8858_4775# a_8768_5167# VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X821 a_7363_4801# VDD.t758 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X822 a_8939_4086# a_9237_4386# a_9173_4478# VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X823 a_7363_4801# a_6760_4775# a_7247_4775# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X824 a_6547_4086# a_6846_4086# a_6781_4112# VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X825 a_9464_3239# a_8402_3239# a_9369_3239# VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X826 VDD.t44 a_4854_3213# a_5561_3239# VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X827 a_4214_4801# VDD.t759 VSS.t142 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X828 x4.X.t0 a_1511_4112# VDD.t353 VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X829 a_4658_4086# a_4926_4296# a_4872_4394# VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.113 ps=1.11 w=0.84 l=0.15
X830 a_8697_4112# x4.X.t69 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.154 ps=1.34 w=0.64 l=0.15
X831 VSS.t605 x7.X a_2979_2366# VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X832 VDD.t244 a_2265_2340# a_2198_2732# VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.174 ps=1.41 w=0.84 l=0.15
X833 a_1508_5167# a_1227_4801# a_1415_4801# VDD.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X834 a_6410_2366# a_6546_2340# a_5991_2340# VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0864 ps=0.91 w=0.64 l=0.15
X835 VSS.t9 a_10681_4086# check[2].t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X836 a_7317_2550# a_6844_2640# a_7561_2366# VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0671 ps=0.75 w=0.36 l=0.15
X837 a_3504_2340# a_3599_2340# VSS.t42 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X838 a_11183_3239# a_10794_3239# a_11075_3605# VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X839 a_7246_3213# x45.Q_N VDD.t249 VDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
R0 D[3].n8 D[3].t2 269.921
R1 D[3].n8 D[3].t3 234.573
R2 D[3].n7 D[3].t1 207.373
R3 D[3].n9 D[3].n8 76.0005
R4 D[3].n14 D[3].t0 34.8148
R5 D[3].n11 D[3] 26.5622
R6 D[3].n12 D[3].n11 19.8539
R7 D[3].n11 D[3].n10 14.6672
R8 D[3] D[3].n7 9.01934
R9 D[3] D[3].n14 8.8299
R10 D[3].n9 D[3] 7.57233
R11 D[3].n7 D[3] 7.45876
R12 D[3].n13 D[3].n12 3.14374
R13 D[3].n12 D[3].n6 2.74043
R14 D[3].n10 D[3].n9 2.70473
R15 D[3].n3 D[3] 2.62982
R16 D[3].n5 D[3].n1 2.26284
R17 D[3].n4 D[3].n3 2.23869
R18 D[3].n10 D[3] 1.9836
R19 D[3].n14 D[3].n13 0.412636
R20 D[3].n6 D[3].n0 0.0232273
R21 D[3].n4 D[3].n2 0.00807576
R22 D[3].n5 D[3].n4 0.00195195
R23 D[3].n6 D[3].n5 0.00194159
R24 VDD.n2145 VDD.t197 1574.59
R25 VDD.n1475 VDD.t486 500.865
R26 VDD.n1513 VDD.t92 500.865
R27 VDD.n1556 VDD.t204 500.865
R28 VDD.n1594 VDD.t557 500.865
R29 VDD.n1637 VDD.t206 500.865
R30 VDD.n914 VDD.t640 500.865
R31 VDD.n1210 VDD.t622 500.865
R32 VDD.n990 VDD.t311 500.865
R33 VDD.n1052 VDD.t595 500.865
R34 VDD.n220 VDD.t278 500.865
R35 VDD.n185 VDD.t438 500.865
R36 VDD.n150 VDD.t116 500.865
R37 VDD.n115 VDD.t240 500.865
R38 VDD.n2261 VDD.t536 500.865
R39 VDD.n2395 VDD.t422 500.865
R40 VDD.n2519 VDD.t547 500.865
R41 VDD.n2643 VDD.t134 500.865
R42 VDD.n2699 VDD.t472 500.865
R43 VDD.n1472 VDD.n1471 440.25
R44 VDD.n1511 VDD.n1510 440.25
R45 VDD.n1553 VDD.n1552 440.25
R46 VDD.n1592 VDD.n1591 440.25
R47 VDD.n1634 VDD.n1633 440.25
R48 VDD.n1285 VDD.n1284 440.25
R49 VDD.n953 VDD.n952 440.25
R50 VDD.n1127 VDD.n1126 440.25
R51 VDD.n1029 VDD.n1028 440.25
R52 VDD.n218 VDD.n217 440.25
R53 VDD.n183 VDD.n182 440.25
R54 VDD.n148 VDD.n147 440.25
R55 VDD.n113 VDD.n112 440.25
R56 VDD.n2273 VDD.n2272 440.25
R57 VDD.n2405 VDD.n2404 440.25
R58 VDD.n2529 VDD.n2528 440.25
R59 VDD.n2653 VDD.n2652 440.25
R60 VDD.n2690 VDD.n2689 440.25
R61 VDD.n288 VDD.t169 397.163
R62 VDD.n377 VDD.t175 397.163
R63 VDD.n466 VDD.t154 397.163
R64 VDD.n555 VDD.t139 397.163
R65 VDD.t172 VDD.n2756 397.144
R66 VDD.t160 VDD.n2592 397.144
R67 VDD.t142 VDD.n2468 397.144
R68 VDD.t178 VDD.n2344 397.144
R69 VDD.n2747 VDD.t157 394.462
R70 VDD.n2583 VDD.t151 394.462
R71 VDD.n2459 VDD.t187 394.462
R72 VDD.n2335 VDD.t181 394.462
R73 VDD.t145 VDD.n296 385.733
R74 VDD.t166 VDD.n385 385.733
R75 VDD.t163 VDD.n474 385.733
R76 VDD.t148 VDD.n563 385.733
R77 VDD.n1673 VDD.t658 374.342
R78 VDD.n1752 VDD.t648 374.342
R79 VDD.n1826 VDD.t650 374.342
R80 VDD.n1905 VDD.t644 374.342
R81 VDD.n1979 VDD.t654 374.342
R82 VDD.n1100 VDD.t646 374.342
R83 VDD.n1179 VDD.t656 374.342
R84 VDD.n1258 VDD.t652 374.342
R85 VDD.n520 VDD.t428 374.342
R86 VDD.n431 VDD.t466 374.342
R87 VDD.n342 VDD.t114 374.342
R88 VDD.n253 VDD.t74 374.342
R89 VDD.n2192 VDD.t138 374.342
R90 VDD.n2315 VDD.t614 374.342
R91 VDD.n2439 VDD.t70 374.342
R92 VDD.n2563 VDD.t674 374.342
R93 VDD.n2781 VDD.t722 374.342
R94 VDD.n1423 VDD.t581 373.63
R95 VDD.n2077 VDD.t539 354.697
R96 VDD.n2259 VDD.t185 326.317
R97 VDD.n2098 VDD.n2092 324.707
R98 VDD.n2098 VDD.n2091 324.707
R99 VDD.n2103 VDD.n2091 324.707
R100 VDD.n2103 VDD.n2085 324.707
R101 VDD.n2109 VDD.n2085 324.707
R102 VDD.n2109 VDD.n2084 324.707
R103 VDD.n2114 VDD.n2084 324.707
R104 VDD.n2114 VDD.n2080 324.707
R105 VDD.n2120 VDD.n2080 324.707
R106 VDD.n2120 VDD.n2079 324.707
R107 VDD.n2125 VDD.n2079 324.707
R108 VDD.n2125 VDD.n2073 324.707
R109 VDD.n2131 VDD.n2073 324.707
R110 VDD.n2131 VDD.n2072 324.707
R111 VDD.n2136 VDD.n2072 324.707
R112 VDD.n2136 VDD.n2065 324.707
R113 VDD.n2142 VDD.n2065 324.707
R114 VDD.n2142 VDD.n2064 324.707
R115 VDD.n2146 VDD.n2064 324.707
R116 VDD.n2156 VDD.n2058 324.707
R117 VDD.n2161 VDD.n2058 324.707
R118 VDD.n2161 VDD.n2054 324.707
R119 VDD.n2167 VDD.n2054 324.707
R120 VDD.n2167 VDD.n2053 324.707
R121 VDD.n2171 VDD.n2053 324.707
R122 VDD.n1666 VDD.n1664 324.707
R123 VDD.n1664 VDD.n1661 324.707
R124 VDD.n1675 VDD.n1661 324.707
R125 VDD.n1675 VDD.n1659 324.707
R126 VDD.n1680 VDD.n1659 324.707
R127 VDD.n1680 VDD.n1655 324.707
R128 VDD.n1689 VDD.n1655 324.707
R129 VDD.n1689 VDD.n1654 324.707
R130 VDD.n1693 VDD.n1654 324.707
R131 VDD.n1693 VDD.n1649 324.707
R132 VDD.n1699 VDD.n1649 324.707
R133 VDD.n1699 VDD.n1647 324.707
R134 VDD.n1702 VDD.n1647 324.707
R135 VDD.n1702 VDD.n1643 324.707
R136 VDD.n1711 VDD.n1643 324.707
R137 VDD.n1711 VDD.n1641 324.707
R138 VDD.n1716 VDD.n1641 324.707
R139 VDD.n1716 VDD.n1636 324.707
R140 VDD.n1722 VDD.n1636 324.707
R141 VDD.n1722 VDD.n1635 324.707
R142 VDD.n1726 VDD.n1635 324.707
R143 VDD.n1726 VDD.n1630 324.707
R144 VDD.n1732 VDD.n1630 324.707
R145 VDD.n1732 VDD.n1628 324.707
R146 VDD.n1737 VDD.n1628 324.707
R147 VDD.n1737 VDD.n1622 324.707
R148 VDD.n1745 VDD.n1622 324.707
R149 VDD.n1745 VDD.n1621 324.707
R150 VDD.n1750 VDD.n1621 324.707
R151 VDD.n1750 VDD.n1617 324.707
R152 VDD.n1757 VDD.n1617 324.707
R153 VDD.n1757 VDD.n1616 324.707
R154 VDD.n1761 VDD.n1616 324.707
R155 VDD.n1761 VDD.n1610 324.707
R156 VDD.n1768 VDD.n1610 324.707
R157 VDD.n1768 VDD.n1608 324.707
R158 VDD.n1772 VDD.n1608 324.707
R159 VDD.n1772 VDD.n1603 324.707
R160 VDD.n1778 VDD.n1603 324.707
R161 VDD.n1778 VDD.n1601 324.707
R162 VDD.n1782 VDD.n1601 324.707
R163 VDD.n1782 VDD.n1596 324.707
R164 VDD.n1791 VDD.n1596 324.707
R165 VDD.n1791 VDD.n1595 324.707
R166 VDD.n1796 VDD.n1595 324.707
R167 VDD.n1796 VDD.n1590 324.707
R168 VDD.n1802 VDD.n1590 324.707
R169 VDD.n1802 VDD.n1589 324.707
R170 VDD.n1807 VDD.n1589 324.707
R171 VDD.n1807 VDD.n1585 324.707
R172 VDD.n1816 VDD.n1585 324.707
R173 VDD.n1816 VDD.n1584 324.707
R174 VDD.n1820 VDD.n1584 324.707
R175 VDD.n1820 VDD.n1580 324.707
R176 VDD.n1828 VDD.n1580 324.707
R177 VDD.n1828 VDD.n1578 324.707
R178 VDD.n1833 VDD.n1578 324.707
R179 VDD.n1833 VDD.n1574 324.707
R180 VDD.n1842 VDD.n1574 324.707
R181 VDD.n1842 VDD.n1573 324.707
R182 VDD.n1846 VDD.n1573 324.707
R183 VDD.n1846 VDD.n1568 324.707
R184 VDD.n1852 VDD.n1568 324.707
R185 VDD.n1852 VDD.n1566 324.707
R186 VDD.n1855 VDD.n1566 324.707
R187 VDD.n1855 VDD.n1562 324.707
R188 VDD.n1864 VDD.n1562 324.707
R189 VDD.n1864 VDD.n1560 324.707
R190 VDD.n1869 VDD.n1560 324.707
R191 VDD.n1869 VDD.n1555 324.707
R192 VDD.n1875 VDD.n1555 324.707
R193 VDD.n1875 VDD.n1554 324.707
R194 VDD.n1879 VDD.n1554 324.707
R195 VDD.n1879 VDD.n1549 324.707
R196 VDD.n1885 VDD.n1549 324.707
R197 VDD.n1885 VDD.n1547 324.707
R198 VDD.n1890 VDD.n1547 324.707
R199 VDD.n1890 VDD.n1541 324.707
R200 VDD.n1898 VDD.n1541 324.707
R201 VDD.n1898 VDD.n1540 324.707
R202 VDD.n1903 VDD.n1540 324.707
R203 VDD.n1903 VDD.n1536 324.707
R204 VDD.n1910 VDD.n1536 324.707
R205 VDD.n1910 VDD.n1535 324.707
R206 VDD.n1914 VDD.n1535 324.707
R207 VDD.n1914 VDD.n1529 324.707
R208 VDD.n1921 VDD.n1529 324.707
R209 VDD.n1921 VDD.n1527 324.707
R210 VDD.n1925 VDD.n1527 324.707
R211 VDD.n1925 VDD.n1522 324.707
R212 VDD.n1931 VDD.n1522 324.707
R213 VDD.n1931 VDD.n1520 324.707
R214 VDD.n1935 VDD.n1520 324.707
R215 VDD.n1935 VDD.n1515 324.707
R216 VDD.n1944 VDD.n1515 324.707
R217 VDD.n1944 VDD.n1514 324.707
R218 VDD.n1949 VDD.n1514 324.707
R219 VDD.n1949 VDD.n1509 324.707
R220 VDD.n1955 VDD.n1509 324.707
R221 VDD.n1955 VDD.n1508 324.707
R222 VDD.n1960 VDD.n1508 324.707
R223 VDD.n1960 VDD.n1504 324.707
R224 VDD.n1969 VDD.n1504 324.707
R225 VDD.n1969 VDD.n1503 324.707
R226 VDD.n1973 VDD.n1503 324.707
R227 VDD.n1973 VDD.n1499 324.707
R228 VDD.n1981 VDD.n1499 324.707
R229 VDD.n1981 VDD.n1497 324.707
R230 VDD.n1986 VDD.n1497 324.707
R231 VDD.n1986 VDD.n1493 324.707
R232 VDD.n1995 VDD.n1493 324.707
R233 VDD.n1995 VDD.n1492 324.707
R234 VDD.n1999 VDD.n1492 324.707
R235 VDD.n1999 VDD.n1487 324.707
R236 VDD.n2005 VDD.n1487 324.707
R237 VDD.n2005 VDD.n1485 324.707
R238 VDD.n2008 VDD.n1485 324.707
R239 VDD.n2008 VDD.n1481 324.707
R240 VDD.n2017 VDD.n1481 324.707
R241 VDD.n2017 VDD.n1479 324.707
R242 VDD.n2022 VDD.n1479 324.707
R243 VDD.n2022 VDD.n1474 324.707
R244 VDD.n2028 VDD.n1474 324.707
R245 VDD.n2028 VDD.n1473 324.707
R246 VDD.n2032 VDD.n1473 324.707
R247 VDD.n2032 VDD.n1468 324.707
R248 VDD.n2038 VDD.n1468 324.707
R249 VDD.n2038 VDD.n1466 324.707
R250 VDD.n2041 VDD.n1466 324.707
R251 VDD.n1036 VDD.n1034 324.707
R252 VDD.n1040 VDD.n1034 324.707
R253 VDD.n1040 VDD.n1026 324.707
R254 VDD.n1046 VDD.n1026 324.707
R255 VDD.n1046 VDD.n1025 324.707
R256 VDD.n1051 VDD.n1025 324.707
R257 VDD.n1051 VDD.n1021 324.707
R258 VDD.n1058 VDD.n1021 324.707
R259 VDD.n1058 VDD.n1020 324.707
R260 VDD.n1063 VDD.n1020 324.707
R261 VDD.n1063 VDD.n1014 324.707
R262 VDD.n1069 VDD.n1014 324.707
R263 VDD.n1069 VDD.n1013 324.707
R264 VDD.n1073 VDD.n1013 324.707
R265 VDD.n1073 VDD.n1009 324.707
R266 VDD.n1081 VDD.n1009 324.707
R267 VDD.n1081 VDD.n1008 324.707
R268 VDD.n1086 VDD.n1008 324.707
R269 VDD.n1086 VDD.n1003 324.707
R270 VDD.n1093 VDD.n1003 324.707
R271 VDD.n1093 VDD.n1002 324.707
R272 VDD.n1098 VDD.n1002 324.707
R273 VDD.n1098 VDD.n998 324.707
R274 VDD.n1108 VDD.n998 324.707
R275 VDD.n1108 VDD.n997 324.707
R276 VDD.n1113 VDD.n997 324.707
R277 VDD.n1113 VDD.n994 324.707
R278 VDD.n1121 VDD.n994 324.707
R279 VDD.n1121 VDD.n993 324.707
R280 VDD.n1125 VDD.n993 324.707
R281 VDD.n1125 VDD.n988 324.707
R282 VDD.n1133 VDD.n988 324.707
R283 VDD.n1133 VDD.n986 324.707
R284 VDD.n1138 VDD.n986 324.707
R285 VDD.n1138 VDD.n982 324.707
R286 VDD.n1146 VDD.n982 324.707
R287 VDD.n1146 VDD.n981 324.707
R288 VDD.n1150 VDD.n981 324.707
R289 VDD.n1150 VDD.n975 324.707
R290 VDD.n1156 VDD.n975 324.707
R291 VDD.n1156 VDD.n974 324.707
R292 VDD.n1161 VDD.n974 324.707
R293 VDD.n1161 VDD.n970 324.707
R294 VDD.n1169 VDD.n970 324.707
R295 VDD.n1169 VDD.n969 324.707
R296 VDD.n1174 VDD.n969 324.707
R297 VDD.n1174 VDD.n965 324.707
R298 VDD.n1181 VDD.n965 324.707
R299 VDD.n1181 VDD.n964 324.707
R300 VDD.n1186 VDD.n964 324.707
R301 VDD.n1186 VDD.n959 324.707
R302 VDD.n1193 VDD.n959 324.707
R303 VDD.n1193 VDD.n958 324.707
R304 VDD.n1198 VDD.n958 324.707
R305 VDD.n1198 VDD.n950 324.707
R306 VDD.n1204 VDD.n950 324.707
R307 VDD.n1204 VDD.n949 324.707
R308 VDD.n1209 VDD.n949 324.707
R309 VDD.n1209 VDD.n945 324.707
R310 VDD.n1216 VDD.n945 324.707
R311 VDD.n1216 VDD.n944 324.707
R312 VDD.n1221 VDD.n944 324.707
R313 VDD.n1221 VDD.n938 324.707
R314 VDD.n1227 VDD.n938 324.707
R315 VDD.n1227 VDD.n937 324.707
R316 VDD.n1231 VDD.n937 324.707
R317 VDD.n1231 VDD.n933 324.707
R318 VDD.n1239 VDD.n933 324.707
R319 VDD.n1239 VDD.n932 324.707
R320 VDD.n1244 VDD.n932 324.707
R321 VDD.n1244 VDD.n927 324.707
R322 VDD.n1251 VDD.n927 324.707
R323 VDD.n1251 VDD.n926 324.707
R324 VDD.n1256 VDD.n926 324.707
R325 VDD.n1256 VDD.n922 324.707
R326 VDD.n1266 VDD.n922 324.707
R327 VDD.n1266 VDD.n921 324.707
R328 VDD.n1271 VDD.n921 324.707
R329 VDD.n1271 VDD.n918 324.707
R330 VDD.n1279 VDD.n918 324.707
R331 VDD.n1279 VDD.n917 324.707
R332 VDD.n1283 VDD.n917 324.707
R333 VDD.n1283 VDD.n912 324.707
R334 VDD.n1291 VDD.n912 324.707
R335 VDD.n1291 VDD.n909 324.707
R336 VDD.n1300 VDD.n909 324.707
R337 VDD.n1454 VDD.n825 324.707
R338 VDD.n1458 VDD.n825 324.707
R339 VDD.n579 VDD.n116 324.707
R340 VDD.n579 VDD.n111 324.707
R341 VDD.n586 VDD.n111 324.707
R342 VDD.n586 VDD.n110 324.707
R343 VDD.n591 VDD.n110 324.707
R344 VDD.n591 VDD.n108 324.707
R345 VDD.n108 VDD.n103 324.707
R346 VDD.n599 VDD.n103 324.707
R347 VDD.n599 VDD.n101 324.707
R348 VDD.n604 VDD.n101 324.707
R349 VDD.n604 VDD.n95 324.707
R350 VDD.n612 VDD.n95 324.707
R351 VDD.n612 VDD.n93 324.707
R352 VDD.n618 VDD.n93 324.707
R353 VDD.n618 VDD.n94 324.707
R354 VDD.n94 VDD.n88 324.707
R355 VDD.n628 VDD.n88 324.707
R356 VDD.n628 VDD.n86 324.707
R357 VDD.n738 VDD.n22 324.707
R358 VDD.n747 VDD.n22 324.707
R359 VDD.n747 VDD.n21 324.707
R360 VDD.n752 VDD.n21 324.707
R361 VDD.n752 VDD.n17 324.707
R362 VDD.n758 VDD.n17 324.707
R363 VDD.n758 VDD.n16 324.707
R364 VDD.n762 VDD.n16 324.707
R365 VDD.n490 VDD.n151 324.707
R366 VDD.n490 VDD.n146 324.707
R367 VDD.n496 VDD.n146 324.707
R368 VDD.n496 VDD.n145 324.707
R369 VDD.n501 VDD.n145 324.707
R370 VDD.n501 VDD.n141 324.707
R371 VDD.n510 VDD.n141 324.707
R372 VDD.n510 VDD.n140 324.707
R373 VDD.n514 VDD.n140 324.707
R374 VDD.n514 VDD.n136 324.707
R375 VDD.n522 VDD.n136 324.707
R376 VDD.n522 VDD.n134 324.707
R377 VDD.n527 VDD.n134 324.707
R378 VDD.n527 VDD.n130 324.707
R379 VDD.n536 VDD.n130 324.707
R380 VDD.n536 VDD.n129 324.707
R381 VDD.n540 VDD.n129 324.707
R382 VDD.n540 VDD.n124 324.707
R383 VDD.n546 VDD.n124 324.707
R384 VDD.n546 VDD.n122 324.707
R385 VDD.n549 VDD.n122 324.707
R386 VDD.n549 VDD.n118 324.707
R387 VDD.n574 VDD.n118 324.707
R388 VDD.n401 VDD.n186 324.707
R389 VDD.n401 VDD.n181 324.707
R390 VDD.n407 VDD.n181 324.707
R391 VDD.n407 VDD.n180 324.707
R392 VDD.n412 VDD.n180 324.707
R393 VDD.n412 VDD.n176 324.707
R394 VDD.n421 VDD.n176 324.707
R395 VDD.n421 VDD.n175 324.707
R396 VDD.n425 VDD.n175 324.707
R397 VDD.n425 VDD.n171 324.707
R398 VDD.n433 VDD.n171 324.707
R399 VDD.n433 VDD.n169 324.707
R400 VDD.n438 VDD.n169 324.707
R401 VDD.n438 VDD.n165 324.707
R402 VDD.n447 VDD.n165 324.707
R403 VDD.n447 VDD.n164 324.707
R404 VDD.n451 VDD.n164 324.707
R405 VDD.n451 VDD.n159 324.707
R406 VDD.n457 VDD.n159 324.707
R407 VDD.n457 VDD.n157 324.707
R408 VDD.n460 VDD.n157 324.707
R409 VDD.n460 VDD.n153 324.707
R410 VDD.n485 VDD.n153 324.707
R411 VDD.n312 VDD.n221 324.707
R412 VDD.n312 VDD.n216 324.707
R413 VDD.n318 VDD.n216 324.707
R414 VDD.n318 VDD.n215 324.707
R415 VDD.n323 VDD.n215 324.707
R416 VDD.n323 VDD.n211 324.707
R417 VDD.n332 VDD.n211 324.707
R418 VDD.n332 VDD.n210 324.707
R419 VDD.n336 VDD.n210 324.707
R420 VDD.n336 VDD.n206 324.707
R421 VDD.n344 VDD.n206 324.707
R422 VDD.n344 VDD.n204 324.707
R423 VDD.n349 VDD.n204 324.707
R424 VDD.n349 VDD.n200 324.707
R425 VDD.n358 VDD.n200 324.707
R426 VDD.n358 VDD.n199 324.707
R427 VDD.n362 VDD.n199 324.707
R428 VDD.n362 VDD.n194 324.707
R429 VDD.n368 VDD.n194 324.707
R430 VDD.n368 VDD.n192 324.707
R431 VDD.n371 VDD.n192 324.707
R432 VDD.n371 VDD.n188 324.707
R433 VDD.n396 VDD.n188 324.707
R434 VDD.n246 VDD.n244 324.707
R435 VDD.n244 VDD.n241 324.707
R436 VDD.n255 VDD.n241 324.707
R437 VDD.n255 VDD.n239 324.707
R438 VDD.n260 VDD.n239 324.707
R439 VDD.n260 VDD.n235 324.707
R440 VDD.n269 VDD.n235 324.707
R441 VDD.n269 VDD.n234 324.707
R442 VDD.n273 VDD.n234 324.707
R443 VDD.n273 VDD.n229 324.707
R444 VDD.n279 VDD.n229 324.707
R445 VDD.n279 VDD.n227 324.707
R446 VDD.n282 VDD.n227 324.707
R447 VDD.n282 VDD.n223 324.707
R448 VDD.n307 VDD.n223 324.707
R449 VDD.n801 VDD.n779 318.858
R450 VDD.n2088 VDD.n2087 315.596
R451 VDD.n786 VDD.n779 315.43
R452 VDD.n801 VDD.n778 315.43
R453 VDD.n806 VDD.n772 315.43
R454 VDD.n816 VDD.n772 315.43
R455 VDD.n816 VDD.n771 315.43
R456 VDD.n820 VDD.n771 315.43
R457 VDD.n1743 VDD.n1742 312.132
R458 VDD.n1822 VDD.n1582 312.132
R459 VDD.n1896 VDD.n1895 312.132
R460 VDD.n1975 VDD.n1501 312.132
R461 VDD.n1669 VDD.n1663 312.132
R462 VDD.n1106 VDD.n1105 312.132
R463 VDD.n1188 VDD.n962 312.132
R464 VDD.n1264 VDD.n1263 312.132
R465 VDD.n516 VDD.n138 312.132
R466 VDD.n427 VDD.n173 312.132
R467 VDD.n338 VDD.n208 312.132
R468 VDD.n249 VDD.n243 312.132
R469 VDD.n2183 VDD.n2176 312.132
R470 VDD.n2298 VDD.n9 312.132
R471 VDD.n2430 VDD.n5 312.132
R472 VDD.n2554 VDD.n1 312.132
R473 VDD.n2790 VDD.n2789 312.132
R474 VDD.n806 VDD.n778 312
R475 VDD.n1438 VDD.n1436 311.387
R476 VDD.n2096 VDD.n2095 307.478
R477 VDD.n1687 VDD.n1686 307.212
R478 VDD.n1763 VDD.n1614 307.212
R479 VDD.n1840 VDD.n1839 307.212
R480 VDD.n1916 VDD.n1533 307.212
R481 VDD.n1993 VDD.n1992 307.212
R482 VDD.n1088 VDD.n1006 307.212
R483 VDD.n1167 VDD.n1166 307.212
R484 VDD.n1246 VDD.n930 307.212
R485 VDD.n534 VDD.n533 307.212
R486 VDD.n445 VDD.n444 307.212
R487 VDD.n356 VDD.n355 307.212
R488 VDD.n267 VDD.n266 307.212
R489 VDD.n2210 VDD.n2206 307.212
R490 VDD.n2331 VDD.n2330 306.985
R491 VDD.n2455 VDD.n2454 306.985
R492 VDD.n2579 VDD.n2578 306.985
R493 VDD.n2764 VDD.n2763 306.985
R494 VDD.n1385 VDD.n1383 306.546
R495 VDD.n1707 VDD.n1706 305.529
R496 VDD.n1786 VDD.n1785 305.529
R497 VDD.n1860 VDD.n1859 305.529
R498 VDD.n1939 VDD.n1938 305.529
R499 VDD.n2013 VDD.n2012 305.529
R500 VDD.n1018 VDD.n1017 305.529
R501 VDD.n1142 VDD.n1141 305.529
R502 VDD.n942 VDD.n941 305.529
R503 VDD.n2249 VDD.n2245 305.529
R504 VDD.n2383 VDD.n2379 305.529
R505 VDD.n2507 VDD.n2503 305.529
R506 VDD.n2631 VDD.n2627 305.529
R507 VDD.n2714 VDD.n2710 305.529
R508 VDD.n571 VDD.n565 305.3
R509 VDD.n482 VDD.n476 305.3
R510 VDD.n393 VDD.n387 305.3
R511 VDD.n304 VDD.n298 305.3
R512 VDD.n1305 VDD.n1304 304.861
R513 VDD.n2266 VDD.t184 289.93
R514 VDD.n1454 VDD.n826 289.413
R515 VDD.n738 VDD.n27 289.413
R516 VDD.n786 VDD.t715 287.635
R517 VDD.t146 VDD.t461 281.096
R518 VDD.t167 VDD.t16 281.096
R519 VDD.t164 VDD.t431 281.096
R520 VDD.t149 VDD.t552 281.096
R521 VDD.n2741 VDD.t173 276.317
R522 VDD.n2598 VDD.t161 276.317
R523 VDD.n2474 VDD.t143 276.317
R524 VDD.n2350 VDD.t179 276.317
R525 VDD.n1294 VDD.n902 264.707
R526 VDD.n1315 VDD.n900 264.707
R527 VDD.n1322 VDD.n892 264.707
R528 VDD.n1335 VDD.n888 264.707
R529 VDD.n1339 VDD.n881 264.707
R530 VDD.n1354 VDD.n879 264.707
R531 VDD.n1364 VDD.n874 264.707
R532 VDD.n1368 VDD.n867 264.707
R533 VDD.n1382 VDD.n865 264.707
R534 VDD.n1388 VDD.n860 264.707
R535 VDD.n1401 VDD.n856 264.707
R536 VDD.n1405 VDD.n849 264.707
R537 VDD.n1422 VDD.n846 264.707
R538 VDD.n1418 VDD.n839 264.707
R539 VDD.n1435 VDD.n837 264.707
R540 VDD.n1441 VDD.n831 264.707
R541 VDD.n646 VDD.n74 264.707
R542 VDD.n658 VDD.n72 264.707
R543 VDD.n666 VDD.n63 264.707
R544 VDD.n680 VDD.n58 264.707
R545 VDD.n684 VDD.n52 264.707
R546 VDD.n696 VDD.n50 264.707
R547 VDD.n704 VDD.n41 264.707
R548 VDD.n718 VDD.n36 264.707
R549 VDD.n722 VDD.n29 264.707
R550 VDD.t257 VDD.t146 249.863
R551 VDD.t57 VDD.t167 249.863
R552 VDD.t662 VDD.t164 249.863
R553 VDD.t675 VDD.t149 249.863
R554 VDD.n1676 VDD.n1660 242.779
R555 VDD.n1692 VDD.n1691 242.779
R556 VDD.n1700 VDD.n1648 242.779
R557 VDD.t304 VDD.n1701 242.779
R558 VDD.n1712 VDD.n1642 242.779
R559 VDD.n1724 VDD.n1723 242.779
R560 VDD.n1733 VDD.n1629 242.779
R561 VDD.n1736 VDD.n1735 242.779
R562 VDD.n1749 VDD.n1747 242.779
R563 VDD.n1769 VDD.n1609 242.779
R564 VDD.n1771 VDD.n1770 242.779
R565 VDD.t525 VDD.n1602 242.779
R566 VDD.n1781 VDD.n1779 242.779
R567 VDD.n1795 VDD.n1794 242.779
R568 VDD.n1806 VDD.n1804 242.779
R569 VDD.n1818 VDD.n1817 242.779
R570 VDD.n1829 VDD.n1579 242.779
R571 VDD.n1845 VDD.n1844 242.779
R572 VDD.n1853 VDD.n1567 242.779
R573 VDD.t322 VDD.n1854 242.779
R574 VDD.n1865 VDD.n1561 242.779
R575 VDD.n1877 VDD.n1876 242.779
R576 VDD.n1886 VDD.n1548 242.779
R577 VDD.n1889 VDD.n1888 242.779
R578 VDD.n1902 VDD.n1900 242.779
R579 VDD.n1922 VDD.n1528 242.779
R580 VDD.n1924 VDD.n1923 242.779
R581 VDD.t220 VDD.n1521 242.779
R582 VDD.n1934 VDD.n1932 242.779
R583 VDD.n1948 VDD.n1947 242.779
R584 VDD.n1959 VDD.n1957 242.779
R585 VDD.n1971 VDD.n1970 242.779
R586 VDD.n1982 VDD.n1498 242.779
R587 VDD.n1998 VDD.n1997 242.779
R588 VDD.n2006 VDD.n1486 242.779
R589 VDD.t530 VDD.n2007 242.779
R590 VDD.n2018 VDD.n1480 242.779
R591 VDD.n2030 VDD.n2029 242.779
R592 VDD.n2039 VDD.n1467 242.779
R593 VDD.n2113 VDD.n2111 241.436
R594 VDD.n2122 VDD.n2121 241.436
R595 VDD.n2124 VDD.n2123 241.436
R596 VDD.n256 VDD.n240 239.452
R597 VDD.n272 VDD.n271 239.452
R598 VDD.n280 VDD.n228 239.452
R599 VDD.t0 VDD.n281 239.452
R600 VDD.n308 VDD.n222 239.452
R601 VDD.n311 VDD.n310 239.452
R602 VDD.n322 VDD.n320 239.452
R603 VDD.n334 VDD.n333 239.452
R604 VDD.n345 VDD.n205 239.452
R605 VDD.n361 VDD.n360 239.452
R606 VDD.n369 VDD.n193 239.452
R607 VDD.t347 VDD.n370 239.452
R608 VDD.n397 VDD.n187 239.452
R609 VDD.n400 VDD.n399 239.452
R610 VDD.n411 VDD.n409 239.452
R611 VDD.n423 VDD.n422 239.452
R612 VDD.n434 VDD.n170 239.452
R613 VDD.n450 VDD.n449 239.452
R614 VDD.n458 VDD.n158 239.452
R615 VDD.t679 VDD.n459 239.452
R616 VDD.n486 VDD.n152 239.452
R617 VDD.n489 VDD.n488 239.452
R618 VDD.n500 VDD.n498 239.452
R619 VDD.n512 VDD.n511 239.452
R620 VDD.n523 VDD.n135 239.452
R621 VDD.n539 VDD.n538 239.452
R622 VDD.n547 VDD.n123 239.452
R623 VDD.t64 VDD.n548 239.452
R624 VDD.n575 VDD.n117 239.452
R625 VDD.n578 VDD.n577 239.452
R626 VDD.n590 VDD.n588 239.452
R627 VDD.n600 VDD.n102 239.452
R628 VDD.n601 VDD.n600 239.452
R629 VDD.n1039 VDD.n1038 237.5
R630 VDD.n1050 VDD.n1048 237.5
R631 VDD.n1062 VDD.n1061 237.5
R632 VDD.n1070 VDD.t253 237.5
R633 VDD.n1072 VDD.n1071 237.5
R634 VDD.n1083 VDD.n1082 237.5
R635 VDD.n1097 VDD.n1096 237.5
R636 VDD.n1123 VDD.n1122 237.5
R637 VDD.n1134 VDD.n987 237.5
R638 VDD.n1148 VDD.n1147 237.5
R639 VDD.t54 VDD.n1149 237.5
R640 VDD.n1158 VDD.n1157 237.5
R641 VDD.n1160 VDD.n1159 237.5
R642 VDD.n1183 VDD.n1182 237.5
R643 VDD.n1197 VDD.n1196 237.5
R644 VDD.n1208 VDD.n1206 237.5
R645 VDD.n1220 VDD.n1219 237.5
R646 VDD.n1228 VDD.t611 237.5
R647 VDD.n1230 VDD.n1229 237.5
R648 VDD.n1241 VDD.n1240 237.5
R649 VDD.n1255 VDD.n1254 237.5
R650 VDD.n1281 VDD.n1280 237.5
R651 VDD.n1292 VDD.n911 237.5
R652 VDD.n1456 VDD.n1455 237.5
R653 VDD.n1300 VDD.n910 232.941
R654 VDD.n2101 VDD.t308 230.94
R655 VDD.n1457 VDD.t62 229.756
R656 VDD.n634 VDD.n86 229.412
R657 VDD.n642 VDD.n81 229.412
R658 VDD.n297 VDD.t145 229.072
R659 VDD.n386 VDD.t166 229.072
R660 VDD.n475 VDD.t163 229.072
R661 VDD.n564 VDD.t148 229.072
R662 VDD.t190 VDD.t207 221.667
R663 VDD.t304 VDD.t72 221.667
R664 VDD.t558 VDD.t739 221.667
R665 VDD.t331 VDD.t525 221.667
R666 VDD.t314 VDD.t201 221.667
R667 VDD.t322 VDD.t87 221.667
R668 VDD.t89 VDD.t484 221.667
R669 VDD.t199 VDD.t220 221.667
R670 VDD.t332 VDD.t487 221.667
R671 VDD.t530 VDD.t216 221.667
R672 VDD.n2113 VDD.t247 220.442
R673 VDD.t197 VDD.t193 220.442
R674 VDD.t524 VDD.t279 218.631
R675 VDD.t0 VDD.t502 218.631
R676 VDD.t30 VDD.t439 218.631
R677 VDD.t347 VDD.t209 218.631
R678 VDD.t97 VDD.t117 218.631
R679 VDD.t679 VDD.t481 218.631
R680 VDD.t283 VDD.t237 218.631
R681 VDD.t64 VDD.t436 218.631
R682 VDD.t374 VDD.t380 218.631
R683 VDD.t253 VDD.t520 216.849
R684 VDD.t592 VDD.t68 216.849
R685 VDD.t54 VDD.t700 216.849
R686 VDD.t11 VDD.t312 216.849
R687 VDD.t611 VDD.t272 216.849
R688 VDD.t619 VDD.t666 216.849
R689 VDD.t4 VDD.n2110 209.946
R690 VDD.t538 VDD.n2122 209.946
R691 VDD.t731 VDD.n1690 208.472
R692 VDD.n1760 VDD.t617 208.472
R693 VDD.t629 VDD.n1843 208.472
R694 VDD.n1913 VDD.t384 208.472
R695 VDD.t105 VDD.n1996 208.472
R696 VDD.n613 VDD.t358 208.22
R697 VDD.t356 VDD.n614 208.22
R698 VDD.n2265 VDD.t750 208.013
R699 VDD.t170 VDD.n270 205.617
R700 VDD.t176 VDD.n359 205.617
R701 VDD.t155 VDD.n448 205.617
R702 VDD.t140 VDD.n537 205.617
R703 VDD.n1085 VDD.t83 203.94
R704 VDD.n1170 VDD.t516 203.94
R705 VDD.n1243 VDD.t250 203.94
R706 VDD.n105 VDD.t361 201.19
R707 VDD.n2796 VDD 200
R708 VDD.n2 VDD 200
R709 VDD.n6 VDD 200
R710 VDD.n10 VDD 200
R711 VDD.n2112 VDD.t501 199.448
R712 VDD.n2168 VDD 199.448
R713 VDD.n737 VDD.t596 197.809
R714 VDD.n759 VDD 197.809
R715 VDD.n1112 VDD 196.196
R716 VDD.n1194 VDD 196.196
R717 VDD.n1270 VDD 196.196
R718 VDD.n1713 VDD.t493 195.279
R719 VDD.n1723 VDD.t205 195.279
R720 VDD.t725 VDD.n1780 195.279
R721 VDD.n1795 VDD.t556 195.279
R722 VDD.n1866 VDD.t229 195.279
R723 VDD.n1876 VDD.t203 195.279
R724 VDD.t35 VDD.n1933 195.279
R725 VDD.n1948 VDD.t91 195.279
R726 VDD.n2019 VDD.t590 195.279
R727 VDD.n2029 VDD.t485 195.279
R728 VDD.n695 VDD.n694 195.206
R729 VDD.n817 VDD 195.136
R730 VDD.n1295 VDD.n901 193.614
R731 VDD.n1314 VDD.n1313 193.614
R732 VDD.n1353 VDD.n1350 193.614
R733 VDD.n1419 VDD.n838 193.614
R734 VDD.n311 VDD.t277 192.603
R735 VDD.n400 VDD.t437 192.603
R736 VDD.n489 VDD.t115 192.603
R737 VDD.n578 VDD.t239 192.603
R738 VDD.n1050 VDD.t594 191.034
R739 VDD.t264 VDD.n1060 191.034
R740 VDD.t310 VDD.n1134 191.034
R741 VDD.n1136 VDD.t20 191.034
R742 VDD.n1208 VDD.t621 191.034
R743 VDD.t131 VDD.n1218 191.034
R744 VDD.t639 VDD.n1292 191.034
R745 VDD.t574 VDD.n51 190
R746 VDD.t372 VDD.n602 187.398
R747 VDD.n617 VDD.t366 187.398
R748 VDD.n831 VDD.n830 185
R749 VDD.n1443 VDD.n831 185
R750 VDD.n1439 VDD.n1435 185
R751 VDD.n1435 VDD.n1434 185
R752 VDD.n840 VDD.n839 185
R753 VDD.n839 VDD.n838 185
R754 VDD.n1424 VDD.n1422 185
R755 VDD.n1422 VDD.n1421 185
R756 VDD.n850 VDD.n849 185
R757 VDD.n849 VDD.n848 185
R758 VDD.n1401 VDD.n1400 185
R759 VDD.n1402 VDD.n1401 185
R760 VDD.n860 VDD.n859 185
R761 VDD.n1390 VDD.n860 185
R762 VDD.n1386 VDD.n1382 185
R763 VDD.n1382 VDD.n1381 185
R764 VDD.n868 VDD.n867 185
R765 VDD.n867 VDD.n866 185
R766 VDD.n1364 VDD.n1363 185
R767 VDD.n1365 VDD.n1364 185
R768 VDD.n1354 VDD.n1353 185
R769 VDD.n882 VDD.n881 185
R770 VDD.n881 VDD.n880 185
R771 VDD.n1335 VDD.n1334 185
R772 VDD.n1336 VDD.n1335 185
R773 VDD.n892 VDD.n891 185
R774 VDD.n1324 VDD.n892 185
R775 VDD.n1316 VDD.n1315 185
R776 VDD.n1315 VDD.n1314 185
R777 VDD.n903 VDD.n902 185
R778 VDD.n902 VDD.n901 185
R779 VDD.n910 VDD.n905 185
R780 VDD.n1298 VDD.n910 185
R781 VDD.n30 VDD.n29 185
R782 VDD.n29 VDD.n28 185
R783 VDD.n718 VDD.n717 185
R784 VDD.n719 VDD.n718 185
R785 VDD.n41 VDD.n40 185
R786 VDD.n706 VDD.n41 185
R787 VDD.n697 VDD.n696 185
R788 VDD.n696 VDD.n695 185
R789 VDD.n53 VDD.n52 185
R790 VDD.n52 VDD.n51 185
R791 VDD.n680 VDD.n679 185
R792 VDD.n681 VDD.n680 185
R793 VDD.n63 VDD.n62 185
R794 VDD.n668 VDD.n63 185
R795 VDD.n659 VDD.n658 185
R796 VDD.n658 VDD.n657 185
R797 VDD.n75 VDD.n74 185
R798 VDD.n74 VDD.n73 185
R799 VDD.n642 VDD.n641 185
R800 VDD.n643 VDD.n642 185
R801 VDD.n635 VDD.n634 185
R802 VDD.n634 VDD.n633 185
R803 VDD.t566 VDD.n705 182.192
R804 VDD.n2133 VDD.t537 181.077
R805 VDD.t184 VDD.n2265 179.094
R806 VDD.t624 VDD.n866 178.125
R807 VDD.n736 VDD.t602 176.987
R808 VDD.n785 VDD.t711 174.595
R809 VDD.n2071 VDD.n2070 174.595
R810 VDD.n716 VDD.n37 174.595
R811 VDD.n698 VDD.n49 174.595
R812 VDD.n678 VDD.n59 174.595
R813 VDD.n660 VDD.n71 174.595
R814 VDD.n78 VDD.n77 174.595
R815 VDD.n85 VDD.n84 174.595
R816 VDD.n626 VDD.n89 174.595
R817 VDD.n620 VDD.n619 174.595
R818 VDD.n98 VDD.n97 174.595
R819 VDD.n606 VDD.n605 174.595
R820 VDD.n1678 VDD.t475 171.529
R821 VDD.t28 VDD.n1759 171.529
R822 VDD.n1831 VDD.t95 171.529
R823 VDD.t119 VDD.n1912 171.529
R824 VDD.n1984 VDD.t245 171.529
R825 VDD.n2766 VDD.t542 171.054
R826 VDD.n2573 VDD.t477 171.054
R827 VDD.n2449 VDD.t328 171.054
R828 VDD.n2325 VDD.t582 171.054
R829 VDD.n1336 VDD.t401 170.381
R830 VDD.n1626 VDD.n1625 169.184
R831 VDD.n1811 VDD.n1810 169.184
R832 VDD.n1545 VDD.n1544 169.184
R833 VDD.n1964 VDD.n1963 169.184
R834 VDD.n1464 VDD.n1463 169.184
R835 VDD.n1117 VDD.n1116 169.184
R836 VDD.n956 VDD.n955 169.184
R837 VDD.n1275 VDD.n1274 169.184
R838 VDD.n1032 VDD.n1031 169.184
R839 VDD.n594 VDD.n107 169.184
R840 VDD.n505 VDD.n504 169.184
R841 VDD.n416 VDD.n415 169.184
R842 VDD.n327 VDD.n326 169.184
R843 VDD.n2288 VDD.n2284 169.184
R844 VDD.n2420 VDD.n2416 169.184
R845 VDD.n2544 VDD.n2540 169.184
R846 VDD.n2668 VDD.n2664 169.184
R847 VDD.n2677 VDD.n2673 169.184
R848 VDD.n258 VDD.t390 169.179
R849 VDD.n347 VDD.t273 169.179
R850 VDD.n436 VDD.t703 169.179
R851 VDD.n525 VDD.t510 169.179
R852 VDD.n681 VDD.t354 169.179
R853 VDD.t341 VDD.n1084 167.799
R854 VDD.n1171 VDD.t445 167.799
R855 VDD.t499 VDD.n1242 167.799
R856 VDD.n603 VDD.t360 166.576
R857 VDD.n616 VDD.t352 166.576
R858 VDD.n1651 VDD.n1650 166.542
R859 VDD.n1607 VDD.n1606 166.542
R860 VDD.n1570 VDD.n1569 166.542
R861 VDD.n1526 VDD.n1525 166.542
R862 VDD.n1489 VDD.n1488 166.542
R863 VDD.n1075 VDD.n1074 166.542
R864 VDD.n978 VDD.n977 166.542
R865 VDD.n1233 VDD.n1232 166.542
R866 VDD.n1357 VDD.n1356 166.542
R867 VDD.n126 VDD.n125 166.542
R868 VDD.n161 VDD.n160 166.542
R869 VDD.n196 VDD.n195 166.542
R870 VDD.n231 VDD.n230 166.542
R871 VDD.n2221 VDD.n2220 166.542
R872 VDD.n2355 VDD.n2354 166.542
R873 VDD.n2479 VDD.n2478 166.542
R874 VDD.n2603 VDD.n2602 166.542
R875 VDD.n2736 VDD.n2735 166.542
R876 VDD.n2057 VDD.n2056 166.381
R877 VDD.n777 VDD.n776 166.381
R878 VDD.n20 VDD.n19 166.381
R879 VDD.n2051 VDD.n2050 166.006
R880 VDD.n14 VDD.n13 166.006
R881 VDD.n2143 VDD.t413 165.332
R882 VDD.n2145 VDD.t415 165.332
R883 VDD.n1391 VDD.t400 165.218
R884 VDD.n2061 VDD.n2060 164.453
R885 VDD.n25 VDD.n24 164.453
R886 VDD.n2147 VDD.t416 163.582
R887 VDD.n770 VDD.n769 162.47
R888 VDD.n707 VDD.t570 161.37
R889 VDD.n799 VDD.n781 160.918
R890 VDD.n2132 VDD.t698 160.083
R891 VDD.n31 VDD.t577 159.46
R892 VDD.n1725 VDD.t564 158.333
R893 VDD.n1803 VDD.t51 158.333
R894 VDD.n1878 VDD.t441 158.333
R895 VDD.n1956 VDD.t423 158.333
R896 VDD.n2031 VDD.t425 158.333
R897 VDD.n1338 VDD.t77 157.474
R898 VDD.n1365 VDD.t637 157.474
R899 VDD.t398 VDD.n1433 157.474
R900 VDD.n2135 VDD.t79 157.459
R901 VDD.t195 VDD.n2157 157.459
R902 VDD.n319 VDD.t288 156.165
R903 VDD.n408 VDD.t109 156.165
R904 VDD.n497 VDD.t294 156.165
R905 VDD.n587 VDD.t40 156.165
R906 VDD.t598 VDD.n748 156.165
R907 VDD.t49 VDD.n1047 154.892
R908 VDD.n1124 VDD.t296 154.892
R909 VDD.t455 VDD.n1205 154.892
R910 VDD.n1282 VDD.t449 154.892
R911 VDD.n1715 VDD.t733 153.056
R912 VDD.n1792 VDD.t615 153.056
R913 VDD.n1868 VDD.t627 153.056
R914 VDD.n1945 VDD.t386 153.056
R915 VDD.n2021 VDD.t107 153.056
R916 VDD.n824 VDD.t63 152.88
R917 VDD.n2757 VDD.t172 152.694
R918 VDD.n295 VDD.n294 152
R919 VDD.n384 VDD.n383 152
R920 VDD.n473 VDD.n472 152
R921 VDD.n562 VDD.n561 152
R922 VDD.n2593 VDD.t160 151.811
R923 VDD.n2469 VDD.t142 151.811
R924 VDD.t713 VDD.n802 151.487
R925 VDD.t81 VDD.n1059 149.728
R926 VDD.n1137 VDD.t514 149.728
R927 VDD.t248 VDD.n1217 149.728
R928 VDD.n1299 VDD.t669 149.728
R929 VDD.n1324 VDD.t350 149.728
R930 VDD.n2345 VDD.t178 149.322
R931 VDD.n668 VDD.t364 148.357
R932 VDD.n739 VDD.t597 148.195
R933 VDD.t580 VDD.n1417 147.148
R934 VDD.n1455 VDD 147.148
R935 VDD.t697 VDD.n2101 146.962
R936 VDD.n2149 VDD.t198 145.868
R937 VDD.n615 VDD.t362 145.754
R938 VDD.n737 VDD 145.754
R939 VDD.t305 VDD.n1678 145.139
R940 VDD.t495 VDD.n1629 145.139
R941 VDD.n1759 VDD.t526 145.139
R942 VDD.n1804 VDD.t727 145.139
R943 VDD.t325 VDD.n1831 145.139
R944 VDD.t231 VDD.n1548 145.139
R945 VDD.n1912 VDD.t217 145.139
R946 VDD.n1957 VDD.t31 145.139
R947 VDD.t529 VDD.n1984 145.139
R948 VDD.t588 VDD.n1467 145.139
R949 VDD.n2276 VDD.t223 144.738
R950 VDD.n1404 VDD.t349 144.565
R951 VDD.t417 VDD.n2134 144.338
R952 VDD.n2144 VDD.t411 144.338
R953 VDD.t1 VDD.n258 143.151
R954 VDD.n320 VDD.t459 143.151
R955 VDD.t348 VDD.n347 143.151
R956 VDD.n409 VDD.t14 143.151
R957 VDD.t680 VDD.n436 143.151
R958 VDD.n498 VDD.t429 143.151
R959 VDD.t65 VDD.n525 143.151
R960 VDD.n588 VDD.t550 143.151
R961 VDD.n784 VDD.t716 142.571
R962 VDD.t483 VDD.n1714 142.5
R963 VDD.n1793 VDD.t406 142.5
R964 VDD.t397 VDD.n1867 142.5
R965 VDD.n1946 VDD.t8 142.5
R966 VDD.t612 VDD.n2020 142.5
R967 VDD.n1038 VDD.t266 141.984
R968 VDD.n1084 VDD.t252 141.984
R969 VDD.t24 VDD.n1123 141.984
R970 VDD.t53 VDD.n1171 141.984
R971 VDD.n1196 VDD.t129 141.984
R972 VDD.n1242 VDD.t610 141.984
R973 VDD.t45 VDD.n1281 141.984
R974 VDD.n309 VDD.t257 140.548
R975 VDD.n398 VDD.t57 140.548
R976 VDD.n487 VDD.t662 140.548
R977 VDD.n576 VDD.t675 140.548
R978 VDD.n721 VDD.t576 140.548
R979 VDD.n1049 VDD.t270 139.403
R980 VDD.t321 VDD.n1135 139.403
R981 VDD.n1207 VDD.t659 139.403
R982 VDD.t740 VDD.n1293 139.403
R983 VDD.t306 VDD.n1660 137.222
R984 VDD.n1701 VDD.t473 137.222
R985 VDD.n1747 VDD.t527 137.222
R986 VDD.t26 VDD.n1602 137.222
R987 VDD.t323 VDD.n1579 137.222
R988 VDD.n1854 VDD.t93 137.222
R989 VDD.n1900 VDD.t218 137.222
R990 VDD.t121 VDD.n1521 137.222
R991 VDD.t531 VDD.n1498 137.222
R992 VDD.n2007 VDD.t243 137.222
R993 VDD.n1381 VDD.t667 136.821
R994 VDD.t578 VDD.n1442 136.821
R995 VDD.n2100 VDD.t518 136.464
R996 VDD.t191 VDD.n2158 136.464
R997 VDD.t2 VDD.n240 135.343
R998 VDD.n281 VDD.t388 135.343
R999 VDD.t345 VDD.n205 135.343
R1000 VDD.n370 VDD.t275 135.343
R1001 VDD.t681 VDD.n170 135.343
R1002 VDD.n459 VDD.t701 135.343
R1003 VDD.t66 VDD.n135 135.343
R1004 VDD.n548 VDD.t512 135.343
R1005 VDD.t600 VDD.n749 135.343
R1006 VDD.n2041 VDD.t677 135.118
R1007 VDD.n2756 VDD.t748 134.986
R1008 VDD.n2592 VDD.t747 134.986
R1009 VDD.n2468 VDD.t755 134.986
R1010 VDD.n2344 VDD.t759 134.986
R1011 VDD.n288 VDD.t757 134.966
R1012 VDD.n377 VDD.t745 134.966
R1013 VDD.n466 VDD.t751 134.966
R1014 VDD.n555 VDD.t756 134.966
R1015 VDD.n1734 VDD.t491 134.583
R1016 VDD.t729 VDD.n1805 134.583
R1017 VDD.n1887 VDD.t233 134.583
R1018 VDD.t33 VDD.n1958 134.583
R1019 VDD.n2040 VDD.t586 134.583
R1020 VDD.n2747 VDD.t749 134.484
R1021 VDD.n2583 VDD.t754 134.484
R1022 VDD.n2459 VDD.t758 134.484
R1023 VDD.n2335 VDD.t743 134.484
R1024 VDD.t343 VDD.n1070 134.239
R1025 VDD.n1096 VDD.t254 134.239
R1026 VDD.n1149 VDD.t447 134.239
R1027 VDD.t55 VDD.n1183 134.239
R1028 VDD.t497 VDD.n1228 134.239
R1029 VDD.n1254 VDD.t608 134.239
R1030 VDD.n295 VDD.t753 133.5
R1031 VDD.n384 VDD.t744 133.5
R1032 VDD.n473 VDD.t746 133.5
R1033 VDD.n562 VDD.t752 133.5
R1034 VDD.t463 VDD.n321 132.74
R1035 VDD.t18 VDD.n410 132.74
R1036 VDD.t433 VDD.n499 132.74
R1037 VDD.t554 VDD.n589 132.74
R1038 VDD.t641 VDD.n1036 132.363
R1039 VDD.t268 VDD.n1037 131.659
R1040 VDD.n1111 VDD.t22 131.659
R1041 VDD.t127 VDD.n1195 131.659
R1042 VDD.n1269 VDD.t43 131.659
R1043 VDD.t709 VDD.n803 130.946
R1044 VDD.n657 VDD.t376 127.534
R1045 VDD.n1677 VDD.t657 126.668
R1046 VDD.n1736 VDD.t60 126.668
R1047 VDD.t647 VDD.n1748 126.668
R1048 VDD.n1817 VDD.t221 126.668
R1049 VDD.n1830 VDD.t649 126.668
R1050 VDD.n1889 VDD.t339 126.668
R1051 VDD.t643 VDD.n1901 126.668
R1052 VDD.n1970 VDD.t741 126.668
R1053 VDD.n1983 VDD.t653 126.668
R1054 VDD.n2102 VDD.t623 125.968
R1055 VDD.t560 VDD.n2159 125.968
R1056 VDD.t562 VDD.n2168 125.968
R1057 VDD.n2170 VDD.t281 125.968
R1058 VDD.n257 VDD.t73 124.933
R1059 VDD.n333 VDD.t6 124.933
R1060 VDD.n346 VDD.t113 124.933
R1061 VDD.n422 VDD.t85 124.933
R1062 VDD.n435 VDD.t465 124.933
R1063 VDD.n511 VDD.t38 124.933
R1064 VDD.n524 VDD.t427 124.933
R1065 VDD.t125 VDD.n102 124.933
R1066 VDD.t382 VDD.n629 124.933
R1067 VDD.t660 VDD.n750 124.933
R1068 VDD.t211 VDD.n759 124.933
R1069 VDD.n761 VDD.t235 124.933
R1070 VDD.n1679 VDD.t71 124.028
R1071 VDD.n1758 VDD.t330 124.028
R1072 VDD.n1832 VDD.t88 124.028
R1073 VDD.n1911 VDD.t200 124.028
R1074 VDD.n1985 VDD.t215 124.028
R1075 VDD.t645 VDD.n1095 123.913
R1076 VDD.n1112 VDD.t664 123.913
R1077 VDD.n1172 VDD.t655 123.913
R1078 VDD.t467 VDD.n1194 123.913
R1079 VDD.t651 VDD.n1253 123.913
R1080 VDD.n1270 VDD.t58 123.913
R1081 VDD VDD.t689 123.684
R1082 VDD.t625 VDD 123.684
R1083 VDD.t683 VDD 123.684
R1084 VDD.t685 VDD 123.684
R1085 VDD.t693 VDD 123.684
R1086 VDD.t453 VDD.n804 123.243
R1087 VDD.t606 VDD.n817 123.243
R1088 VDD.n819 VDD.t604 123.243
R1089 VDD.n259 VDD.t503 122.329
R1090 VDD.n348 VDD.t210 122.329
R1091 VDD.n437 VDD.t482 122.329
R1092 VDD.n526 VDD.t435 122.329
R1093 VDD.n2068 VDD.n2067 121.769
R1094 VDD.t521 VDD.n1094 121.332
R1095 VDD VDD.t522 121.332
R1096 VDD.n1173 VDD.t699 121.332
R1097 VDD.t548 VDD 121.332
R1098 VDD.t271 VDD.n1252 121.332
R1099 VDD VDD.t9 121.332
R1100 VDD.t71 VDD.n1677 118.751
R1101 VDD.n1748 VDD.t330 118.751
R1102 VDD.t88 VDD.n1830 118.751
R1103 VDD.n1901 VDD.t200 118.751
R1104 VDD.t215 VDD.n1983 118.751
R1105 VDD.n2774 VDD.t124 118.421
R1106 VDD.n2565 VDD.t489 118.421
R1107 VDD.n2441 VDD.t407 118.421
R1108 VDD.n2317 VDD.t504 118.421
R1109 VDD.n2194 VDD.t723 118.421
R1110 VDD.t503 VDD.n257 117.124
R1111 VDD.t210 VDD.n346 117.124
R1112 VDD.t482 VDD.n435 117.124
R1113 VDD.t435 VDD.n524 117.124
R1114 VDD.n1095 VDD.t521 116.168
R1115 VDD.t699 VDD.n1172 116.168
R1116 VDD.n1253 VDD.t271 116.168
R1117 VDD.t290 VDD.n1665 116.112
R1118 VDD.t657 VDD.n1676 116.112
R1119 VDD.t60 VDD.n1734 116.112
R1120 VDD.n1746 VDD.t213 116.112
R1121 VDD.n1749 VDD.t647 116.112
R1122 VDD.n1805 VDD.t221 116.112
R1123 VDD.n1819 VDD.t402 116.112
R1124 VDD.t649 VDD.n1829 116.112
R1125 VDD.t339 VDD.n1887 116.112
R1126 VDD.n1899 VDD.t409 116.112
R1127 VDD.n1902 VDD.t643 116.112
R1128 VDD.n1958 VDD.t741 116.112
R1129 VDD.n1972 VDD.t631 116.112
R1130 VDD.t653 VDD.n1982 116.112
R1131 VDD.t677 VDD.n2040 116.112
R1132 VDD.n2674 VDD.t457 115.79
R1133 VDD.n2778 VDD.t721 115.79
R1134 VDD.t689 VDD.n2793 115.79
R1135 VDD.n2665 VDD.t241 115.79
R1136 VDD.n2560 VDD.t673 115.79
R1137 VDD.n2551 VDD.t625 115.79
R1138 VDD.n2541 VDD.t451 115.79
R1139 VDD.n2436 VDD.t69 115.79
R1140 VDD.n2427 VDD.t683 115.79
R1141 VDD.n2417 VDD.t719 115.79
R1142 VDD.n2312 VDD.t613 115.79
R1143 VDD.n2295 VDD.t685 115.79
R1144 VDD.n2285 VDD.t717 115.79
R1145 VDD.n2189 VDD.t137 115.79
R1146 VDD.n2180 VDD.t693 115.79
R1147 VDD.n2099 VDD.t404 115.471
R1148 VDD.t623 VDD.n2100 115.471
R1149 VDD.n2160 VDD.t560 115.471
R1150 VDD.n2169 VDD.t562 115.471
R1151 VDD.t281 VDD.n2169 115.471
R1152 VDD.t633 VDD.n245 114.522
R1153 VDD.t73 VDD.n256 114.522
R1154 VDD.n321 VDD.t6 114.522
R1155 VDD.n335 VDD.t695 114.522
R1156 VDD.t113 VDD.n345 114.522
R1157 VDD.n410 VDD.t85 114.522
R1158 VDD.n424 VDD.t691 114.522
R1159 VDD.t465 VDD.n434 114.522
R1160 VDD.n499 VDD.t38 114.522
R1161 VDD.n513 VDD.t687 114.522
R1162 VDD.t427 VDD.n523 114.522
R1163 VDD.n589 VDD.t125 114.522
R1164 VDD.n630 VDD.t382 114.522
R1165 VDD.n751 VDD.t660 114.522
R1166 VDD.n760 VDD.t211 114.522
R1167 VDD.t235 VDD.n760 114.522
R1168 VDD.n1037 VDD.t641 113.588
R1169 VDD.n1097 VDD.t645 113.588
R1170 VDD.t522 VDD.n1109 113.588
R1171 VDD.t664 VDD.n1111 113.588
R1172 VDD.n1182 VDD.t655 113.588
R1173 VDD.n1185 VDD.t548 113.588
R1174 VDD.n1195 VDD.t467 113.588
R1175 VDD.n1255 VDD.t651 113.588
R1176 VDD.t9 VDD.n1267 113.588
R1177 VDD.t58 VDD.n1269 113.588
R1178 VDD.n805 VDD.t453 112.974
R1179 VDD.n818 VDD.t606 112.974
R1180 VDD.t604 VDD.n818 112.974
R1181 VDD.t491 VDD.n1733 108.195
R1182 VDD.n1806 VDD.t729 108.195
R1183 VDD.t233 VDD.n1886 108.195
R1184 VDD.n1959 VDD.t33 108.195
R1185 VDD.t586 VDD.n2039 108.195
R1186 VDD.n2679 VDD.t262 107.895
R1187 VDD.n2660 VDD.t337 107.895
R1188 VDD.n2536 VDD.t317 107.895
R1189 VDD.n2412 VDD.t99 107.895
R1190 VDD.n2280 VDD.t227 107.895
R1191 VDD.n322 VDD.t463 106.713
R1192 VDD.n411 VDD.t18 106.713
R1193 VDD.n500 VDD.t433 106.713
R1194 VDD.n590 VDD.t554 106.713
R1195 VDD.t368 VDD.n73 106.713
R1196 VDD.n1039 VDD.t268 105.843
R1197 VDD.n1122 VDD.t22 105.843
R1198 VDD.n1197 VDD.t127 105.843
R1199 VDD.n1280 VDD.t43 105.843
R1200 VDD.n1665 VDD.t306 105.556
R1201 VDD.t473 VDD.n1700 105.556
R1202 VDD.t527 VDD.n1746 105.556
R1203 VDD.n1771 VDD.t26 105.556
R1204 VDD.n1819 VDD.t323 105.556
R1205 VDD.t93 VDD.n1853 105.556
R1206 VDD.t218 VDD.n1899 105.556
R1207 VDD.n1924 VDD.t121 105.556
R1208 VDD.n1972 VDD.t531 105.556
R1209 VDD.t243 VDD.n2006 105.556
R1210 VDD.n2731 VDD.t540 105.263
R1211 VDD.n2793 VDD.t285 105.263
R1212 VDD.n2608 VDD.t479 105.263
R1213 VDD.n2551 VDD.t707 105.263
R1214 VDD.n2484 VDD.t326 105.263
R1215 VDD.n2427 VDD.t735 105.263
R1216 VDD.n2360 VDD.t584 105.263
R1217 VDD.n2295 VDD.t300 105.263
R1218 VDD.n2226 VDD.t394 105.263
R1219 VDD.n2180 VDD.t506 105.263
R1220 VDD.t518 VDD.n2099 104.972
R1221 VDD.n2160 VDD.t191 104.972
R1222 VDD.n245 VDD.t2 104.111
R1223 VDD.t388 VDD.n280 104.111
R1224 VDD.n335 VDD.t345 104.111
R1225 VDD.t275 VDD.n369 104.111
R1226 VDD.n424 VDD.t681 104.111
R1227 VDD.t701 VDD.n458 104.111
R1228 VDD.n513 VDD.t66 104.111
R1229 VDD.t512 VDD.n547 104.111
R1230 VDD.t370 VDD.n630 104.111
R1231 VDD.n751 VDD.t600 104.111
R1232 VDD.n1072 VDD.t343 103.261
R1233 VDD.n1109 VDD.t254 103.261
R1234 VDD.n1157 VDD.t447 103.261
R1235 VDD.n1185 VDD.t55 103.261
R1236 VDD.n1230 VDD.t497 103.261
R1237 VDD.n1267 VDD.t608 103.261
R1238 VDD.n805 VDD.t709 102.704
R1239 VDD.n1390 VDD.t75 100.68
R1240 VDD.n1715 VDD.t483 100.278
R1241 VDD.t406 VDD.n1792 100.278
R1242 VDD.n1868 VDD.t397 100.278
R1243 VDD.t8 VDD.n1945 100.278
R1244 VDD.n2021 VDD.t612 100.278
R1245 VDD.n2706 VDD.t42 100.001
R1246 VDD.n2633 VDD.t636 100.001
R1247 VDD.n2509 VDD.t635 100.001
R1248 VDD.n2385 VDD.t256 100.001
R1249 VDD.n2251 VDD.t663 100.001
R1250 VDD.n1059 VDD.t270 98.0983
R1251 VDD.n1137 VDD.t321 98.0983
R1252 VDD.n1217 VDD.t659 98.0983
R1253 VDD.n1299 VDD.t740 98.0983
R1254 VDD.n1679 VDD.t305 97.6394
R1255 VDD.n1725 VDD.t495 97.6394
R1256 VDD.t526 VDD.n1758 97.6394
R1257 VDD.t727 VDD.n1803 97.6394
R1258 VDD.n1832 VDD.t325 97.6394
R1259 VDD.n1878 VDD.t231 97.6394
R1260 VDD.t217 VDD.n1911 97.6394
R1261 VDD.t31 VDD.n1956 97.6394
R1262 VDD.n1985 VDD.t529 97.6394
R1263 VDD.n2031 VDD.t588 97.6394
R1264 VDD.n2687 VDD.t260 97.3689
R1265 VDD.n2770 VDD.t284 97.3689
R1266 VDD.n2650 VDD.t333 97.3689
R1267 VDD.n2569 VDD.t705 97.3689
R1268 VDD.n2526 VDD.t315 97.3689
R1269 VDD.n2445 VDD.t737 97.3689
R1270 VDD.n2402 VDD.t101 97.3689
R1271 VDD.n2321 VDD.t302 97.3689
R1272 VDD.n2198 VDD.t508 97.3689
R1273 VDD.n2135 VDD.t417 97.0999
R1274 VDD.t411 VDD.n2143 97.0999
R1275 VDD.n259 VDD.t1 96.3019
R1276 VDD.t459 VDD.n319 96.3019
R1277 VDD.n348 VDD.t348 96.3019
R1278 VDD.t14 VDD.n408 96.3019
R1279 VDD.n437 VDD.t680 96.3019
R1280 VDD.t429 VDD.n497 96.3019
R1281 VDD.n526 VDD.t65 96.3019
R1282 VDD.t550 VDD.n587 96.3019
R1283 VDD.n1047 VDD.t266 95.5168
R1284 VDD.n1094 VDD.t252 95.5168
R1285 VDD.n1124 VDD.t24 95.5168
R1286 VDD.n1173 VDD.t53 95.5168
R1287 VDD.n1205 VDD.t129 95.5168
R1288 VDD.n1252 VDD.t610 95.5168
R1289 VDD.n1282 VDD.t45 95.5168
R1290 VDD.n2102 VDD.t697 94.4756
R1291 VDD.n629 VDD.t362 93.6991
R1292 VDD.t75 VDD.n1389 92.9353
R1293 VDD.n787 VDD.n786 92.5005
R1294 VDD.n771 VDD.n770 92.5005
R1295 VDD.n818 VDD.n771 92.5005
R1296 VDD.n816 VDD.n815 92.5005
R1297 VDD.n817 VDD.n816 92.5005
R1298 VDD.n808 VDD.n772 92.5005
R1299 VDD.n804 VDD.n772 92.5005
R1300 VDD.n807 VDD.n806 92.5005
R1301 VDD.n806 VDD.n805 92.5005
R1302 VDD.n782 VDD.n778 92.5005
R1303 VDD.n803 VDD.n778 92.5005
R1304 VDD.n801 VDD.n800 92.5005
R1305 VDD.n802 VDD.n801 92.5005
R1306 VDD.n821 VDD.n820 92.5005
R1307 VDD.n820 VDD.n819 92.5005
R1308 VDD.n791 VDD.n779 92.5005
R1309 VDD.n785 VDD.n779 92.5005
R1310 VDD.n1446 VDD.n1445 92.5005
R1311 VDD.n833 VDD.n832 92.5005
R1312 VDD.n1432 VDD.n1431 92.5005
R1313 VDD.n1420 VDD.n847 92.5005
R1314 VDD.n1416 VDD.n1415 92.5005
R1315 VDD.n1403 VDD.n855 92.5005
R1316 VDD.n1393 VDD.n1392 92.5005
R1317 VDD.n862 VDD.n861 92.5005
R1318 VDD.n1379 VDD.n1378 92.5005
R1319 VDD.n1366 VDD.n873 92.5005
R1320 VDD.n1352 VDD.n878 92.5005
R1321 VDD.n1349 VDD.n1348 92.5005
R1322 VDD.n1337 VDD.n887 92.5005
R1323 VDD.n1327 VDD.n1326 92.5005
R1324 VDD.n894 VDD.n893 92.5005
R1325 VDD.n1312 VDD.n1311 92.5005
R1326 VDD.n1297 VDD.n1296 92.5005
R1327 VDD.n1447 VDD.n1446 92.5005
R1328 VDD.n1431 VDD.n1430 92.5005
R1329 VDD.n1415 VDD.n1414 92.5005
R1330 VDD.n855 VDD.n853 92.5005
R1331 VDD.n1394 VDD.n1393 92.5005
R1332 VDD.n1378 VDD.n1377 92.5005
R1333 VDD.n873 VDD.n871 92.5005
R1334 VDD.n1348 VDD.n1347 92.5005
R1335 VDD.n887 VDD.n885 92.5005
R1336 VDD.n1328 VDD.n1327 92.5005
R1337 VDD.n895 VDD.n894 92.5005
R1338 VDD.n1311 VDD.n1310 92.5005
R1339 VDD.n734 VDD.n733 92.5005
R1340 VDD.n720 VDD.n35 92.5005
R1341 VDD.n709 VDD.n708 92.5005
R1342 VDD.n43 VDD.n42 92.5005
R1343 VDD.n693 VDD.n692 92.5005
R1344 VDD.n682 VDD.n57 92.5005
R1345 VDD.n671 VDD.n670 92.5005
R1346 VDD.n65 VDD.n64 92.5005
R1347 VDD.n655 VDD.n654 92.5005
R1348 VDD.n644 VDD.n80 92.5005
R1349 VDD.n733 VDD.n732 92.5005
R1350 VDD.n35 VDD.n33 92.5005
R1351 VDD.n710 VDD.n709 92.5005
R1352 VDD.n44 VDD.n43 92.5005
R1353 VDD.n692 VDD.n691 92.5005
R1354 VDD.n57 VDD.n55 92.5005
R1355 VDD.n672 VDD.n671 92.5005
R1356 VDD.n66 VDD.n65 92.5005
R1357 VDD.n654 VDD.n653 92.5005
R1358 VDD.n640 VDD.n80 92.5005
R1359 VDD.n1686 VDD.t732 91.4648
R1360 VDD.n1706 VDD.t494 91.4648
R1361 VDD.n1706 VDD.t734 91.4648
R1362 VDD.n1614 VDD.t618 91.4648
R1363 VDD.n1785 VDD.t726 91.4648
R1364 VDD.n1785 VDD.t616 91.4648
R1365 VDD.n1839 VDD.t630 91.4648
R1366 VDD.n1859 VDD.t230 91.4648
R1367 VDD.n1859 VDD.t628 91.4648
R1368 VDD.n1533 VDD.t385 91.4648
R1369 VDD.n1938 VDD.t36 91.4648
R1370 VDD.n1938 VDD.t387 91.4648
R1371 VDD.n1992 VDD.t106 91.4648
R1372 VDD.n2012 VDD.t591 91.4648
R1373 VDD.n2012 VDD.t108 91.4648
R1374 VDD.n1017 VDD.t82 91.4648
R1375 VDD.n1017 VDD.t265 91.4648
R1376 VDD.n1006 VDD.t84 91.4648
R1377 VDD.n1141 VDD.t515 91.4648
R1378 VDD.n1141 VDD.t21 91.4648
R1379 VDD.n1166 VDD.t517 91.4648
R1380 VDD.n941 VDD.t249 91.4648
R1381 VDD.n941 VDD.t132 91.4648
R1382 VDD.n930 VDD.t251 91.4648
R1383 VDD.n1304 VDD.t670 91.4648
R1384 VDD.n1304 VDD.t48 91.4648
R1385 VDD.n1383 VDD.t668 91.4648
R1386 VDD.n565 VDD.t553 91.4648
R1387 VDD.n565 VDD.t150 91.4648
R1388 VDD.n533 VDD.t141 91.4648
R1389 VDD.n476 VDD.t432 91.4648
R1390 VDD.n476 VDD.t165 91.4648
R1391 VDD.n444 VDD.t156 91.4648
R1392 VDD.n387 VDD.t17 91.4648
R1393 VDD.n387 VDD.t168 91.4648
R1394 VDD.n355 VDD.t177 91.4648
R1395 VDD.n298 VDD.t462 91.4648
R1396 VDD.n298 VDD.t147 91.4648
R1397 VDD.n266 VDD.t171 91.4648
R1398 VDD.n2206 VDD.t444 91.4648
R1399 VDD.n2245 VDD.t672 91.4648
R1400 VDD.n2245 VDD.t226 91.4648
R1401 VDD.n2330 VDD.t180 91.4648
R1402 VDD.n2379 VDD.t183 91.4648
R1403 VDD.n2379 VDD.t104 91.4648
R1404 VDD.n2454 VDD.t144 91.4648
R1405 VDD.n2503 VDD.t189 91.4648
R1406 VDD.n2503 VDD.t320 91.4648
R1407 VDD.n2578 VDD.t162 91.4648
R1408 VDD.n2627 VDD.t153 91.4648
R1409 VDD.n2627 VDD.t336 91.4648
R1410 VDD.n2763 VDD.t174 91.4648
R1411 VDD.n2710 VDD.t159 91.4648
R1412 VDD.n2710 VDD.t259 91.4648
R1413 VDD.t733 VDD.n1713 89.7227
R1414 VDD.n1780 VDD.t615 89.7227
R1415 VDD.t627 VDD.n1866 89.7227
R1416 VDD.n1933 VDD.t386 89.7227
R1417 VDD.t107 VDD.n2019 89.7227
R1418 VDD.n2711 VDD.t158 89.4742
R1419 VDD.n2628 VDD.t152 89.4742
R1420 VDD.n2504 VDD.t188 89.4742
R1421 VDD.n2380 VDD.t182 89.4742
R1422 VDD.n2246 VDD.t671 89.4742
R1423 VDD.n645 VDD.t368 88.4936
R1424 VDD.n1060 VDD.t81 87.7722
R1425 VDD.t514 VDD.n1136 87.7722
R1426 VDD.n1218 VDD.t248 87.7722
R1427 VDD.n2265 VDD 87.6875
R1428 VDD.n1686 VDD.t476 86.7743
R1429 VDD.n1650 VDD.t474 86.7743
R1430 VDD.n1614 VDD.t29 86.7743
R1431 VDD.n1606 VDD.t27 86.7743
R1432 VDD.n1839 VDD.t96 86.7743
R1433 VDD.n1569 VDD.t94 86.7743
R1434 VDD.n1533 VDD.t120 86.7743
R1435 VDD.n1525 VDD.t122 86.7743
R1436 VDD.n1992 VDD.t246 86.7743
R1437 VDD.n1488 VDD.t244 86.7743
R1438 VDD.n1074 VDD.t344 86.7743
R1439 VDD.n1006 VDD.t342 86.7743
R1440 VDD.n977 VDD.t448 86.7743
R1441 VDD.n1166 VDD.t446 86.7743
R1442 VDD.n1232 VDD.t498 86.7743
R1443 VDD.n930 VDD.t500 86.7743
R1444 VDD.n1356 VDD.t78 86.7743
R1445 VDD.n1383 VDD.t76 86.7743
R1446 VDD.n533 VDD.t511 86.7743
R1447 VDD.n125 VDD.t513 86.7743
R1448 VDD.n444 VDD.t704 86.7743
R1449 VDD.n160 VDD.t702 86.7743
R1450 VDD.n355 VDD.t274 86.7743
R1451 VDD.n195 VDD.t276 86.7743
R1452 VDD.n266 VDD.t391 86.7743
R1453 VDD.n230 VDD.t389 86.7743
R1454 VDD.n2220 VDD.t395 86.7743
R1455 VDD.n2206 VDD.t393 86.7743
R1456 VDD.n2330 VDD.t583 86.7743
R1457 VDD.n2354 VDD.t585 86.7743
R1458 VDD.n2454 VDD.t329 86.7743
R1459 VDD.n2478 VDD.t327 86.7743
R1460 VDD.n2578 VDD.t478 86.7743
R1461 VDD.n2602 VDD.t480 86.7743
R1462 VDD.n2763 VDD.t543 86.7743
R1463 VDD.n2735 VDD.t541 86.7743
R1464 VDD.n643 VDD.t378 85.8909
R1465 VDD.n803 VDD.t713 84.7302
R1466 VDD.t564 VDD.n1724 84.4449
R1467 VDD.n1794 VDD.t51 84.4449
R1468 VDD.t441 VDD.n1877 84.4449
R1469 VDD.n1947 VDD.t423 84.4449
R1470 VDD.t425 VDD.n2030 84.4449
R1471 VDD.n2693 VDD.t292 84.211
R1472 VDD.n2646 VDD.t12 84.211
R1473 VDD.n2522 VDD.t298 84.211
R1474 VDD.n2398 VDD.t111 84.211
R1475 VDD.t79 VDD.n2133 83.9784
R1476 VDD.n2158 VDD.t195 83.9784
R1477 VDD.n310 VDD.t288 83.2882
R1478 VDD.n399 VDD.t109 83.2882
R1479 VDD.n488 VDD.t294 83.2882
R1480 VDD.n577 VDD.t40 83.2882
R1481 VDD.n631 VDD.t378 83.2882
R1482 VDD.n749 VDD.t598 83.2882
R1483 VDD.n1048 VDD.t49 82.6092
R1484 VDD.t296 VDD.n987 82.6092
R1485 VDD.n1206 VDD.t455 82.6092
R1486 VDD.t449 VDD.n911 82.6092
R1487 VDD.n2123 VDD.t698 81.3541
R1488 VDD VDD.t290 79.1672
R1489 VDD VDD.t213 79.1672
R1490 VDD.t402 VDD 79.1672
R1491 VDD VDD.t409 79.1672
R1492 VDD.t631 VDD 79.1672
R1493 VDD VDD.t404 78.7298
R1494 VDD VDD.t633 78.0827
R1495 VDD.t695 VDD 78.0827
R1496 VDD.t691 VDD 78.0827
R1497 VDD.t687 VDD 78.0827
R1498 VDD.n2134 VDD.t413 76.1055
R1499 VDD.t415 VDD.n2144 76.1055
R1500 VDD.n296 VDD.n287 75.2776
R1501 VDD.n385 VDD.n376 75.2776
R1502 VDD.n474 VDD.n465 75.2776
R1503 VDD.n563 VDD.n554 75.2776
R1504 VDD.t360 VDD.n601 72.8772
R1505 VDD.t352 VDD.n615 72.8772
R1506 VDD.n1690 VDD.t475 71.2505
R1507 VDD.n1760 VDD.t28 71.2505
R1508 VDD.n1843 VDD.t95 71.2505
R1509 VDD.n1913 VDD.t119 71.2505
R1510 VDD.n1996 VDD.t245 71.2505
R1511 VDD.n2207 VDD.t392 71.0531
R1512 VDD.n270 VDD.t390 70.2745
R1513 VDD.n359 VDD.t273 70.2745
R1514 VDD.n448 VDD.t703 70.2745
R1515 VDD.n537 VDD.t510 70.2745
R1516 VDD.n1085 VDD.t341 69.7016
R1517 VDD.t445 VDD.n1170 69.7016
R1518 VDD.n1243 VDD.t499 69.7016
R1519 VDD.t376 VDD.n656 67.6717
R1520 VDD VDD.n735 67.6717
R1521 VDD.n633 VDD.t370 65.069
R1522 VDD.n802 VDD.t711 64.1897
R1523 VDD.n1471 VDD.t426 63.1021
R1524 VDD.n1510 VDD.t424 63.1021
R1525 VDD.n1552 VDD.t442 63.1021
R1526 VDD.n1591 VDD.t52 63.1021
R1527 VDD.n1633 VDD.t565 63.1021
R1528 VDD.n1284 VDD.t450 63.1021
R1529 VDD.n952 VDD.t456 63.1021
R1530 VDD.n1126 VDD.t297 63.1021
R1531 VDD.n1028 VDD.t50 63.1021
R1532 VDD.n217 VDD.t289 63.1021
R1533 VDD.n182 VDD.t110 63.1021
R1534 VDD.n147 VDD.t295 63.1021
R1535 VDD.n112 VDD.t41 63.1021
R1536 VDD.n2272 VDD.t186 63.1021
R1537 VDD.n2404 VDD.t112 63.1021
R1538 VDD.n2528 VDD.t299 63.1021
R1539 VDD.n2652 VDD.t13 63.1021
R1540 VDD.n2689 VDD.t293 63.1021
R1541 VDD.n2157 VDD.t193 62.9839
R1542 VDD.n748 VDD.t602 62.4663
R1543 VDD.n2070 VDD.t80 61.563
R1544 VDD.t537 VDD.n2132 60.3596
R1545 VDD.n634 VDD.n87 60.0005
R1546 VDD.n1625 VDD.t492 58.4849
R1547 VDD.n1810 VDD.t730 58.4849
R1548 VDD.n1544 VDD.t234 58.4849
R1549 VDD.n1963 VDD.t34 58.4849
R1550 VDD.n1463 VDD.t587 58.4849
R1551 VDD.n1116 VDD.t23 58.4849
R1552 VDD.n955 VDD.t128 58.4849
R1553 VDD.n1274 VDD.t44 58.4849
R1554 VDD.n1031 VDD.t269 58.4849
R1555 VDD.n107 VDD.t555 58.4849
R1556 VDD.n504 VDD.t434 58.4849
R1557 VDD.n415 VDD.t19 58.4849
R1558 VDD.n326 VDD.t464 58.4849
R1559 VDD.n2284 VDD.t228 58.4849
R1560 VDD.n2416 VDD.t100 58.4849
R1561 VDD.n2540 VDD.t318 58.4849
R1562 VDD.n2664 VDD.t338 58.4849
R1563 VDD.n2673 VDD.t263 58.4849
R1564 VDD.n1357 VDD.n1355 57.7084
R1565 VDD.t667 VDD.n1380 56.794
R1566 VDD.n1443 VDD.t578 56.794
R1567 VDD.n2304 VDD.n2303 56.4711
R1568 VDD.n2092 VDD 55.6885
R1569 VDD.t576 VDD.n28 54.658
R1570 VDD.n603 VDD.t372 52.0553
R1571 VDD.t366 VDD.n616 52.0553
R1572 VDD.t349 VDD.n848 49.0494
R1573 VDD.t493 VDD.n1712 47.5005
R1574 VDD.n1714 VDD.t205 47.5005
R1575 VDD.n1781 VDD.t725 47.5005
R1576 VDD.t556 VDD.n1793 47.5005
R1577 VDD.t229 VDD.n1865 47.5005
R1578 VDD.n1867 VDD.t203 47.5005
R1579 VDD.n1934 VDD.t35 47.5005
R1580 VDD.t91 VDD.n1946 47.5005
R1581 VDD.t590 VDD.n2018 47.5005
R1582 VDD.n2020 VDD.t485 47.5005
R1583 VDD.n2702 VDD.t471 47.3689
R1584 VDD.n2716 VDD.t258 47.3689
R1585 VDD.n2637 VDD.t133 47.3689
R1586 VDD.n2623 VDD.t335 47.3689
R1587 VDD.n2513 VDD.t546 47.3689
R1588 VDD.n2499 VDD.t319 47.3689
R1589 VDD.n2389 VDD.t421 47.3689
R1590 VDD.n2375 VDD.t103 47.3689
R1591 VDD.n2255 VDD.t535 47.3689
R1592 VDD.n2241 VDD.t225 47.3689
R1593 VDD.t461 VDD.n308 46.8498
R1594 VDD.t277 VDD.n309 46.8498
R1595 VDD.t16 VDD.n397 46.8498
R1596 VDD.t437 VDD.n398 46.8498
R1597 VDD.t431 VDD.n486 46.8498
R1598 VDD.t115 VDD.n487 46.8498
R1599 VDD.t552 VDD.n575 46.8498
R1600 VDD.t239 VDD.n576 46.8498
R1601 VDD.t364 VDD.n667 46.8498
R1602 VDD.t594 VDD.n1049 46.4679
R1603 VDD.n1062 VDD.t264 46.4679
R1604 VDD.n1135 VDD.t310 46.4679
R1605 VDD.n1147 VDD.t20 46.4679
R1606 VDD.t621 VDD.n1207 46.4679
R1607 VDD.n1220 VDD.t131 46.4679
R1608 VDD.n1293 VDD.t639 46.4679
R1609 VDD.n1421 VDD.t580 46.4679
R1610 VDD.n2170 VDD 44.6138
R1611 VDD.n633 VDD.n632 44.2471
R1612 VDD.n761 VDD 44.2471
R1613 VDD.t350 VDD.n1323 43.8864
R1614 VDD.n1457 VDD 43.8864
R1615 VDD.n819 VDD 43.6491
R1616 VDD.n2067 VDD.t414 42.3555
R1617 VDD VDD.n2795 42.1058
R1618 VDD.n2550 VDD 42.1058
R1619 VDD.n2426 VDD 42.1058
R1620 VDD.n2306 VDD.n2305 42.1058
R1621 VDD.n2294 VDD 42.1058
R1622 VDD.n2179 VDD 42.1058
R1623 VDD.n2121 VDD.t501 41.9894
R1624 VDD.n2159 VDD 41.9894
R1625 VDD.t596 VDD.n736 41.6443
R1626 VDD.n750 VDD 41.6443
R1627 VDD.n2095 VDD.t405 41.5552
R1628 VDD.n2095 VDD.t519 41.5552
R1629 VDD.n2087 VDD.t309 41.5552
R1630 VDD.n2087 VDD.t5 41.5552
R1631 VDD.n1742 VDD.t214 41.5552
R1632 VDD.n1742 VDD.t528 41.5552
R1633 VDD.n1582 VDD.t403 41.5552
R1634 VDD.n1582 VDD.t324 41.5552
R1635 VDD.n1895 VDD.t410 41.5552
R1636 VDD.n1895 VDD.t219 41.5552
R1637 VDD.n1501 VDD.t632 41.5552
R1638 VDD.n1501 VDD.t532 41.5552
R1639 VDD.n1663 VDD.t291 41.5552
R1640 VDD.n1663 VDD.t307 41.5552
R1641 VDD.n1105 VDD.t255 41.5552
R1642 VDD.n1105 VDD.t523 41.5552
R1643 VDD.n962 VDD.t56 41.5552
R1644 VDD.n962 VDD.t549 41.5552
R1645 VDD.n1263 VDD.t609 41.5552
R1646 VDD.n1263 VDD.t10 41.5552
R1647 VDD.n1436 VDD.t399 41.5552
R1648 VDD.n1436 VDD.t579 41.5552
R1649 VDD.n138 VDD.t688 41.5552
R1650 VDD.n138 VDD.t67 41.5552
R1651 VDD.n173 VDD.t692 41.5552
R1652 VDD.n173 VDD.t682 41.5552
R1653 VDD.n208 VDD.t696 41.5552
R1654 VDD.n208 VDD.t346 41.5552
R1655 VDD.n243 VDD.t634 41.5552
R1656 VDD.n243 VDD.t3 41.5552
R1657 VDD.n2176 VDD.t507 41.5552
R1658 VDD.n2176 VDD.t694 41.5552
R1659 VDD.n9 VDD.t301 41.5552
R1660 VDD.n9 VDD.t686 41.5552
R1661 VDD.n5 VDD.t736 41.5552
R1662 VDD.n5 VDD.t684 41.5552
R1663 VDD.n1 VDD.t708 41.5552
R1664 VDD.n1 VDD.t626 41.5552
R1665 VDD.n2789 VDD.t286 41.5552
R1666 VDD.n2789 VDD.t690 41.5552
R1667 VDD VDD.n1110 41.3048
R1668 VDD.n1184 VDD 41.3048
R1669 VDD VDD.n1268 41.3048
R1670 VDD.t715 VDD.n785 41.0816
R1671 VDD.n804 VDD 41.0816
R1672 VDD.n1650 VDD.t208 38.6969
R1673 VDD.n1606 VDD.t559 38.6969
R1674 VDD.n1569 VDD.t202 38.6969
R1675 VDD.n1525 VDD.t90 38.6969
R1676 VDD.n1488 VDD.t488 38.6969
R1677 VDD.n1074 VDD.t593 38.6969
R1678 VDD.n977 VDD.t313 38.6969
R1679 VDD.n1232 VDD.t620 38.6969
R1680 VDD.n1356 VDD.t638 38.6969
R1681 VDD.n125 VDD.t238 38.6969
R1682 VDD.n160 VDD.t118 38.6969
R1683 VDD.n195 VDD.t440 38.6969
R1684 VDD.n230 VDD.t280 38.6969
R1685 VDD.n2220 VDD.t534 38.6969
R1686 VDD.n2354 VDD.t420 38.6969
R1687 VDD.n2478 VDD.t545 38.6969
R1688 VDD.n2602 VDD.t136 38.6969
R1689 VDD.n2735 VDD.t470 38.6969
R1690 VDD.n2050 VDD.t563 36.1587
R1691 VDD.n2050 VDD.t282 36.1587
R1692 VDD.n769 VDD.t607 36.1587
R1693 VDD.n769 VDD.t605 36.1587
R1694 VDD.n13 VDD.t212 36.1587
R1695 VDD.n13 VDD.t236 36.1587
R1696 VDD.t77 VDD.n880 36.1418
R1697 VDD.n1351 VDD.t637 36.1418
R1698 VDD.n1434 VDD.t398 36.1418
R1699 VDD.n1311 VDD.n900 35.2946
R1700 VDD.n1322 VDD.n894 35.2946
R1701 VDD.n1327 VDD.n888 35.2946
R1702 VDD.n1339 VDD.n887 35.2946
R1703 VDD.n1348 VDD.n879 35.2946
R1704 VDD.n878 VDD.n874 35.2946
R1705 VDD.n1368 VDD.n873 35.2946
R1706 VDD.n1378 VDD.n865 35.2946
R1707 VDD.n1393 VDD.n856 35.2946
R1708 VDD.n1405 VDD.n855 35.2946
R1709 VDD.n1415 VDD.n846 35.2946
R1710 VDD.n1431 VDD.n837 35.2946
R1711 VDD.n1446 VDD.n826 35.2946
R1712 VDD.n87 VDD.n81 35.2946
R1713 VDD.n646 VDD.n80 35.2946
R1714 VDD.n654 VDD.n72 35.2946
R1715 VDD.n666 VDD.n65 35.2946
R1716 VDD.n671 VDD.n58 35.2946
R1717 VDD.n684 VDD.n57 35.2946
R1718 VDD.n692 VDD.n50 35.2946
R1719 VDD.n704 VDD.n43 35.2946
R1720 VDD.n709 VDD.n36 35.2946
R1721 VDD.n722 VDD.n35 35.2946
R1722 VDD.n733 VDD.n27 35.2946
R1723 VDD.n1691 VDD.t731 34.3061
R1724 VDD.t617 VDD.n1609 34.3061
R1725 VDD.n1844 VDD.t629 34.3061
R1726 VDD.t384 VDD.n1528 34.3061
R1727 VDD.n1997 VDD.t105 34.3061
R1728 VDD.n2212 VDD.t443 34.211
R1729 VDD.n271 VDD.t170 33.8361
R1730 VDD.n360 VDD.t176 33.8361
R1731 VDD.n449 VDD.t155 33.8361
R1732 VDD.n538 VDD.t140 33.8361
R1733 VDD.n719 VDD.t570 33.8361
R1734 VDD.t83 VDD.n1083 33.5603
R1735 VDD.n1159 VDD.t516 33.5603
R1736 VDD.t250 VDD.n1241 33.5603
R1737 VDD.n1625 VDD.t61 31.831
R1738 VDD.n1810 VDD.t222 31.831
R1739 VDD.n1544 VDD.t340 31.831
R1740 VDD.n1963 VDD.t742 31.831
R1741 VDD.n1463 VDD.t678 31.831
R1742 VDD.n1116 VDD.t665 31.831
R1743 VDD.n955 VDD.t468 31.831
R1744 VDD.n1274 VDD.t59 31.831
R1745 VDD.n1031 VDD.t642 31.831
R1746 VDD.n107 VDD.t126 31.831
R1747 VDD.n504 VDD.t39 31.831
R1748 VDD.n415 VDD.t86 31.831
R1749 VDD.n326 VDD.t7 31.831
R1750 VDD.n2284 VDD.t718 31.831
R1751 VDD.n2416 VDD.t720 31.831
R1752 VDD.n2540 VDD.t452 31.831
R1753 VDD.n2664 VDD.t242 31.831
R1754 VDD.n2673 VDD.t458 31.831
R1755 VDD.n2111 VDD.t4 31.4922
R1756 VDD.n2124 VDD.t538 31.4922
R1757 VDD.n602 VDD.t358 31.2334
R1758 VDD.n617 VDD.t356 31.2334
R1759 VDD.n2070 VDD.t418 30.5947
R1760 VDD.n1402 VDD.t400 28.3972
R1761 VDD.n1471 VDD.t589 28.0332
R1762 VDD.n1510 VDD.t32 28.0332
R1763 VDD.n1552 VDD.t232 28.0332
R1764 VDD.n1591 VDD.t728 28.0332
R1765 VDD.n1633 VDD.t496 28.0332
R1766 VDD.n1284 VDD.t46 28.0332
R1767 VDD.n952 VDD.t130 28.0332
R1768 VDD.n1126 VDD.t25 28.0332
R1769 VDD.n1028 VDD.t267 28.0332
R1770 VDD.n217 VDD.t460 28.0332
R1771 VDD.n182 VDD.t15 28.0332
R1772 VDD.n147 VDD.t430 28.0332
R1773 VDD.n112 VDD.t551 28.0332
R1774 VDD.n2272 VDD.t224 28.0332
R1775 VDD.n2404 VDD.t102 28.0332
R1776 VDD.n2528 VDD.t316 28.0332
R1777 VDD.n2652 VDD.t334 28.0332
R1778 VDD.n2689 VDD.t261 28.0332
R1779 VDD.n2067 VDD.t412 26.5955
R1780 VDD.n2060 VDD.t194 26.5955
R1781 VDD.n2060 VDD.t196 26.5955
R1782 VDD.n2056 VDD.t192 26.5955
R1783 VDD.n2056 VDD.t561 26.5955
R1784 VDD.n776 VDD.t710 26.5955
R1785 VDD.n776 VDD.t454 26.5955
R1786 VDD.n781 VDD.t712 26.5955
R1787 VDD.n781 VDD.t714 26.5955
R1788 VDD.n37 VDD.t567 26.5955
R1789 VDD.n37 VDD.t571 26.5955
R1790 VDD.n49 VDD.t569 26.5955
R1791 VDD.n49 VDD.t573 26.5955
R1792 VDD.n59 VDD.t355 26.5955
R1793 VDD.n59 VDD.t575 26.5955
R1794 VDD.n71 VDD.t377 26.5955
R1795 VDD.n71 VDD.t365 26.5955
R1796 VDD.n77 VDD.t379 26.5955
R1797 VDD.n77 VDD.t369 26.5955
R1798 VDD.n84 VDD.t383 26.5955
R1799 VDD.n84 VDD.t371 26.5955
R1800 VDD.n89 VDD.t353 26.5955
R1801 VDD.n89 VDD.t363 26.5955
R1802 VDD.n619 VDD.t357 26.5955
R1803 VDD.n619 VDD.t367 26.5955
R1804 VDD.n97 VDD.t381 26.5955
R1805 VDD.n97 VDD.t375 26.5955
R1806 VDD.n605 VDD.t373 26.5955
R1807 VDD.n605 VDD.t359 26.5955
R1808 VDD.n24 VDD.t603 26.5955
R1809 VDD.n24 VDD.t599 26.5955
R1810 VDD.n19 VDD.t601 26.5955
R1811 VDD.n19 VDD.t661 26.5955
R1812 VDD.n632 VDD.n631 26.0279
R1813 VDD.n645 VDD.n644 26.0279
R1814 VDD.n656 VDD.n655 26.0279
R1815 VDD.n667 VDD.n64 26.0279
R1816 VDD.n670 VDD.n669 26.0279
R1817 VDD.n669 VDD.t354 26.0279
R1818 VDD.n683 VDD.n682 26.0279
R1819 VDD.n705 VDD.n42 26.0279
R1820 VDD.n708 VDD.n707 26.0279
R1821 VDD.n721 VDD.n720 26.0279
R1822 VDD.n735 VDD.n734 26.0279
R1823 VDD.n1297 VDD.n1295 25.8157
R1824 VDD.n1323 VDD.n893 25.8157
R1825 VDD.n1326 VDD.n1325 25.8157
R1826 VDD.n1338 VDD.n1337 25.8157
R1827 VDD.n1350 VDD.n1349 25.8157
R1828 VDD.n1352 VDD.n1351 25.8157
R1829 VDD.n1367 VDD.n1366 25.8157
R1830 VDD.n1380 VDD.n1379 25.8157
R1831 VDD.n1389 VDD.n861 25.8157
R1832 VDD.n1392 VDD.n1391 25.8157
R1833 VDD.n1404 VDD.n1403 25.8157
R1834 VDD.n1417 VDD.n1416 25.8157
R1835 VDD.n1420 VDD.n1419 25.8157
R1836 VDD.n1433 VDD.n1432 25.8157
R1837 VDD.n1442 VDD.n832 25.8157
R1838 VDD.n1445 VDD.n1444 25.8157
R1839 VDD.n1296 VDD.n910 24.7064
R1840 VDD.n1311 VDD.n902 24.7064
R1841 VDD.n1315 VDD.n894 24.7064
R1842 VDD.n1327 VDD.n892 24.7064
R1843 VDD.n1335 VDD.n887 24.7064
R1844 VDD.n1348 VDD.n881 24.7064
R1845 VDD.n1364 VDD.n873 24.7064
R1846 VDD.n1378 VDD.n867 24.7064
R1847 VDD.n1382 VDD.n862 24.7064
R1848 VDD.n1393 VDD.n860 24.7064
R1849 VDD.n1401 VDD.n855 24.7064
R1850 VDD.n1415 VDD.n849 24.7064
R1851 VDD.n1422 VDD.n847 24.7064
R1852 VDD.n1431 VDD.n839 24.7064
R1853 VDD.n1435 VDD.n833 24.7064
R1854 VDD.n1446 VDD.n831 24.7064
R1855 VDD.n642 VDD.n80 24.7064
R1856 VDD.n654 VDD.n74 24.7064
R1857 VDD.n658 VDD.n65 24.7064
R1858 VDD.n671 VDD.n63 24.7064
R1859 VDD.n680 VDD.n57 24.7064
R1860 VDD.n692 VDD.n52 24.7064
R1861 VDD.n696 VDD.n43 24.7064
R1862 VDD.n709 VDD.n41 24.7064
R1863 VDD.n718 VDD.n35 24.7064
R1864 VDD.n733 VDD.n29 24.7064
R1865 VDD.n2155 VDD.n2059 24.1595
R1866 VDD.n1440 VDD.n833 24.0258
R1867 VDD.n847 VDD.n844 24.0139
R1868 VDD.n1296 VDD.n906 23.9985
R1869 VDD.n1387 VDD.n862 23.9985
R1870 VDD.n1313 VDD.t47 23.2342
R1871 VDD.n1325 VDD.t401 23.2342
R1872 VDD.t72 VDD.n1642 21.1116
R1873 VDD.n1779 VDD.t331 21.1116
R1874 VDD.t87 VDD.n1561 21.1116
R1875 VDD.n1932 VDD.t199 21.1116
R1876 VDD.t216 VDD.n1480 21.1116
R1877 VDD.n2720 VDD.t123 21.0531
R1878 VDD.n2619 VDD.t490 21.0531
R1879 VDD.n2495 VDD.t408 21.0531
R1880 VDD.n2371 VDD.t505 21.0531
R1881 VDD.n2237 VDD.t724 21.0531
R1882 VDD.t247 VDD.n2112 20.995
R1883 VDD.t502 VDD.n222 20.8224
R1884 VDD.t209 VDD.n187 20.8224
R1885 VDD.t481 VDD.n152 20.8224
R1886 VDD.t436 VDD.n117 20.8224
R1887 VDD.n1061 VDD.t520 20.6527
R1888 VDD.t700 VDD.n1148 20.6527
R1889 VDD.n1219 VDD.t272 20.6527
R1890 VDD.t669 VDD.n1298 20.6527
R1891 VDD.n1444 VDD 20.6527
R1892 VDD.n2104 VDD.n2090 20.3039
R1893 VDD.n2104 VDD.n2086 20.3039
R1894 VDD.n2108 VDD.n2086 20.3039
R1895 VDD.n2115 VDD.n2083 20.3039
R1896 VDD.n2115 VDD.n2081 20.3039
R1897 VDD.n2119 VDD.n2081 20.3039
R1898 VDD.n2126 VDD.n2074 20.3039
R1899 VDD.n2130 VDD.n2074 20.3039
R1900 VDD.n2130 VDD.n2075 20.3039
R1901 VDD.n2137 VDD.n2066 20.3039
R1902 VDD.n2141 VDD.n2066 20.3039
R1903 VDD.n2147 VDD.n2063 20.3039
R1904 VDD.n2163 VDD.n2162 20.3039
R1905 VDD.n1681 VDD.n1658 20.3039
R1906 VDD.n1681 VDD.n1656 20.3039
R1907 VDD.n1694 VDD.n1653 20.3039
R1908 VDD.n1695 VDD.n1694 20.3039
R1909 VDD.n1698 VDD.n1646 20.3039
R1910 VDD.n1703 VDD.n1646 20.3039
R1911 VDD.n1703 VDD.n1644 20.3039
R1912 VDD.n1710 VDD.n1644 20.3039
R1913 VDD.n1718 VDD.n1717 20.3039
R1914 VDD.n1731 VDD.n1631 20.3039
R1915 VDD.n1738 VDD.n1623 20.3039
R1916 VDD.n1756 VDD.n1618 20.3039
R1917 VDD.n1756 VDD.n1615 20.3039
R1918 VDD.n1767 VDD.n1611 20.3039
R1919 VDD.n1767 VDD.n1612 20.3039
R1920 VDD.n1773 VDD.n1604 20.3039
R1921 VDD.n1777 VDD.n1604 20.3039
R1922 VDD.n1777 VDD.n1600 20.3039
R1923 VDD.n1783 VDD.n1600 20.3039
R1924 VDD.n1790 VDD.n1598 20.3039
R1925 VDD.n1808 VDD.n1588 20.3039
R1926 VDD.n1815 VDD.n1583 20.3039
R1927 VDD.n1834 VDD.n1577 20.3039
R1928 VDD.n1834 VDD.n1575 20.3039
R1929 VDD.n1847 VDD.n1572 20.3039
R1930 VDD.n1848 VDD.n1847 20.3039
R1931 VDD.n1851 VDD.n1565 20.3039
R1932 VDD.n1856 VDD.n1565 20.3039
R1933 VDD.n1856 VDD.n1563 20.3039
R1934 VDD.n1863 VDD.n1563 20.3039
R1935 VDD.n1871 VDD.n1870 20.3039
R1936 VDD.n1884 VDD.n1550 20.3039
R1937 VDD.n1891 VDD.n1542 20.3039
R1938 VDD.n1909 VDD.n1537 20.3039
R1939 VDD.n1909 VDD.n1534 20.3039
R1940 VDD.n1920 VDD.n1530 20.3039
R1941 VDD.n1920 VDD.n1531 20.3039
R1942 VDD.n1926 VDD.n1523 20.3039
R1943 VDD.n1930 VDD.n1523 20.3039
R1944 VDD.n1930 VDD.n1519 20.3039
R1945 VDD.n1936 VDD.n1519 20.3039
R1946 VDD.n1943 VDD.n1517 20.3039
R1947 VDD.n1961 VDD.n1507 20.3039
R1948 VDD.n1968 VDD.n1502 20.3039
R1949 VDD.n1987 VDD.n1496 20.3039
R1950 VDD.n1987 VDD.n1494 20.3039
R1951 VDD.n2000 VDD.n1491 20.3039
R1952 VDD.n2001 VDD.n2000 20.3039
R1953 VDD.n2004 VDD.n1484 20.3039
R1954 VDD.n2009 VDD.n1484 20.3039
R1955 VDD.n2009 VDD.n1482 20.3039
R1956 VDD.n2016 VDD.n1482 20.3039
R1957 VDD.n2024 VDD.n2023 20.3039
R1958 VDD.n2037 VDD.n1469 20.3039
R1959 VDD.n1041 VDD.n1027 20.3039
R1960 VDD.n1057 VDD.n1022 20.3039
R1961 VDD.n1064 VDD.n1015 20.3039
R1962 VDD.n1068 VDD.n1015 20.3039
R1963 VDD.n1068 VDD.n1012 20.3039
R1964 VDD.n1076 VDD.n1012 20.3039
R1965 VDD.n1080 VDD.n1010 20.3039
R1966 VDD.n1080 VDD.n1007 20.3039
R1967 VDD.n1092 VDD.n1004 20.3039
R1968 VDD.n1092 VDD.n1001 20.3039
R1969 VDD.n1114 VDD.n996 20.3039
R1970 VDD.n1120 VDD.n992 20.3039
R1971 VDD.n1139 VDD.n985 20.3039
R1972 VDD.n1145 VDD.n980 20.3039
R1973 VDD.n1151 VDD.n980 20.3039
R1974 VDD.n1151 VDD.n976 20.3039
R1975 VDD.n1155 VDD.n976 20.3039
R1976 VDD.n1162 VDD.n973 20.3039
R1977 VDD.n1162 VDD.n971 20.3039
R1978 VDD.n1175 VDD.n968 20.3039
R1979 VDD.n1175 VDD.n966 20.3039
R1980 VDD.n1192 VDD.n960 20.3039
R1981 VDD.n1199 VDD.n951 20.3039
R1982 VDD.n1215 VDD.n946 20.3039
R1983 VDD.n1222 VDD.n939 20.3039
R1984 VDD.n1226 VDD.n939 20.3039
R1985 VDD.n1226 VDD.n936 20.3039
R1986 VDD.n1234 VDD.n936 20.3039
R1987 VDD.n1238 VDD.n934 20.3039
R1988 VDD.n1238 VDD.n931 20.3039
R1989 VDD.n1250 VDD.n928 20.3039
R1990 VDD.n1250 VDD.n925 20.3039
R1991 VDD.n1272 VDD.n920 20.3039
R1992 VDD.n1278 VDD.n916 20.3039
R1993 VDD.n1301 VDD.n908 20.3039
R1994 VDD.n1453 VDD.n828 20.3039
R1995 VDD.n598 VDD.n104 20.3039
R1996 VDD.n607 VDD.n100 20.3039
R1997 VDD.n611 VDD.n96 20.3039
R1998 VDD.n621 VDD.n92 20.3039
R1999 VDD.n625 VDD.n90 20.3039
R2000 VDD.n754 VDD.n753 20.3039
R2001 VDD.n592 VDD.n109 20.3039
R2002 VDD.n568 VDD.n567 20.3039
R2003 VDD.n509 VDD.n139 20.3039
R2004 VDD.n528 VDD.n133 20.3039
R2005 VDD.n528 VDD.n131 20.3039
R2006 VDD.n541 VDD.n128 20.3039
R2007 VDD.n542 VDD.n541 20.3039
R2008 VDD.n545 VDD.n121 20.3039
R2009 VDD.n550 VDD.n121 20.3039
R2010 VDD.n550 VDD.n119 20.3039
R2011 VDD.n573 VDD.n119 20.3039
R2012 VDD.n502 VDD.n144 20.3039
R2013 VDD.n479 VDD.n478 20.3039
R2014 VDD.n420 VDD.n174 20.3039
R2015 VDD.n439 VDD.n168 20.3039
R2016 VDD.n439 VDD.n166 20.3039
R2017 VDD.n452 VDD.n163 20.3039
R2018 VDD.n453 VDD.n452 20.3039
R2019 VDD.n456 VDD.n156 20.3039
R2020 VDD.n461 VDD.n156 20.3039
R2021 VDD.n461 VDD.n154 20.3039
R2022 VDD.n484 VDD.n154 20.3039
R2023 VDD.n413 VDD.n179 20.3039
R2024 VDD.n390 VDD.n389 20.3039
R2025 VDD.n331 VDD.n209 20.3039
R2026 VDD.n350 VDD.n203 20.3039
R2027 VDD.n350 VDD.n201 20.3039
R2028 VDD.n363 VDD.n198 20.3039
R2029 VDD.n364 VDD.n363 20.3039
R2030 VDD.n367 VDD.n191 20.3039
R2031 VDD.n372 VDD.n191 20.3039
R2032 VDD.n372 VDD.n189 20.3039
R2033 VDD.n395 VDD.n189 20.3039
R2034 VDD.n324 VDD.n214 20.3039
R2035 VDD.n301 VDD.n300 20.3039
R2036 VDD.n261 VDD.n238 20.3039
R2037 VDD.n261 VDD.n236 20.3039
R2038 VDD.n274 VDD.n233 20.3039
R2039 VDD.n275 VDD.n274 20.3039
R2040 VDD.n278 VDD.n226 20.3039
R2041 VDD.n283 VDD.n226 20.3039
R2042 VDD.n283 VDD.n224 20.3039
R2043 VDD.n306 VDD.n224 20.3039
R2044 VDD.n2292 VDD.n2291 20.3039
R2045 VDD.n2424 VDD.n2423 20.3039
R2046 VDD.n2548 VDD.n2547 20.3039
R2047 VDD.n2798 VDD.n2670 20.3039
R2048 VDD.n627 VDD.n85 19.8626
R2049 VDD.n2068 VDD.n2063 19.6419
R2050 VDD.n2075 VDD.n2071 19.2005
R2051 VDD.n2154 VDD.n2057 19.2005
R2052 VDD.n745 VDD.n20 19.2005
R2053 VDD.n1688 VDD.n1656 18.5384
R2054 VDD.n1762 VDD.n1615 18.5384
R2055 VDD.n1841 VDD.n1575 18.5384
R2056 VDD.n1915 VDD.n1534 18.5384
R2057 VDD.n1994 VDD.n1494 18.5384
R2058 VDD.n1087 VDD.n1004 18.5384
R2059 VDD.n1168 VDD.n968 18.5384
R2060 VDD.n1245 VDD.n928 18.5384
R2061 VDD.n535 VDD.n131 18.5384
R2062 VDD.n446 VDD.n166 18.5384
R2063 VDD.n357 VDD.n201 18.5384
R2064 VDD.n268 VDD.n236 18.5384
R2065 VDD.n644 VDD.n643 18.2197
R2066 VDD.n655 VDD.n73 18.2197
R2067 VDD.n657 VDD.n64 18.2197
R2068 VDD.n670 VDD.n668 18.2197
R2069 VDD.n682 VDD.n681 18.2197
R2070 VDD.n693 VDD.n51 18.2197
R2071 VDD.n708 VDD.n706 18.2197
R2072 VDD.n720 VDD.n719 18.2197
R2073 VDD.n734 VDD.n28 18.2197
R2074 VDD.n1298 VDD.n1297 18.0712
R2075 VDD.n1312 VDD.n901 18.0712
R2076 VDD.n1314 VDD.n893 18.0712
R2077 VDD.n1326 VDD.n1324 18.0712
R2078 VDD.n1337 VDD.n1336 18.0712
R2079 VDD.n1349 VDD.n880 18.0712
R2080 VDD.n1353 VDD.n1352 18.0712
R2081 VDD.n1366 VDD.n1365 18.0712
R2082 VDD.n1379 VDD.n866 18.0712
R2083 VDD.n1381 VDD.n861 18.0712
R2084 VDD.n1392 VDD.n1390 18.0712
R2085 VDD.n1403 VDD.n1402 18.0712
R2086 VDD.n1416 VDD.n848 18.0712
R2087 VDD.n1421 VDD.n1420 18.0712
R2088 VDD.n1432 VDD.n838 18.0712
R2089 VDD.n1434 VDD.n832 18.0712
R2090 VDD.n1445 VDD.n1443 18.0712
R2091 VDD.n808 VDD.n807 17.3181
R2092 VDD.n821 VDD.n770 17.3181
R2093 VDD.n2119 VDD.n2078 17.2143
R2094 VDD.n598 VDD.n105 17.2143
R2095 VDD.n627 VDD.n626 17.2143
R2096 VDD.n746 VDD.n23 16.9936
R2097 VDD.n1727 VDD.n1631 16.7993
R2098 VDD.n1801 VDD.n1588 16.7993
R2099 VDD.n1880 VDD.n1550 16.7993
R2100 VDD.n1954 VDD.n1507 16.7993
R2101 VDD.n2033 VDD.n1469 16.7993
R2102 VDD.n1045 VDD.n1027 16.7993
R2103 VDD.n1128 VDD.n992 16.7993
R2104 VDD.n1203 VDD.n951 16.7993
R2105 VDD.n1286 VDD.n916 16.7993
R2106 VDD.n585 VDD.n109 16.7993
R2107 VDD.n495 VDD.n144 16.7993
R2108 VDD.n406 VDD.n179 16.7993
R2109 VDD.n317 VDD.n214 16.7993
R2110 VDD.n2166 VDD 16.7729
R2111 VDD.n757 VDD 16.7729
R2112 VDD.n782 VDD.n777 16.1887
R2113 VDD.n774 VDD.n770 16.1887
R2114 VDD.n694 VDD.t568 15.6169
R2115 VDD.n1367 VDD.t624 15.4896
R2116 VDD.n808 VDD.n773 15.2476
R2117 VDD.n1717 VDD.n1640 15.2281
R2118 VDD.n1790 VDD.n1597 15.2281
R2119 VDD.n1870 VDD.n1559 15.2281
R2120 VDD.n1943 VDD.n1516 15.2281
R2121 VDD.n2023 VDD.n1478 15.2281
R2122 VDD.n1057 VDD.n1019 15.2281
R2123 VDD.n1139 VDD.n983 15.2281
R2124 VDD.n1215 VDD.n943 15.2281
R2125 VDD.n1731 VDD.n1627 15.0074
R2126 VDD.n1808 VDD.n1586 15.0074
R2127 VDD.n1884 VDD.n1546 15.0074
R2128 VDD.n1961 VDD.n1505 15.0074
R2129 VDD.n2037 VDD.n1465 15.0074
R2130 VDD.n1041 VDD.n1033 15.0074
R2131 VDD.n1120 VDD.n995 15.0074
R2132 VDD.n1199 VDD.n957 15.0074
R2133 VDD.n1278 VDD.n919 15.0074
R2134 VDD.n593 VDD.n592 15.0074
R2135 VDD.n502 VDD.n142 15.0074
R2136 VDD.n413 VDD.n177 15.0074
R2137 VDD.n324 VDD.n212 15.0074
R2138 VDD.n1355 VDD.n1354 14.9976
R2139 VDD.n792 VDD.n780 14.8711
R2140 VDD.n1301 VDD.n905 14.566
R2141 VDD.n1453 VDD.n827 14.3453
R2142 VDD.n636 VDD.n635 14.3453
R2143 VDD.n641 VDD.n639 14.3453
R2144 VDD.n740 VDD.n26 14.3453
R2145 VDD.n799 VDD.n798 13.9299
R2146 VDD.n607 VDD.n606 13.6833
R2147 VDD.n620 VDD.n90 13.6833
R2148 VDD.n289 VDD 13.6005
R2149 VDD.n378 VDD 13.6005
R2150 VDD.n467 VDD 13.6005
R2151 VDD.n556 VDD 13.6005
R2152 VDD.n2754 VDD 13.6005
R2153 VDD.n2590 VDD 13.6005
R2154 VDD.n2466 VDD 13.6005
R2155 VDD.n2342 VDD 13.6005
R2156 VDD.n2097 VDD.n2090 13.4626
R2157 VDD.n1668 VDD.n1662 13.4626
R2158 VDD.n1744 VDD.n1620 13.4626
R2159 VDD.n1821 VDD.n1581 13.4626
R2160 VDD.n1897 VDD.n1539 13.4626
R2161 VDD.n1974 VDD.n1500 13.4626
R2162 VDD.n1107 VDD.n999 13.4626
R2163 VDD.n1187 VDD.n963 13.4626
R2164 VDD.n1265 VDD.n923 13.4626
R2165 VDD.n515 VDD.n137 13.4626
R2166 VDD.n426 VDD.n172 13.4626
R2167 VDD.n337 VDD.n207 13.4626
R2168 VDD.n248 VDD.n242 13.4626
R2169 VDD.t207 VDD.n1648 13.1949
R2170 VDD.n1770 VDD.t558 13.1949
R2171 VDD.t201 VDD.n1567 13.1949
R2172 VDD.n1923 VDD.t89 13.1949
R2173 VDD.t487 VDD.n1486 13.1949
R2174 VDD.n2737 VDD.t469 13.1584
R2175 VDD.n2604 VDD.t135 13.1584
R2176 VDD.n2480 VDD.t544 13.1584
R2177 VDD.n2356 VDD.t419 13.1584
R2178 VDD.n2222 VDD.t533 13.1584
R2179 VDD.n2166 VDD.n2052 13.0212
R2180 VDD.n2172 VDD.n2052 13.0212
R2181 VDD.n757 VDD.n15 13.0212
R2182 VDD.n763 VDD.n15 13.0212
R2183 VDD.t279 VDD.n228 13.0142
R2184 VDD.t439 VDD.n193 13.0142
R2185 VDD.t117 VDD.n158 13.0142
R2186 VDD.t237 VDD.n123 13.0142
R2187 VDD.n706 VDD.t566 13.0142
R2188 VDD.n1071 VDD.t592 12.9081
R2189 VDD.t312 VDD.n1158 12.9081
R2190 VDD.n1229 VDD.t619 12.9081
R2191 VDD.n1317 VDD.n1316 12.8005
R2192 VDD.n896 VDD.n891 12.8005
R2193 VDD.n1334 VDD.n1333 12.8005
R2194 VDD.n1342 VDD.n882 12.8005
R2195 VDD.n1363 VDD.n1362 12.8005
R2196 VDD.n1371 VDD.n868 12.8005
R2197 VDD.n1386 VDD.n859 12.8005
R2198 VDD.n1400 VDD.n1399 12.8005
R2199 VDD.n1408 VDD.n850 12.8005
R2200 VDD.n649 VDD.n75 12.8005
R2201 VDD.n67 VDD.n62 12.8005
R2202 VDD.n687 VDD.n53 12.8005
R2203 VDD.n45 VDD.n40 12.8005
R2204 VDD.n725 VDD.n30 12.8005
R2205 VDD.n2097 VDD.n2093 12.5798
R2206 VDD.n1674 VDD.n1662 12.5798
R2207 VDD.n1674 VDD.n1658 12.5798
R2208 VDD.n1738 VDD.n1627 12.5798
R2209 VDD.n1744 VDD.n1623 12.5798
R2210 VDD.n1751 VDD.n1620 12.5798
R2211 VDD.n1751 VDD.n1618 12.5798
R2212 VDD.n1815 VDD.n1586 12.5798
R2213 VDD.n1821 VDD.n1583 12.5798
R2214 VDD.n1827 VDD.n1581 12.5798
R2215 VDD.n1827 VDD.n1577 12.5798
R2216 VDD.n1891 VDD.n1546 12.5798
R2217 VDD.n1897 VDD.n1542 12.5798
R2218 VDD.n1904 VDD.n1539 12.5798
R2219 VDD.n1904 VDD.n1537 12.5798
R2220 VDD.n1968 VDD.n1505 12.5798
R2221 VDD.n1974 VDD.n1502 12.5798
R2222 VDD.n1980 VDD.n1500 12.5798
R2223 VDD.n1980 VDD.n1496 12.5798
R2224 VDD.n2042 VDD.n1465 12.5798
R2225 VDD.n1668 VDD.n1667 12.5798
R2226 VDD.n1099 VDD.n1001 12.5798
R2227 VDD.n1099 VDD.n999 12.5798
R2228 VDD.n1107 VDD.n996 12.5798
R2229 VDD.n1114 VDD.n995 12.5798
R2230 VDD.n1180 VDD.n966 12.5798
R2231 VDD.n1180 VDD.n963 12.5798
R2232 VDD.n1187 VDD.n960 12.5798
R2233 VDD.n1192 VDD.n957 12.5798
R2234 VDD.n1257 VDD.n925 12.5798
R2235 VDD.n1257 VDD.n923 12.5798
R2236 VDD.n1265 VDD.n920 12.5798
R2237 VDD.n1272 VDD.n919 12.5798
R2238 VDD.n1035 VDD.n1033 12.5798
R2239 VDD.n593 VDD.n104 12.5798
R2240 VDD.n568 VDD.n564 12.5798
R2241 VDD.n509 VDD.n142 12.5798
R2242 VDD.n515 VDD.n139 12.5798
R2243 VDD.n521 VDD.n137 12.5798
R2244 VDD.n521 VDD.n133 12.5798
R2245 VDD.n479 VDD.n475 12.5798
R2246 VDD.n420 VDD.n177 12.5798
R2247 VDD.n426 VDD.n174 12.5798
R2248 VDD.n432 VDD.n172 12.5798
R2249 VDD.n432 VDD.n168 12.5798
R2250 VDD.n390 VDD.n386 12.5798
R2251 VDD.n331 VDD.n212 12.5798
R2252 VDD.n337 VDD.n209 12.5798
R2253 VDD.n343 VDD.n207 12.5798
R2254 VDD.n343 VDD.n203 12.5798
R2255 VDD.n301 VDD.n297 12.5798
R2256 VDD.n254 VDD.n242 12.5798
R2257 VDD.n254 VDD.n238 12.5798
R2258 VDD.n248 VDD.n247 12.5798
R2259 VDD.n2088 VDD.n2083 12.1384
R2260 VDD.n717 VDD.n716 12.1384
R2261 VDD.n1439 VDD.n834 11.6971
R2262 VDD.n661 VDD.n660 11.2557
R2263 VDD.n1666 VDD 11.0898
R2264 VDD.n246 VDD 11.0536
R2265 VDD.n296 VDD.n295 10.9416
R2266 VDD.n385 VDD.n384 10.9416
R2267 VDD.n474 VDD.n473 10.9416
R2268 VDD.n563 VDD.n562 10.9416
R2269 VDD.n1424 VDD.n843 10.8143
R2270 VDD.n828 VDD.n824 10.8143
R2271 VDD.n2110 VDD.t308 10.4977
R2272 VDD.t380 VDD.n613 10.4115
R2273 VDD.n614 VDD.t374 10.4115
R2274 VDD.t568 VDD.n693 10.4115
R2275 VDD.t572 VDD.n42 10.4115
R2276 VDD.n790 VDD.n784 10.1652
R2277 VDD.n611 VDD.n98 10.1522
R2278 VDD.n98 VDD.n92 10.1522
R2279 VDD.n1459 VDD.n824 9.49016
R2280 VDD.n2149 VDD.n2059 9.41227
R2281 VDD.n1451 VDD.n827 9.3005
R2282 VDD.n1448 VDD.n829 9.3005
R2283 VDD.n1448 VDD.n826 9.3005
R2284 VDD.n1444 VDD.n826 9.3005
R2285 VDD.n1439 VDD.n836 9.3005
R2286 VDD.n1442 VDD.n1441 9.3005
R2287 VDD.n1439 VDD.n835 9.3005
R2288 VDD.n1429 VDD.n1428 9.3005
R2289 VDD.n1429 VDD.n837 9.3005
R2290 VDD.n1433 VDD.n837 9.3005
R2291 VDD.n1426 VDD.n834 9.3005
R2292 VDD.n1424 VDD.n845 9.3005
R2293 VDD.n1419 VDD.n1418 9.3005
R2294 VDD.n1425 VDD.n1424 9.3005
R2295 VDD.n1413 VDD.n1412 9.3005
R2296 VDD.n1413 VDD.n846 9.3005
R2297 VDD.n1417 VDD.n846 9.3005
R2298 VDD.n1410 VDD.n843 9.3005
R2299 VDD.n1406 VDD.n854 9.3005
R2300 VDD.n1406 VDD.n1405 9.3005
R2301 VDD.n1405 VDD.n1404 9.3005
R2302 VDD.n1409 VDD.n1408 9.3005
R2303 VDD.n1396 VDD.n1395 9.3005
R2304 VDD.n1395 VDD.n856 9.3005
R2305 VDD.n1391 VDD.n856 9.3005
R2306 VDD.n1399 VDD.n1398 9.3005
R2307 VDD.n1386 VDD.n864 9.3005
R2308 VDD.n1389 VDD.n1388 9.3005
R2309 VDD.n1386 VDD.n858 9.3005
R2310 VDD.n1376 VDD.n1375 9.3005
R2311 VDD.n1376 VDD.n865 9.3005
R2312 VDD.n1380 VDD.n865 9.3005
R2313 VDD.n1373 VDD.n863 9.3005
R2314 VDD.n1369 VDD.n872 9.3005
R2315 VDD.n1369 VDD.n1368 9.3005
R2316 VDD.n1368 VDD.n1367 9.3005
R2317 VDD.n1372 VDD.n1371 9.3005
R2318 VDD.n1359 VDD.n1358 9.3005
R2319 VDD.n1358 VDD.n874 9.3005
R2320 VDD.n1351 VDD.n874 9.3005
R2321 VDD.n1362 VDD.n1361 9.3005
R2322 VDD.n1346 VDD.n1345 9.3005
R2323 VDD.n1346 VDD.n879 9.3005
R2324 VDD.n1350 VDD.n879 9.3005
R2325 VDD.n877 VDD.n876 9.3005
R2326 VDD.n1340 VDD.n886 9.3005
R2327 VDD.n1340 VDD.n1339 9.3005
R2328 VDD.n1339 VDD.n1338 9.3005
R2329 VDD.n1343 VDD.n1342 9.3005
R2330 VDD.n1330 VDD.n1329 9.3005
R2331 VDD.n1329 VDD.n888 9.3005
R2332 VDD.n1325 VDD.n888 9.3005
R2333 VDD.n1333 VDD.n1332 9.3005
R2334 VDD.n1321 VDD.n1320 9.3005
R2335 VDD.n1322 VDD.n1321 9.3005
R2336 VDD.n1323 VDD.n1322 9.3005
R2337 VDD.n896 VDD.n890 9.3005
R2338 VDD.n1309 VDD.n1308 9.3005
R2339 VDD.n1309 VDD.n900 9.3005
R2340 VDD.n1313 VDD.n900 9.3005
R2341 VDD.n1318 VDD.n1317 9.3005
R2342 VDD.n1306 VDD.n1303 9.3005
R2343 VDD.n1295 VDD.n1294 9.3005
R2344 VDD.n1307 VDD.n1306 9.3005
R2345 VDD.n810 VDD.n773 9.3005
R2346 VDD.n790 VDD.n789 9.3005
R2347 VDD.n295 VDD.n293 9.3005
R2348 VDD.n384 VDD.n382 9.3005
R2349 VDD.n473 VDD.n471 9.3005
R2350 VDD.n562 VDD.n560 9.3005
R2351 VDD.n727 VDD.n26 9.3005
R2352 VDD.n731 VDD.n730 9.3005
R2353 VDD.n731 VDD.n27 9.3005
R2354 VDD.n735 VDD.n27 9.3005
R2355 VDD.n723 VDD.n34 9.3005
R2356 VDD.n723 VDD.n722 9.3005
R2357 VDD.n722 VDD.n721 9.3005
R2358 VDD.n726 VDD.n725 9.3005
R2359 VDD.n712 VDD.n711 9.3005
R2360 VDD.n711 VDD.n36 9.3005
R2361 VDD.n707 VDD.n36 9.3005
R2362 VDD.n715 VDD.n714 9.3005
R2363 VDD.n703 VDD.n702 9.3005
R2364 VDD.n704 VDD.n703 9.3005
R2365 VDD.n705 VDD.n704 9.3005
R2366 VDD.n45 VDD.n39 9.3005
R2367 VDD.n690 VDD.n689 9.3005
R2368 VDD.n690 VDD.n50 9.3005
R2369 VDD.n694 VDD.n50 9.3005
R2370 VDD.n700 VDD.n699 9.3005
R2371 VDD.n685 VDD.n56 9.3005
R2372 VDD.n685 VDD.n684 9.3005
R2373 VDD.n684 VDD.n683 9.3005
R2374 VDD.n688 VDD.n687 9.3005
R2375 VDD.n674 VDD.n673 9.3005
R2376 VDD.n673 VDD.n58 9.3005
R2377 VDD.n669 VDD.n58 9.3005
R2378 VDD.n677 VDD.n676 9.3005
R2379 VDD.n665 VDD.n664 9.3005
R2380 VDD.n666 VDD.n665 9.3005
R2381 VDD.n667 VDD.n666 9.3005
R2382 VDD.n67 VDD.n61 9.3005
R2383 VDD.n652 VDD.n651 9.3005
R2384 VDD.n652 VDD.n72 9.3005
R2385 VDD.n656 VDD.n72 9.3005
R2386 VDD.n662 VDD.n661 9.3005
R2387 VDD.n647 VDD.n79 9.3005
R2388 VDD.n647 VDD.n646 9.3005
R2389 VDD.n646 VDD.n645 9.3005
R2390 VDD.n650 VDD.n649 9.3005
R2391 VDD.n639 VDD.n81 9.3005
R2392 VDD.n631 VDD.n81 9.3005
R2393 VDD.n2310 VDD.n2308 9.3005
R2394 VDD.n2308 VDD.n2307 9.3005
R2395 VDD.n1718 VDD.n1637 9.11136
R2396 VDD.n1598 VDD.n1594 9.11136
R2397 VDD.n1871 VDD.n1556 9.11136
R2398 VDD.n1517 VDD.n1513 9.11136
R2399 VDD.n2024 VDD.n1475 9.11136
R2400 VDD.n1052 VDD.n1022 9.11136
R2401 VDD.n990 VDD.n985 9.11136
R2402 VDD.n1210 VDD.n946 9.11136
R2403 VDD.n914 VDD.n908 9.11136
R2404 VDD.n567 VDD.n115 9.11136
R2405 VDD.n478 VDD.n150 9.11136
R2406 VDD.n389 VDD.n185 9.11136
R2407 VDD.n300 VDD.n220 9.11136
R2408 VDD.n2155 VDD.n2154 9.04877
R2409 VDD.n746 VDD.n745 9.04877
R2410 VDD.n290 VDD.n288 8.91563
R2411 VDD.n379 VDD.n377 8.91563
R2412 VDD.n468 VDD.n466 8.91563
R2413 VDD.n557 VDD.n555 8.91563
R2414 VDD.n1721 VDD.n1638 8.78856
R2415 VDD.n1798 VDD.n1797 8.78856
R2416 VDD.n1874 VDD.n1557 8.78856
R2417 VDD.n1951 VDD.n1950 8.78856
R2418 VDD.n2027 VDD.n1476 8.78856
R2419 VDD.n1053 VDD.n1024 8.78856
R2420 VDD.n1132 VDD.n989 8.78856
R2421 VDD.n1211 VDD.n948 8.78856
R2422 VDD.n1290 VDD.n913 8.78856
R2423 VDD.n581 VDD.n580 8.78856
R2424 VDD.n492 VDD.n491 8.78856
R2425 VDD.n403 VDD.n402 8.78856
R2426 VDD.n314 VDD.n313 8.78856
R2427 VDD.n1710 VDD.n1640 8.6074
R2428 VDD.n1783 VDD.n1597 8.6074
R2429 VDD.n1863 VDD.n1559 8.6074
R2430 VDD.n1936 VDD.n1516 8.6074
R2431 VDD.n2016 VDD.n1478 8.6074
R2432 VDD.n1064 VDD.n1019 8.6074
R2433 VDD.n1145 VDD.n983 8.6074
R2434 VDD.n1222 VDD.n943 8.6074
R2435 VDD.n698 VDD.n697 8.6074
R2436 VDD.n573 VDD.n572 8.6074
R2437 VDD.n484 VDD.n483 8.6074
R2438 VDD.n395 VDD.n394 8.6074
R2439 VDD.n306 VDD.n305 8.6074
R2440 VDD.n1034 VDD.n1033 8.47522
R2441 VDD.n593 VDD.n108 8.47522
R2442 VDD.n142 VDD.n141 8.47522
R2443 VDD.n177 VDD.n176 8.47522
R2444 VDD.n212 VDD.n211 8.47522
R2445 VDD.n2676 VDD.n2675 8.47522
R2446 VDD.n1466 VDD.n1465 8.47518
R2447 VDD.n1505 VDD.n1504 8.47518
R2448 VDD.n1547 VDD.n1546 8.47518
R2449 VDD.n1586 VDD.n1585 8.47518
R2450 VDD.n1628 VDD.n1627 8.47518
R2451 VDD.n919 VDD.n918 8.47518
R2452 VDD.n958 VDD.n957 8.47518
R2453 VDD.n995 VDD.n994 8.47518
R2454 VDD.n2287 VDD.n2286 8.47518
R2455 VDD.n2419 VDD.n2418 8.47518
R2456 VDD.n2543 VDD.n2542 8.47518
R2457 VDD.n2667 VDD.n2666 8.47518
R2458 VDD.n2053 VDD.n2052 8.47281
R2459 VDD.n1668 VDD.n1664 8.47281
R2460 VDD.n248 VDD.n244 8.47281
R2461 VDD.n2156 VDD.n2155 8.47276
R2462 VDD.n1974 VDD.n1973 8.47276
R2463 VDD.n1898 VDD.n1897 8.47276
R2464 VDD.n1821 VDD.n1820 8.47276
R2465 VDD.n1745 VDD.n1744 8.47276
R2466 VDD.n1266 VDD.n1265 8.47276
R2467 VDD.n1187 VDD.n1186 8.47276
R2468 VDD.n1108 VDD.n1107 8.47276
R2469 VDD.n16 VDD.n15 8.47276
R2470 VDD.n747 VDD.n746 8.47276
R2471 VDD.n515 VDD.n514 8.47276
R2472 VDD.n426 VDD.n425 8.47276
R2473 VDD.n337 VDD.n336 8.47276
R2474 VDD.n2182 VDD.n2181 8.47276
R2475 VDD.n2297 VDD.n2296 8.47276
R2476 VDD.n2429 VDD.n2428 8.47276
R2477 VDD.n2553 VDD.n2552 8.47276
R2478 VDD.n2792 VDD.n2791 8.47276
R2479 VDD.n2098 VDD.n2097 8.47181
R2480 VDD.n2314 VDD.n2313 8.47164
R2481 VDD.n2438 VDD.n2437 8.47164
R2482 VDD.n2562 VDD.n2561 8.47164
R2483 VDD.n2780 VDD.n2779 8.47164
R2484 VDD.n1981 VDD.n1980 8.4716
R2485 VDD.n1904 VDD.n1903 8.4716
R2486 VDD.n1828 VDD.n1827 8.4716
R2487 VDD.n1751 VDD.n1750 8.4716
R2488 VDD.n1675 VDD.n1674 8.4716
R2489 VDD.n1257 VDD.n1256 8.4716
R2490 VDD.n1181 VDD.n1180 8.4716
R2491 VDD.n1099 VDD.n1098 8.4716
R2492 VDD.n522 VDD.n521 8.4716
R2493 VDD.n433 VDD.n432 8.4716
R2494 VDD.n344 VDD.n343 8.4716
R2495 VDD.n255 VDD.n254 8.4716
R2496 VDD.n2191 VDD.n2190 8.4716
R2497 VDD.n2079 VDD.n2078 8.47092
R2498 VDD.n2248 VDD.n2247 8.47011
R2499 VDD.n1479 VDD.n1478 8.47007
R2500 VDD.n1995 VDD.n1994 8.47007
R2501 VDD.n1516 VDD.n1515 8.47007
R2502 VDD.n1915 VDD.n1914 8.47007
R2503 VDD.n1560 VDD.n1559 8.47007
R2504 VDD.n1842 VDD.n1841 8.47007
R2505 VDD.n1597 VDD.n1596 8.47007
R2506 VDD.n1762 VDD.n1761 8.47007
R2507 VDD.n1641 VDD.n1640 8.47007
R2508 VDD.n1689 VDD.n1688 8.47007
R2509 VDD.n1245 VDD.n1244 8.47007
R2510 VDD.n944 VDD.n943 8.47007
R2511 VDD.n1169 VDD.n1168 8.47007
R2512 VDD.n983 VDD.n982 8.47007
R2513 VDD.n1087 VDD.n1086 8.47007
R2514 VDD.n1020 VDD.n1019 8.47007
R2515 VDD.n536 VDD.n535 8.47007
R2516 VDD.n447 VDD.n446 8.47007
R2517 VDD.n358 VDD.n357 8.47007
R2518 VDD.n269 VDD.n268 8.47007
R2519 VDD.n2209 VDD.n2208 8.47007
R2520 VDD.n2382 VDD.n2381 8.47007
R2521 VDD.n2506 VDD.n2505 8.47007
R2522 VDD.n2630 VDD.n2629 8.47007
R2523 VDD.n2713 VDD.n2712 8.47007
R2524 VDD.n2147 VDD.n2146 8.45089
R2525 VDD.n2146 VDD.n2145 8.45089
R2526 VDD.n2144 VDD.n2064 8.45089
R2527 VDD.n2143 VDD.n2142 8.45089
R2528 VDD.n2134 VDD.n2065 8.45089
R2529 VDD.n2136 VDD.n2135 8.45089
R2530 VDD.n2133 VDD.n2072 8.45089
R2531 VDD.n2132 VDD.n2131 8.45089
R2532 VDD.n2123 VDD.n2073 8.45089
R2533 VDD.n2125 VDD.n2124 8.45089
R2534 VDD.n2122 VDD.n2079 8.45089
R2535 VDD.n2121 VDD.n2120 8.45089
R2536 VDD.n2112 VDD.n2080 8.45089
R2537 VDD.n2114 VDD.n2113 8.45089
R2538 VDD.n2111 VDD.n2084 8.45089
R2539 VDD.n2110 VDD.n2109 8.45089
R2540 VDD.n2101 VDD.n2085 8.45089
R2541 VDD.n2103 VDD.n2102 8.45089
R2542 VDD.n2100 VDD.n2091 8.45089
R2543 VDD.n2099 VDD.n2098 8.45089
R2544 VDD.n2167 VDD.n2166 8.45089
R2545 VDD.n2168 VDD.n2167 8.45089
R2546 VDD.n2159 VDD.n2054 8.45089
R2547 VDD.n2161 VDD.n2160 8.45089
R2548 VDD.n2158 VDD.n2058 8.45089
R2549 VDD.n2157 VDD.n2156 8.45089
R2550 VDD.n2169 VDD.n2053 8.45089
R2551 VDD.n2172 VDD.n2171 8.45089
R2552 VDD.n2171 VDD.n2170 8.45089
R2553 VDD.n2042 VDD.n2041 8.45089
R2554 VDD.n2040 VDD.n1466 8.45089
R2555 VDD.n2039 VDD.n2038 8.45089
R2556 VDD.n1468 VDD.n1467 8.45089
R2557 VDD.n2032 VDD.n2031 8.45089
R2558 VDD.n2030 VDD.n1473 8.45089
R2559 VDD.n2029 VDD.n2028 8.45089
R2560 VDD.n2020 VDD.n1474 8.45089
R2561 VDD.n2022 VDD.n2021 8.45089
R2562 VDD.n2019 VDD.n1479 8.45089
R2563 VDD.n2018 VDD.n2017 8.45089
R2564 VDD.n1481 VDD.n1480 8.45089
R2565 VDD.n2008 VDD.t530 8.45089
R2566 VDD.n2007 VDD.n1485 8.45089
R2567 VDD.n2006 VDD.n2005 8.45089
R2568 VDD.n1487 VDD.n1486 8.45089
R2569 VDD.n1999 VDD.n1998 8.45089
R2570 VDD.n1997 VDD.n1492 8.45089
R2571 VDD.n1996 VDD.n1995 8.45089
R2572 VDD.n1984 VDD.n1493 8.45089
R2573 VDD.n1986 VDD.n1985 8.45089
R2574 VDD.n1983 VDD.n1497 8.45089
R2575 VDD.n1982 VDD.n1981 8.45089
R2576 VDD.n1499 VDD.n1498 8.45089
R2577 VDD.n1973 VDD.n1972 8.45089
R2578 VDD.n1971 VDD.n1503 8.45089
R2579 VDD.n1970 VDD.n1969 8.45089
R2580 VDD.n1958 VDD.n1504 8.45089
R2581 VDD.n1960 VDD.n1959 8.45089
R2582 VDD.n1957 VDD.n1508 8.45089
R2583 VDD.n1956 VDD.n1955 8.45089
R2584 VDD.n1947 VDD.n1509 8.45089
R2585 VDD.n1949 VDD.n1948 8.45089
R2586 VDD.n1946 VDD.n1514 8.45089
R2587 VDD.n1945 VDD.n1944 8.45089
R2588 VDD.n1933 VDD.n1515 8.45089
R2589 VDD.n1935 VDD.n1934 8.45089
R2590 VDD.n1932 VDD.n1520 8.45089
R2591 VDD.t220 VDD.n1931 8.45089
R2592 VDD.n1522 VDD.n1521 8.45089
R2593 VDD.n1925 VDD.n1924 8.45089
R2594 VDD.n1923 VDD.n1527 8.45089
R2595 VDD.n1922 VDD.n1921 8.45089
R2596 VDD.n1529 VDD.n1528 8.45089
R2597 VDD.n1914 VDD.n1913 8.45089
R2598 VDD.n1912 VDD.n1535 8.45089
R2599 VDD.n1911 VDD.n1910 8.45089
R2600 VDD.n1901 VDD.n1536 8.45089
R2601 VDD.n1903 VDD.n1902 8.45089
R2602 VDD.n1900 VDD.n1540 8.45089
R2603 VDD.n1899 VDD.n1898 8.45089
R2604 VDD.n1888 VDD.n1541 8.45089
R2605 VDD.n1890 VDD.n1889 8.45089
R2606 VDD.n1887 VDD.n1547 8.45089
R2607 VDD.n1886 VDD.n1885 8.45089
R2608 VDD.n1549 VDD.n1548 8.45089
R2609 VDD.n1879 VDD.n1878 8.45089
R2610 VDD.n1877 VDD.n1554 8.45089
R2611 VDD.n1876 VDD.n1875 8.45089
R2612 VDD.n1867 VDD.n1555 8.45089
R2613 VDD.n1869 VDD.n1868 8.45089
R2614 VDD.n1866 VDD.n1560 8.45089
R2615 VDD.n1865 VDD.n1864 8.45089
R2616 VDD.n1562 VDD.n1561 8.45089
R2617 VDD.n1855 VDD.t322 8.45089
R2618 VDD.n1854 VDD.n1566 8.45089
R2619 VDD.n1853 VDD.n1852 8.45089
R2620 VDD.n1568 VDD.n1567 8.45089
R2621 VDD.n1846 VDD.n1845 8.45089
R2622 VDD.n1844 VDD.n1573 8.45089
R2623 VDD.n1843 VDD.n1842 8.45089
R2624 VDD.n1831 VDD.n1574 8.45089
R2625 VDD.n1833 VDD.n1832 8.45089
R2626 VDD.n1830 VDD.n1578 8.45089
R2627 VDD.n1829 VDD.n1828 8.45089
R2628 VDD.n1580 VDD.n1579 8.45089
R2629 VDD.n1820 VDD.n1819 8.45089
R2630 VDD.n1818 VDD.n1584 8.45089
R2631 VDD.n1817 VDD.n1816 8.45089
R2632 VDD.n1805 VDD.n1585 8.45089
R2633 VDD.n1807 VDD.n1806 8.45089
R2634 VDD.n1804 VDD.n1589 8.45089
R2635 VDD.n1803 VDD.n1802 8.45089
R2636 VDD.n1794 VDD.n1590 8.45089
R2637 VDD.n1796 VDD.n1795 8.45089
R2638 VDD.n1793 VDD.n1595 8.45089
R2639 VDD.n1792 VDD.n1791 8.45089
R2640 VDD.n1780 VDD.n1596 8.45089
R2641 VDD.n1782 VDD.n1781 8.45089
R2642 VDD.n1779 VDD.n1601 8.45089
R2643 VDD.t525 VDD.n1778 8.45089
R2644 VDD.n1603 VDD.n1602 8.45089
R2645 VDD.n1772 VDD.n1771 8.45089
R2646 VDD.n1770 VDD.n1608 8.45089
R2647 VDD.n1769 VDD.n1768 8.45089
R2648 VDD.n1610 VDD.n1609 8.45089
R2649 VDD.n1761 VDD.n1760 8.45089
R2650 VDD.n1759 VDD.n1616 8.45089
R2651 VDD.n1758 VDD.n1757 8.45089
R2652 VDD.n1748 VDD.n1617 8.45089
R2653 VDD.n1750 VDD.n1749 8.45089
R2654 VDD.n1747 VDD.n1621 8.45089
R2655 VDD.n1746 VDD.n1745 8.45089
R2656 VDD.n1735 VDD.n1622 8.45089
R2657 VDD.n1737 VDD.n1736 8.45089
R2658 VDD.n1734 VDD.n1628 8.45089
R2659 VDD.n1733 VDD.n1732 8.45089
R2660 VDD.n1630 VDD.n1629 8.45089
R2661 VDD.n1726 VDD.n1725 8.45089
R2662 VDD.n1724 VDD.n1635 8.45089
R2663 VDD.n1723 VDD.n1722 8.45089
R2664 VDD.n1714 VDD.n1636 8.45089
R2665 VDD.n1716 VDD.n1715 8.45089
R2666 VDD.n1713 VDD.n1641 8.45089
R2667 VDD.n1712 VDD.n1711 8.45089
R2668 VDD.n1643 VDD.n1642 8.45089
R2669 VDD.n1702 VDD.t304 8.45089
R2670 VDD.n1701 VDD.n1647 8.45089
R2671 VDD.n1700 VDD.n1699 8.45089
R2672 VDD.n1649 VDD.n1648 8.45089
R2673 VDD.n1693 VDD.n1692 8.45089
R2674 VDD.n1691 VDD.n1654 8.45089
R2675 VDD.n1690 VDD.n1689 8.45089
R2676 VDD.n1678 VDD.n1655 8.45089
R2677 VDD.n1680 VDD.n1679 8.45089
R2678 VDD.n1677 VDD.n1659 8.45089
R2679 VDD.n1676 VDD.n1675 8.45089
R2680 VDD.n1661 VDD.n1660 8.45089
R2681 VDD.n1665 VDD.n1664 8.45089
R2682 VDD.n1667 VDD.n1666 8.45089
R2683 VDD.n1459 VDD.n1458 8.45089
R2684 VDD.n1458 VDD.n1457 8.45089
R2685 VDD.n1456 VDD.n825 8.45089
R2686 VDD.n1455 VDD.n1454 8.45089
R2687 VDD.n1300 VDD.n1299 8.45089
R2688 VDD.n1293 VDD.n909 8.45089
R2689 VDD.n1292 VDD.n1291 8.45089
R2690 VDD.n912 VDD.n911 8.45089
R2691 VDD.n1283 VDD.n1282 8.45089
R2692 VDD.n1281 VDD.n917 8.45089
R2693 VDD.n1280 VDD.n1279 8.45089
R2694 VDD.n1269 VDD.n918 8.45089
R2695 VDD.n1271 VDD.n1270 8.45089
R2696 VDD.n1268 VDD.n921 8.45089
R2697 VDD.n1267 VDD.n1266 8.45089
R2698 VDD.n1254 VDD.n922 8.45089
R2699 VDD.n1256 VDD.n1255 8.45089
R2700 VDD.n1253 VDD.n926 8.45089
R2701 VDD.n1252 VDD.n1251 8.45089
R2702 VDD.n1242 VDD.n927 8.45089
R2703 VDD.n1244 VDD.n1243 8.45089
R2704 VDD.n1241 VDD.n932 8.45089
R2705 VDD.n1240 VDD.n1239 8.45089
R2706 VDD.n1229 VDD.n933 8.45089
R2707 VDD.n1231 VDD.n1230 8.45089
R2708 VDD.n1228 VDD.n937 8.45089
R2709 VDD.t611 VDD.n1227 8.45089
R2710 VDD.n1219 VDD.n938 8.45089
R2711 VDD.n1221 VDD.n1220 8.45089
R2712 VDD.n1218 VDD.n944 8.45089
R2713 VDD.n1217 VDD.n1216 8.45089
R2714 VDD.n1207 VDD.n945 8.45089
R2715 VDD.n1209 VDD.n1208 8.45089
R2716 VDD.n1206 VDD.n949 8.45089
R2717 VDD.n1205 VDD.n1204 8.45089
R2718 VDD.n1196 VDD.n950 8.45089
R2719 VDD.n1198 VDD.n1197 8.45089
R2720 VDD.n1195 VDD.n958 8.45089
R2721 VDD.n1194 VDD.n1193 8.45089
R2722 VDD.n1184 VDD.n959 8.45089
R2723 VDD.n1186 VDD.n1185 8.45089
R2724 VDD.n1183 VDD.n964 8.45089
R2725 VDD.n1182 VDD.n1181 8.45089
R2726 VDD.n1172 VDD.n965 8.45089
R2727 VDD.n1174 VDD.n1173 8.45089
R2728 VDD.n1171 VDD.n969 8.45089
R2729 VDD.n1170 VDD.n1169 8.45089
R2730 VDD.n1159 VDD.n970 8.45089
R2731 VDD.n1161 VDD.n1160 8.45089
R2732 VDD.n1158 VDD.n974 8.45089
R2733 VDD.n1157 VDD.n1156 8.45089
R2734 VDD.n1149 VDD.n975 8.45089
R2735 VDD.n1150 VDD.t54 8.45089
R2736 VDD.n1148 VDD.n981 8.45089
R2737 VDD.n1147 VDD.n1146 8.45089
R2738 VDD.n1136 VDD.n982 8.45089
R2739 VDD.n1138 VDD.n1137 8.45089
R2740 VDD.n1135 VDD.n986 8.45089
R2741 VDD.n1134 VDD.n1133 8.45089
R2742 VDD.n988 VDD.n987 8.45089
R2743 VDD.n1125 VDD.n1124 8.45089
R2744 VDD.n1123 VDD.n993 8.45089
R2745 VDD.n1122 VDD.n1121 8.45089
R2746 VDD.n1111 VDD.n994 8.45089
R2747 VDD.n1113 VDD.n1112 8.45089
R2748 VDD.n1110 VDD.n997 8.45089
R2749 VDD.n1109 VDD.n1108 8.45089
R2750 VDD.n1096 VDD.n998 8.45089
R2751 VDD.n1098 VDD.n1097 8.45089
R2752 VDD.n1095 VDD.n1002 8.45089
R2753 VDD.n1094 VDD.n1093 8.45089
R2754 VDD.n1084 VDD.n1003 8.45089
R2755 VDD.n1086 VDD.n1085 8.45089
R2756 VDD.n1083 VDD.n1008 8.45089
R2757 VDD.n1082 VDD.n1081 8.45089
R2758 VDD.n1071 VDD.n1009 8.45089
R2759 VDD.n1073 VDD.n1072 8.45089
R2760 VDD.n1070 VDD.n1013 8.45089
R2761 VDD.t253 VDD.n1069 8.45089
R2762 VDD.n1061 VDD.n1014 8.45089
R2763 VDD.n1063 VDD.n1062 8.45089
R2764 VDD.n1060 VDD.n1020 8.45089
R2765 VDD.n1059 VDD.n1058 8.45089
R2766 VDD.n1049 VDD.n1021 8.45089
R2767 VDD.n1051 VDD.n1050 8.45089
R2768 VDD.n1048 VDD.n1025 8.45089
R2769 VDD.n1047 VDD.n1046 8.45089
R2770 VDD.n1038 VDD.n1026 8.45089
R2771 VDD.n1040 VDD.n1039 8.45089
R2772 VDD.n1037 VDD.n1034 8.45089
R2773 VDD.n1036 VDD.n1035 8.45089
R2774 VDD.n763 VDD.n762 8.45089
R2775 VDD.n762 VDD.n761 8.45089
R2776 VDD.n760 VDD.n16 8.45089
R2777 VDD.n759 VDD.n758 8.45089
R2778 VDD.n750 VDD.n17 8.45089
R2779 VDD.n752 VDD.n751 8.45089
R2780 VDD.n749 VDD.n21 8.45089
R2781 VDD.n748 VDD.n747 8.45089
R2782 VDD.n736 VDD.n22 8.45089
R2783 VDD.n738 VDD.n737 8.45089
R2784 VDD.n630 VDD.n86 8.45089
R2785 VDD.n629 VDD.n628 8.45089
R2786 VDD.n615 VDD.n88 8.45089
R2787 VDD.n616 VDD.n94 8.45089
R2788 VDD.n618 VDD.n617 8.45089
R2789 VDD.n614 VDD.n93 8.45089
R2790 VDD.n613 VDD.n612 8.45089
R2791 VDD.n602 VDD.n95 8.45089
R2792 VDD.n604 VDD.n603 8.45089
R2793 VDD.n601 VDD.n101 8.45089
R2794 VDD.n600 VDD.n599 8.45089
R2795 VDD.n103 VDD.n102 8.45089
R2796 VDD.n589 VDD.n108 8.45089
R2797 VDD.n591 VDD.n590 8.45089
R2798 VDD.n588 VDD.n110 8.45089
R2799 VDD.n587 VDD.n586 8.45089
R2800 VDD.n577 VDD.n111 8.45089
R2801 VDD.n579 VDD.n578 8.45089
R2802 VDD.n576 VDD.n116 8.45089
R2803 VDD.n574 VDD.n573 8.45089
R2804 VDD.n575 VDD.n574 8.45089
R2805 VDD.n118 VDD.n117 8.45089
R2806 VDD.n549 VDD.t64 8.45089
R2807 VDD.n548 VDD.n122 8.45089
R2808 VDD.n547 VDD.n546 8.45089
R2809 VDD.n124 VDD.n123 8.45089
R2810 VDD.n540 VDD.n539 8.45089
R2811 VDD.n538 VDD.n129 8.45089
R2812 VDD.n537 VDD.n536 8.45089
R2813 VDD.n525 VDD.n130 8.45089
R2814 VDD.n527 VDD.n526 8.45089
R2815 VDD.n524 VDD.n134 8.45089
R2816 VDD.n523 VDD.n522 8.45089
R2817 VDD.n136 VDD.n135 8.45089
R2818 VDD.n514 VDD.n513 8.45089
R2819 VDD.n512 VDD.n140 8.45089
R2820 VDD.n511 VDD.n510 8.45089
R2821 VDD.n499 VDD.n141 8.45089
R2822 VDD.n501 VDD.n500 8.45089
R2823 VDD.n498 VDD.n145 8.45089
R2824 VDD.n497 VDD.n496 8.45089
R2825 VDD.n488 VDD.n146 8.45089
R2826 VDD.n490 VDD.n489 8.45089
R2827 VDD.n487 VDD.n151 8.45089
R2828 VDD.n485 VDD.n484 8.45089
R2829 VDD.n486 VDD.n485 8.45089
R2830 VDD.n153 VDD.n152 8.45089
R2831 VDD.n460 VDD.t679 8.45089
R2832 VDD.n459 VDD.n157 8.45089
R2833 VDD.n458 VDD.n457 8.45089
R2834 VDD.n159 VDD.n158 8.45089
R2835 VDD.n451 VDD.n450 8.45089
R2836 VDD.n449 VDD.n164 8.45089
R2837 VDD.n448 VDD.n447 8.45089
R2838 VDD.n436 VDD.n165 8.45089
R2839 VDD.n438 VDD.n437 8.45089
R2840 VDD.n435 VDD.n169 8.45089
R2841 VDD.n434 VDD.n433 8.45089
R2842 VDD.n171 VDD.n170 8.45089
R2843 VDD.n425 VDD.n424 8.45089
R2844 VDD.n423 VDD.n175 8.45089
R2845 VDD.n422 VDD.n421 8.45089
R2846 VDD.n410 VDD.n176 8.45089
R2847 VDD.n412 VDD.n411 8.45089
R2848 VDD.n409 VDD.n180 8.45089
R2849 VDD.n408 VDD.n407 8.45089
R2850 VDD.n399 VDD.n181 8.45089
R2851 VDD.n401 VDD.n400 8.45089
R2852 VDD.n398 VDD.n186 8.45089
R2853 VDD.n396 VDD.n395 8.45089
R2854 VDD.n397 VDD.n396 8.45089
R2855 VDD.n188 VDD.n187 8.45089
R2856 VDD.n371 VDD.t347 8.45089
R2857 VDD.n370 VDD.n192 8.45089
R2858 VDD.n369 VDD.n368 8.45089
R2859 VDD.n194 VDD.n193 8.45089
R2860 VDD.n362 VDD.n361 8.45089
R2861 VDD.n360 VDD.n199 8.45089
R2862 VDD.n359 VDD.n358 8.45089
R2863 VDD.n347 VDD.n200 8.45089
R2864 VDD.n349 VDD.n348 8.45089
R2865 VDD.n346 VDD.n204 8.45089
R2866 VDD.n345 VDD.n344 8.45089
R2867 VDD.n206 VDD.n205 8.45089
R2868 VDD.n336 VDD.n335 8.45089
R2869 VDD.n334 VDD.n210 8.45089
R2870 VDD.n333 VDD.n332 8.45089
R2871 VDD.n321 VDD.n211 8.45089
R2872 VDD.n323 VDD.n322 8.45089
R2873 VDD.n320 VDD.n215 8.45089
R2874 VDD.n319 VDD.n318 8.45089
R2875 VDD.n310 VDD.n216 8.45089
R2876 VDD.n312 VDD.n311 8.45089
R2877 VDD.n309 VDD.n221 8.45089
R2878 VDD.n307 VDD.n306 8.45089
R2879 VDD.n308 VDD.n307 8.45089
R2880 VDD.n223 VDD.n222 8.45089
R2881 VDD.n282 VDD.t0 8.45089
R2882 VDD.n281 VDD.n227 8.45089
R2883 VDD.n280 VDD.n279 8.45089
R2884 VDD.n229 VDD.n228 8.45089
R2885 VDD.n273 VDD.n272 8.45089
R2886 VDD.n271 VDD.n234 8.45089
R2887 VDD.n270 VDD.n269 8.45089
R2888 VDD.n258 VDD.n235 8.45089
R2889 VDD.n260 VDD.n259 8.45089
R2890 VDD.n257 VDD.n239 8.45089
R2891 VDD.n256 VDD.n255 8.45089
R2892 VDD.n241 VDD.n240 8.45089
R2893 VDD.n245 VDD.n244 8.45089
R2894 VDD.n247 VDD.n246 8.45089
R2895 VDD.n2178 VDD.n2177 8.45089
R2896 VDD.n2179 VDD.n2178 8.45089
R2897 VDD.n2181 VDD.n2180 8.45089
R2898 VDD.n2186 VDD.n2185 8.45089
R2899 VDD.n2190 VDD.n2189 8.45089
R2900 VDD.n2195 VDD.n2194 8.45089
R2901 VDD.n2199 VDD.n2198 8.45089
R2902 VDD.n2203 VDD.n2202 8.45089
R2903 VDD.n2208 VDD.n2207 8.45089
R2904 VDD.n2213 VDD.n2212 8.45089
R2905 VDD.n2217 VDD.n2216 8.45089
R2906 VDD.n2223 VDD.n2222 8.45089
R2907 VDD.n2227 VDD.n2226 8.45089
R2908 VDD.n2231 VDD.n2230 8.45089
R2909 VDD.n2234 VDD.t509 8.45089
R2910 VDD.n2238 VDD.n2237 8.45089
R2911 VDD.n2242 VDD.n2241 8.45089
R2912 VDD.n2247 VDD.n2246 8.45089
R2913 VDD.n2252 VDD.n2251 8.45089
R2914 VDD.n2256 VDD.n2255 8.45089
R2915 VDD.n2260 VDD.n2259 8.45089
R2916 VDD.n2278 VDD.n2277 8.45089
R2917 VDD.n2277 VDD.n2276 8.45089
R2918 VDD.n2281 VDD.n2280 8.45089
R2919 VDD.n2286 VDD.n2285 8.45089
R2920 VDD.n11 VDD.n10 8.45089
R2921 VDD.n2294 VDD.n2293 8.45089
R2922 VDD.n2296 VDD.n2295 8.45089
R2923 VDD.n2313 VDD.n2312 8.45089
R2924 VDD.n2318 VDD.n2317 8.45089
R2925 VDD.n2322 VDD.n2321 8.45089
R2926 VDD.n2326 VDD.n2325 8.45089
R2927 VDD.n2352 VDD.n2351 8.45089
R2928 VDD.n2351 VDD.n2350 8.45089
R2929 VDD.n2357 VDD.n2356 8.45089
R2930 VDD.n2361 VDD.n2360 8.45089
R2931 VDD.n2365 VDD.n2364 8.45089
R2932 VDD.n2368 VDD.t303 8.45089
R2933 VDD.n2372 VDD.n2371 8.45089
R2934 VDD.n2376 VDD.n2375 8.45089
R2935 VDD.n2381 VDD.n2380 8.45089
R2936 VDD.n2386 VDD.n2385 8.45089
R2937 VDD.n2390 VDD.n2389 8.45089
R2938 VDD.n2394 VDD.n2393 8.45089
R2939 VDD.n2399 VDD.n2398 8.45089
R2940 VDD.n2403 VDD.n2402 8.45089
R2941 VDD.n2409 VDD.n2408 8.45089
R2942 VDD.n2413 VDD.n2412 8.45089
R2943 VDD.n2418 VDD.n2417 8.45089
R2944 VDD.n7 VDD.n6 8.45089
R2945 VDD.n2426 VDD.n2425 8.45089
R2946 VDD.n2428 VDD.n2427 8.45089
R2947 VDD.n2433 VDD.n2432 8.45089
R2948 VDD.n2437 VDD.n2436 8.45089
R2949 VDD.n2442 VDD.n2441 8.45089
R2950 VDD.n2446 VDD.n2445 8.45089
R2951 VDD.n2450 VDD.n2449 8.45089
R2952 VDD.n2476 VDD.n2475 8.45089
R2953 VDD.n2475 VDD.n2474 8.45089
R2954 VDD.n2481 VDD.n2480 8.45089
R2955 VDD.n2485 VDD.n2484 8.45089
R2956 VDD.n2489 VDD.n2488 8.45089
R2957 VDD.n2492 VDD.t738 8.45089
R2958 VDD.n2496 VDD.n2495 8.45089
R2959 VDD.n2500 VDD.n2499 8.45089
R2960 VDD.n2505 VDD.n2504 8.45089
R2961 VDD.n2510 VDD.n2509 8.45089
R2962 VDD.n2514 VDD.n2513 8.45089
R2963 VDD.n2518 VDD.n2517 8.45089
R2964 VDD.n2523 VDD.n2522 8.45089
R2965 VDD.n2527 VDD.n2526 8.45089
R2966 VDD.n2533 VDD.n2532 8.45089
R2967 VDD.n2537 VDD.n2536 8.45089
R2968 VDD.n2542 VDD.n2541 8.45089
R2969 VDD.n3 VDD.n2 8.45089
R2970 VDD.n2550 VDD.n2549 8.45089
R2971 VDD.n2552 VDD.n2551 8.45089
R2972 VDD.n2557 VDD.n2556 8.45089
R2973 VDD.n2561 VDD.n2560 8.45089
R2974 VDD.n2566 VDD.n2565 8.45089
R2975 VDD.n2570 VDD.n2569 8.45089
R2976 VDD.n2574 VDD.n2573 8.45089
R2977 VDD.n2600 VDD.n2599 8.45089
R2978 VDD.n2599 VDD.n2598 8.45089
R2979 VDD.n2605 VDD.n2604 8.45089
R2980 VDD.n2609 VDD.n2608 8.45089
R2981 VDD.n2613 VDD.n2612 8.45089
R2982 VDD.n2616 VDD.t706 8.45089
R2983 VDD.n2620 VDD.n2619 8.45089
R2984 VDD.n2624 VDD.n2623 8.45089
R2985 VDD.n2629 VDD.n2628 8.45089
R2986 VDD.n2634 VDD.n2633 8.45089
R2987 VDD.n2638 VDD.n2637 8.45089
R2988 VDD.n2642 VDD.n2641 8.45089
R2989 VDD.n2647 VDD.n2646 8.45089
R2990 VDD.n2651 VDD.n2650 8.45089
R2991 VDD.n2657 VDD.n2656 8.45089
R2992 VDD.n2661 VDD.n2660 8.45089
R2993 VDD.n2666 VDD.n2665 8.45089
R2994 VDD.n2797 VDD.n2796 8.45089
R2995 VDD.n2795 VDD.n2794 8.45089
R2996 VDD.n2793 VDD.n2792 8.45089
R2997 VDD.n2784 VDD.n2783 8.45089
R2998 VDD.n2779 VDD.n2778 8.45089
R2999 VDD.n2775 VDD.n2774 8.45089
R3000 VDD.n2771 VDD.n2770 8.45089
R3001 VDD.n2767 VDD.n2766 8.45089
R3002 VDD.n2743 VDD.n2742 8.45089
R3003 VDD.n2742 VDD.n2741 8.45089
R3004 VDD.n2738 VDD.n2737 8.45089
R3005 VDD.n2732 VDD.n2731 8.45089
R3006 VDD.n2728 VDD.n2727 8.45089
R3007 VDD.n2724 VDD.t287 8.45089
R3008 VDD.n2721 VDD.n2720 8.45089
R3009 VDD.n2717 VDD.n2716 8.45089
R3010 VDD.n2712 VDD.n2711 8.45089
R3011 VDD.n2707 VDD.n2706 8.45089
R3012 VDD.n2703 VDD.n2702 8.45089
R3013 VDD.n2698 VDD.n2697 8.45089
R3014 VDD.n2694 VDD.n2693 8.45089
R3015 VDD.n2688 VDD.n2687 8.45089
R3016 VDD.n2684 VDD.n2683 8.45089
R3017 VDD.n2680 VDD.n2679 8.45089
R3018 VDD.n2675 VDD.n2674 8.45089
R3019 VDD.n2672 VDD.n2671 8.45089
R3020 VDD.n2163 VDD.n2054 8.45089
R3021 VDD.n2162 VDD.n2161 8.45089
R3022 VDD.n2154 VDD.n2058 8.45089
R3023 VDD.n2064 VDD.n2063 8.45089
R3024 VDD.n2142 VDD.n2141 8.45089
R3025 VDD.n2066 VDD.n2065 8.45089
R3026 VDD.n2137 VDD.n2136 8.45089
R3027 VDD.n2075 VDD.n2072 8.45089
R3028 VDD.n2131 VDD.n2130 8.45089
R3029 VDD.n2074 VDD.n2073 8.45089
R3030 VDD.n2126 VDD.n2125 8.45089
R3031 VDD.n2120 VDD.n2119 8.45089
R3032 VDD.n2081 VDD.n2080 8.45089
R3033 VDD.n2115 VDD.n2114 8.45089
R3034 VDD.n2084 VDD.n2083 8.45089
R3035 VDD.n2109 VDD.n2108 8.45089
R3036 VDD.n2086 VDD.n2085 8.45089
R3037 VDD.n2104 VDD.n2103 8.45089
R3038 VDD.n2091 VDD.n2090 8.45089
R3039 VDD.n2093 VDD.n2092 8.45089
R3040 VDD.n2038 VDD.n2037 8.45089
R3041 VDD.n1469 VDD.n1468 8.45089
R3042 VDD.n2033 VDD.n2032 8.45089
R3043 VDD.n1476 VDD.n1473 8.45089
R3044 VDD.n2028 VDD.n2027 8.45089
R3045 VDD.n2024 VDD.n1474 8.45089
R3046 VDD.n2023 VDD.n2022 8.45089
R3047 VDD.n2017 VDD.n2016 8.45089
R3048 VDD.n1482 VDD.n1481 8.45089
R3049 VDD.n2009 VDD.n2008 8.45089
R3050 VDD.n1485 VDD.n1484 8.45089
R3051 VDD.n2005 VDD.n2004 8.45089
R3052 VDD.n2001 VDD.n1487 8.45089
R3053 VDD.n2000 VDD.n1999 8.45089
R3054 VDD.n1492 VDD.n1491 8.45089
R3055 VDD.n1494 VDD.n1493 8.45089
R3056 VDD.n1987 VDD.n1986 8.45089
R3057 VDD.n1497 VDD.n1496 8.45089
R3058 VDD.n1500 VDD.n1499 8.45089
R3059 VDD.n1503 VDD.n1502 8.45089
R3060 VDD.n1969 VDD.n1968 8.45089
R3061 VDD.n1961 VDD.n1960 8.45089
R3062 VDD.n1508 VDD.n1507 8.45089
R3063 VDD.n1955 VDD.n1954 8.45089
R3064 VDD.n1951 VDD.n1509 8.45089
R3065 VDD.n1950 VDD.n1949 8.45089
R3066 VDD.n1517 VDD.n1514 8.45089
R3067 VDD.n1944 VDD.n1943 8.45089
R3068 VDD.n1936 VDD.n1935 8.45089
R3069 VDD.n1520 VDD.n1519 8.45089
R3070 VDD.n1931 VDD.n1930 8.45089
R3071 VDD.n1523 VDD.n1522 8.45089
R3072 VDD.n1926 VDD.n1925 8.45089
R3073 VDD.n1531 VDD.n1527 8.45089
R3074 VDD.n1921 VDD.n1920 8.45089
R3075 VDD.n1530 VDD.n1529 8.45089
R3076 VDD.n1535 VDD.n1534 8.45089
R3077 VDD.n1910 VDD.n1909 8.45089
R3078 VDD.n1537 VDD.n1536 8.45089
R3079 VDD.n1540 VDD.n1539 8.45089
R3080 VDD.n1542 VDD.n1541 8.45089
R3081 VDD.n1891 VDD.n1890 8.45089
R3082 VDD.n1885 VDD.n1884 8.45089
R3083 VDD.n1550 VDD.n1549 8.45089
R3084 VDD.n1880 VDD.n1879 8.45089
R3085 VDD.n1557 VDD.n1554 8.45089
R3086 VDD.n1875 VDD.n1874 8.45089
R3087 VDD.n1871 VDD.n1555 8.45089
R3088 VDD.n1870 VDD.n1869 8.45089
R3089 VDD.n1864 VDD.n1863 8.45089
R3090 VDD.n1563 VDD.n1562 8.45089
R3091 VDD.n1856 VDD.n1855 8.45089
R3092 VDD.n1566 VDD.n1565 8.45089
R3093 VDD.n1852 VDD.n1851 8.45089
R3094 VDD.n1848 VDD.n1568 8.45089
R3095 VDD.n1847 VDD.n1846 8.45089
R3096 VDD.n1573 VDD.n1572 8.45089
R3097 VDD.n1575 VDD.n1574 8.45089
R3098 VDD.n1834 VDD.n1833 8.45089
R3099 VDD.n1578 VDD.n1577 8.45089
R3100 VDD.n1581 VDD.n1580 8.45089
R3101 VDD.n1584 VDD.n1583 8.45089
R3102 VDD.n1816 VDD.n1815 8.45089
R3103 VDD.n1808 VDD.n1807 8.45089
R3104 VDD.n1589 VDD.n1588 8.45089
R3105 VDD.n1802 VDD.n1801 8.45089
R3106 VDD.n1798 VDD.n1590 8.45089
R3107 VDD.n1797 VDD.n1796 8.45089
R3108 VDD.n1598 VDD.n1595 8.45089
R3109 VDD.n1791 VDD.n1790 8.45089
R3110 VDD.n1783 VDD.n1782 8.45089
R3111 VDD.n1601 VDD.n1600 8.45089
R3112 VDD.n1778 VDD.n1777 8.45089
R3113 VDD.n1604 VDD.n1603 8.45089
R3114 VDD.n1773 VDD.n1772 8.45089
R3115 VDD.n1612 VDD.n1608 8.45089
R3116 VDD.n1768 VDD.n1767 8.45089
R3117 VDD.n1611 VDD.n1610 8.45089
R3118 VDD.n1616 VDD.n1615 8.45089
R3119 VDD.n1757 VDD.n1756 8.45089
R3120 VDD.n1618 VDD.n1617 8.45089
R3121 VDD.n1621 VDD.n1620 8.45089
R3122 VDD.n1623 VDD.n1622 8.45089
R3123 VDD.n1738 VDD.n1737 8.45089
R3124 VDD.n1732 VDD.n1731 8.45089
R3125 VDD.n1631 VDD.n1630 8.45089
R3126 VDD.n1727 VDD.n1726 8.45089
R3127 VDD.n1638 VDD.n1635 8.45089
R3128 VDD.n1722 VDD.n1721 8.45089
R3129 VDD.n1718 VDD.n1636 8.45089
R3130 VDD.n1717 VDD.n1716 8.45089
R3131 VDD.n1711 VDD.n1710 8.45089
R3132 VDD.n1644 VDD.n1643 8.45089
R3133 VDD.n1703 VDD.n1702 8.45089
R3134 VDD.n1647 VDD.n1646 8.45089
R3135 VDD.n1699 VDD.n1698 8.45089
R3136 VDD.n1695 VDD.n1649 8.45089
R3137 VDD.n1694 VDD.n1693 8.45089
R3138 VDD.n1654 VDD.n1653 8.45089
R3139 VDD.n1656 VDD.n1655 8.45089
R3140 VDD.n1681 VDD.n1680 8.45089
R3141 VDD.n1659 VDD.n1658 8.45089
R3142 VDD.n1662 VDD.n1661 8.45089
R3143 VDD.n828 VDD.n825 8.45089
R3144 VDD.n1454 VDD.n1453 8.45089
R3145 VDD.n1301 VDD.n1300 8.45089
R3146 VDD.n909 VDD.n908 8.45089
R3147 VDD.n1291 VDD.n1290 8.45089
R3148 VDD.n913 VDD.n912 8.45089
R3149 VDD.n1286 VDD.n1283 8.45089
R3150 VDD.n917 VDD.n916 8.45089
R3151 VDD.n1279 VDD.n1278 8.45089
R3152 VDD.n1272 VDD.n1271 8.45089
R3153 VDD.n921 VDD.n920 8.45089
R3154 VDD.n923 VDD.n922 8.45089
R3155 VDD.n926 VDD.n925 8.45089
R3156 VDD.n1251 VDD.n1250 8.45089
R3157 VDD.n928 VDD.n927 8.45089
R3158 VDD.n932 VDD.n931 8.45089
R3159 VDD.n1239 VDD.n1238 8.45089
R3160 VDD.n934 VDD.n933 8.45089
R3161 VDD.n1234 VDD.n1231 8.45089
R3162 VDD.n937 VDD.n936 8.45089
R3163 VDD.n1227 VDD.n1226 8.45089
R3164 VDD.n939 VDD.n938 8.45089
R3165 VDD.n1222 VDD.n1221 8.45089
R3166 VDD.n1216 VDD.n1215 8.45089
R3167 VDD.n946 VDD.n945 8.45089
R3168 VDD.n1211 VDD.n1209 8.45089
R3169 VDD.n949 VDD.n948 8.45089
R3170 VDD.n1204 VDD.n1203 8.45089
R3171 VDD.n951 VDD.n950 8.45089
R3172 VDD.n1199 VDD.n1198 8.45089
R3173 VDD.n1193 VDD.n1192 8.45089
R3174 VDD.n960 VDD.n959 8.45089
R3175 VDD.n964 VDD.n963 8.45089
R3176 VDD.n966 VDD.n965 8.45089
R3177 VDD.n1175 VDD.n1174 8.45089
R3178 VDD.n969 VDD.n968 8.45089
R3179 VDD.n971 VDD.n970 8.45089
R3180 VDD.n1162 VDD.n1161 8.45089
R3181 VDD.n974 VDD.n973 8.45089
R3182 VDD.n1156 VDD.n1155 8.45089
R3183 VDD.n976 VDD.n975 8.45089
R3184 VDD.n1151 VDD.n1150 8.45089
R3185 VDD.n981 VDD.n980 8.45089
R3186 VDD.n1146 VDD.n1145 8.45089
R3187 VDD.n1139 VDD.n1138 8.45089
R3188 VDD.n986 VDD.n985 8.45089
R3189 VDD.n1133 VDD.n1132 8.45089
R3190 VDD.n989 VDD.n988 8.45089
R3191 VDD.n1128 VDD.n1125 8.45089
R3192 VDD.n993 VDD.n992 8.45089
R3193 VDD.n1121 VDD.n1120 8.45089
R3194 VDD.n1114 VDD.n1113 8.45089
R3195 VDD.n997 VDD.n996 8.45089
R3196 VDD.n999 VDD.n998 8.45089
R3197 VDD.n1002 VDD.n1001 8.45089
R3198 VDD.n1093 VDD.n1092 8.45089
R3199 VDD.n1004 VDD.n1003 8.45089
R3200 VDD.n1008 VDD.n1007 8.45089
R3201 VDD.n1081 VDD.n1080 8.45089
R3202 VDD.n1010 VDD.n1009 8.45089
R3203 VDD.n1076 VDD.n1073 8.45089
R3204 VDD.n1013 VDD.n1012 8.45089
R3205 VDD.n1069 VDD.n1068 8.45089
R3206 VDD.n1015 VDD.n1014 8.45089
R3207 VDD.n1064 VDD.n1063 8.45089
R3208 VDD.n1058 VDD.n1057 8.45089
R3209 VDD.n1022 VDD.n1021 8.45089
R3210 VDD.n1053 VDD.n1051 8.45089
R3211 VDD.n1025 VDD.n1024 8.45089
R3212 VDD.n1046 VDD.n1045 8.45089
R3213 VDD.n1027 VDD.n1026 8.45089
R3214 VDD.n1041 VDD.n1040 8.45089
R3215 VDD.n758 VDD.n757 8.45089
R3216 VDD.n754 VDD.n17 8.45089
R3217 VDD.n753 VDD.n752 8.45089
R3218 VDD.n745 VDD.n21 8.45089
R3219 VDD.n23 VDD.n22 8.45089
R3220 VDD.n740 VDD.n738 8.45089
R3221 VDD.n636 VDD.n86 8.45089
R3222 VDD.n628 VDD.n627 8.45089
R3223 VDD.n625 VDD.n88 8.45089
R3224 VDD.n94 VDD.n90 8.45089
R3225 VDD.n621 VDD.n618 8.45089
R3226 VDD.n93 VDD.n92 8.45089
R3227 VDD.n612 VDD.n611 8.45089
R3228 VDD.n96 VDD.n95 8.45089
R3229 VDD.n607 VDD.n604 8.45089
R3230 VDD.n101 VDD.n100 8.45089
R3231 VDD.n599 VDD.n598 8.45089
R3232 VDD.n104 VDD.n103 8.45089
R3233 VDD.n592 VDD.n591 8.45089
R3234 VDD.n110 VDD.n109 8.45089
R3235 VDD.n586 VDD.n585 8.45089
R3236 VDD.n581 VDD.n111 8.45089
R3237 VDD.n580 VDD.n579 8.45089
R3238 VDD.n567 VDD.n116 8.45089
R3239 VDD.n119 VDD.n118 8.45089
R3240 VDD.n550 VDD.n549 8.45089
R3241 VDD.n122 VDD.n121 8.45089
R3242 VDD.n546 VDD.n545 8.45089
R3243 VDD.n542 VDD.n124 8.45089
R3244 VDD.n541 VDD.n540 8.45089
R3245 VDD.n129 VDD.n128 8.45089
R3246 VDD.n131 VDD.n130 8.45089
R3247 VDD.n528 VDD.n527 8.45089
R3248 VDD.n134 VDD.n133 8.45089
R3249 VDD.n137 VDD.n136 8.45089
R3250 VDD.n140 VDD.n139 8.45089
R3251 VDD.n510 VDD.n509 8.45089
R3252 VDD.n502 VDD.n501 8.45089
R3253 VDD.n145 VDD.n144 8.45089
R3254 VDD.n496 VDD.n495 8.45089
R3255 VDD.n492 VDD.n146 8.45089
R3256 VDD.n491 VDD.n490 8.45089
R3257 VDD.n478 VDD.n151 8.45089
R3258 VDD.n154 VDD.n153 8.45089
R3259 VDD.n461 VDD.n460 8.45089
R3260 VDD.n157 VDD.n156 8.45089
R3261 VDD.n457 VDD.n456 8.45089
R3262 VDD.n453 VDD.n159 8.45089
R3263 VDD.n452 VDD.n451 8.45089
R3264 VDD.n164 VDD.n163 8.45089
R3265 VDD.n166 VDD.n165 8.45089
R3266 VDD.n439 VDD.n438 8.45089
R3267 VDD.n169 VDD.n168 8.45089
R3268 VDD.n172 VDD.n171 8.45089
R3269 VDD.n175 VDD.n174 8.45089
R3270 VDD.n421 VDD.n420 8.45089
R3271 VDD.n413 VDD.n412 8.45089
R3272 VDD.n180 VDD.n179 8.45089
R3273 VDD.n407 VDD.n406 8.45089
R3274 VDD.n403 VDD.n181 8.45089
R3275 VDD.n402 VDD.n401 8.45089
R3276 VDD.n389 VDD.n186 8.45089
R3277 VDD.n189 VDD.n188 8.45089
R3278 VDD.n372 VDD.n371 8.45089
R3279 VDD.n192 VDD.n191 8.45089
R3280 VDD.n368 VDD.n367 8.45089
R3281 VDD.n364 VDD.n194 8.45089
R3282 VDD.n363 VDD.n362 8.45089
R3283 VDD.n199 VDD.n198 8.45089
R3284 VDD.n201 VDD.n200 8.45089
R3285 VDD.n350 VDD.n349 8.45089
R3286 VDD.n204 VDD.n203 8.45089
R3287 VDD.n207 VDD.n206 8.45089
R3288 VDD.n210 VDD.n209 8.45089
R3289 VDD.n332 VDD.n331 8.45089
R3290 VDD.n324 VDD.n323 8.45089
R3291 VDD.n215 VDD.n214 8.45089
R3292 VDD.n318 VDD.n317 8.45089
R3293 VDD.n314 VDD.n216 8.45089
R3294 VDD.n313 VDD.n312 8.45089
R3295 VDD.n300 VDD.n221 8.45089
R3296 VDD.n224 VDD.n223 8.45089
R3297 VDD.n283 VDD.n282 8.45089
R3298 VDD.n227 VDD.n226 8.45089
R3299 VDD.n279 VDD.n278 8.45089
R3300 VDD.n275 VDD.n229 8.45089
R3301 VDD.n274 VDD.n273 8.45089
R3302 VDD.n234 VDD.n233 8.45089
R3303 VDD.n236 VDD.n235 8.45089
R3304 VDD.n261 VDD.n260 8.45089
R3305 VDD.n239 VDD.n238 8.45089
R3306 VDD.n242 VDD.n241 8.45089
R3307 VDD.n2187 VDD.n2186 8.45089
R3308 VDD.n2196 VDD.n2195 8.45089
R3309 VDD.n2200 VDD.n2199 8.45089
R3310 VDD.n2204 VDD.n2203 8.45089
R3311 VDD.n2214 VDD.n2213 8.45089
R3312 VDD.n2218 VDD.n2217 8.45089
R3313 VDD.n2224 VDD.n2223 8.45089
R3314 VDD.n2228 VDD.n2227 8.45089
R3315 VDD.n2232 VDD.n2231 8.45089
R3316 VDD.n2235 VDD.n2234 8.45089
R3317 VDD.n2239 VDD.n2238 8.45089
R3318 VDD.n2243 VDD.n2242 8.45089
R3319 VDD.n2253 VDD.n2252 8.45089
R3320 VDD.n2257 VDD.n2256 8.45089
R3321 VDD.n2262 VDD.n2260 8.45089
R3322 VDD.n2282 VDD.n2281 8.45089
R3323 VDD.n2291 VDD.n11 8.45089
R3324 VDD.n2293 VDD.n2292 8.45089
R3325 VDD.n2319 VDD.n2318 8.45089
R3326 VDD.n2323 VDD.n2322 8.45089
R3327 VDD.n2327 VDD.n2326 8.45089
R3328 VDD.n2358 VDD.n2357 8.45089
R3329 VDD.n2362 VDD.n2361 8.45089
R3330 VDD.n2366 VDD.n2365 8.45089
R3331 VDD.n2369 VDD.n2368 8.45089
R3332 VDD.n2373 VDD.n2372 8.45089
R3333 VDD.n2377 VDD.n2376 8.45089
R3334 VDD.n2387 VDD.n2386 8.45089
R3335 VDD.n2391 VDD.n2390 8.45089
R3336 VDD.n2396 VDD.n2394 8.45089
R3337 VDD.n2400 VDD.n2399 8.45089
R3338 VDD.n2406 VDD.n2403 8.45089
R3339 VDD.n2410 VDD.n2409 8.45089
R3340 VDD.n2414 VDD.n2413 8.45089
R3341 VDD.n2423 VDD.n7 8.45089
R3342 VDD.n2425 VDD.n2424 8.45089
R3343 VDD.n2434 VDD.n2433 8.45089
R3344 VDD.n2443 VDD.n2442 8.45089
R3345 VDD.n2447 VDD.n2446 8.45089
R3346 VDD.n2451 VDD.n2450 8.45089
R3347 VDD.n2482 VDD.n2481 8.45089
R3348 VDD.n2486 VDD.n2485 8.45089
R3349 VDD.n2490 VDD.n2489 8.45089
R3350 VDD.n2493 VDD.n2492 8.45089
R3351 VDD.n2497 VDD.n2496 8.45089
R3352 VDD.n2501 VDD.n2500 8.45089
R3353 VDD.n2511 VDD.n2510 8.45089
R3354 VDD.n2515 VDD.n2514 8.45089
R3355 VDD.n2520 VDD.n2518 8.45089
R3356 VDD.n2524 VDD.n2523 8.45089
R3357 VDD.n2530 VDD.n2527 8.45089
R3358 VDD.n2534 VDD.n2533 8.45089
R3359 VDD.n2538 VDD.n2537 8.45089
R3360 VDD.n2547 VDD.n3 8.45089
R3361 VDD.n2549 VDD.n2548 8.45089
R3362 VDD.n2558 VDD.n2557 8.45089
R3363 VDD.n2567 VDD.n2566 8.45089
R3364 VDD.n2571 VDD.n2570 8.45089
R3365 VDD.n2575 VDD.n2574 8.45089
R3366 VDD.n2606 VDD.n2605 8.45089
R3367 VDD.n2610 VDD.n2609 8.45089
R3368 VDD.n2614 VDD.n2613 8.45089
R3369 VDD.n2617 VDD.n2616 8.45089
R3370 VDD.n2621 VDD.n2620 8.45089
R3371 VDD.n2625 VDD.n2624 8.45089
R3372 VDD.n2635 VDD.n2634 8.45089
R3373 VDD.n2639 VDD.n2638 8.45089
R3374 VDD.n2644 VDD.n2642 8.45089
R3375 VDD.n2648 VDD.n2647 8.45089
R3376 VDD.n2654 VDD.n2651 8.45089
R3377 VDD.n2658 VDD.n2657 8.45089
R3378 VDD.n2662 VDD.n2661 8.45089
R3379 VDD.n2798 VDD.n2797 8.45089
R3380 VDD.n2794 VDD.n2670 8.45089
R3381 VDD.n2785 VDD.n2784 8.45089
R3382 VDD.n2776 VDD.n2775 8.45089
R3383 VDD.n2772 VDD.n2771 8.45089
R3384 VDD.n2768 VDD.n2767 8.45089
R3385 VDD.n2739 VDD.n2738 8.45089
R3386 VDD.n2733 VDD.n2732 8.45089
R3387 VDD.n2729 VDD.n2728 8.45089
R3388 VDD.n2725 VDD.n2724 8.45089
R3389 VDD.n2722 VDD.n2721 8.45089
R3390 VDD.n2718 VDD.n2717 8.45089
R3391 VDD.n2708 VDD.n2707 8.45089
R3392 VDD.n2704 VDD.n2703 8.45089
R3393 VDD.n2700 VDD.n2698 8.45089
R3394 VDD.n2695 VDD.n2694 8.45089
R3395 VDD.n2691 VDD.n2688 8.45089
R3396 VDD.n2685 VDD.n2684 8.45089
R3397 VDD.n2681 VDD.n2680 8.45089
R3398 VDD.n1638 VDD.n1634 8.31095
R3399 VDD.n1798 VDD.n1592 8.31095
R3400 VDD.n1557 VDD.n1553 8.31095
R3401 VDD.n1951 VDD.n1511 8.31095
R3402 VDD.n1476 VDD.n1472 8.31095
R3403 VDD.n1029 VDD.n1024 8.31095
R3404 VDD.n1127 VDD.n989 8.31095
R3405 VDD.n953 VDD.n948 8.31095
R3406 VDD.n1285 VDD.n913 8.31095
R3407 VDD.n581 VDD.n113 8.31095
R3408 VDD.n492 VDD.n148 8.31095
R3409 VDD.n403 VDD.n183 8.31095
R3410 VDD.n314 VDD.n218 8.31095
R3411 VDD.n2108 VDD.n2088 8.16602
R3412 VDD.n2126 VDD.n2078 8.16602
R3413 VDD.n2748 VDD.n2747 8.00414
R3414 VDD.n2584 VDD.n2583 8.00414
R3415 VDD.n2460 VDD.n2459 8.00414
R3416 VDD.n2336 VDD.n2335 8.00414
R3417 VDD.n1692 VDD.t190 7.91717
R3418 VDD.t739 VDD.n1769 7.91717
R3419 VDD.n1845 VDD.t314 7.91717
R3420 VDD.t484 VDD.n1922 7.91717
R3421 VDD.n1998 VDD.t332 7.91717
R3422 VDD.n2741 VDD.t396 7.89524
R3423 VDD.n2598 VDD.t351 7.89524
R3424 VDD.n2474 VDD.t676 7.89524
R3425 VDD.n2350 VDD.t37 7.89524
R3426 VDD.n2216 VDD.t98 7.89524
R3427 VDD.n272 VDD.t524 7.80872
R3428 VDD.n361 VDD.t30 7.80872
R3429 VDD.n450 VDD.t97 7.80872
R3430 VDD.n539 VDD.t283 7.80872
R3431 VDD.n695 VDD.t572 7.80872
R3432 VDD.n1082 VDD.t68 7.74507
R3433 VDD.n1160 VDD.t11 7.74507
R3434 VDD.n1240 VDD.t666 7.74507
R3435 VDD.t62 VDD.n1456 7.74507
R3436 VDD.n678 VDD.n677 7.72464
R3437 VDD.n1355 VDD.n878 7.70756
R3438 VDD.n2756 VDD.n2755 6.95412
R3439 VDD.n2592 VDD.n2591 6.95412
R3440 VDD.n2468 VDD.n2467 6.95412
R3441 VDD.n2344 VDD.n2343 6.95412
R3442 VDD.n1424 VDD.n840 6.84188
R3443 VDD.n1439 VDD.n830 6.84188
R3444 VDD.n606 VDD.n96 6.62119
R3445 VDD.n621 VDD.n620 6.62119
R3446 VDD.n787 VDD.n784 6.4005
R3447 VDD.n1440 VDD.n1439 6.33153
R3448 VDD.n1424 VDD.n844 6.32841
R3449 VDD.n1306 VDD.n906 6.32433
R3450 VDD.n1387 VDD.n1386 6.32433
R3451 VDD.n739 VDD.n23 5.51774
R3452 VDD.n1688 VDD.n1653 5.29705
R3453 VDD.n1762 VDD.n1611 5.29705
R3454 VDD.n1841 VDD.n1572 5.29705
R3455 VDD.n1915 VDD.n1530 5.29705
R3456 VDD.n1994 VDD.n1491 5.29705
R3457 VDD.n1087 VDD.n1007 5.29705
R3458 VDD.n1168 VDD.n971 5.29705
R3459 VDD.n1245 VDD.n931 5.29705
R3460 VDD.n535 VDD.n128 5.29705
R3461 VDD.n446 VDD.n163 5.29705
R3462 VDD.n357 VDD.n198 5.29705
R3463 VDD.n268 VDD.n233 5.29705
R3464 VDD.n683 VDD.t574 5.20598
R3465 VDD.n679 VDD.n678 5.07636
R3466 VDD.n294 VDD 5.04292
R3467 VDD.n383 VDD 5.04292
R3468 VDD.n472 VDD 5.04292
R3469 VDD.n561 VDD 5.04292
R3470 VDD.n2150 VDD.n2149 5.02697
R3471 VDD.n2151 VDD.n2059 4.6505
R3472 VDD.n899 VDD.n898 4.6505
R3473 VDD.n1319 VDD.n897 4.6505
R3474 VDD.n1331 VDD.n889 4.6505
R3475 VDD.n1341 VDD.n884 4.6505
R3476 VDD.n1344 VDD.n883 4.6505
R3477 VDD.n1360 VDD.n875 4.6505
R3478 VDD.n1370 VDD.n870 4.6505
R3479 VDD.n1374 VDD.n869 4.6505
R3480 VDD.n1397 VDD.n857 4.6505
R3481 VDD.n1407 VDD.n852 4.6505
R3482 VDD.n1411 VDD.n851 4.6505
R3483 VDD.n1427 VDD.n841 4.6505
R3484 VDD.n1450 VDD.n1449 4.6505
R3485 VDD.n791 VDD.n783 4.6505
R3486 VDD.n822 VDD.n821 4.6505
R3487 VDD.n798 VDD.n797 4.6505
R3488 VDD.n807 VDD.n775 4.6505
R3489 VDD.n809 VDD.n808 4.6505
R3490 VDD.n815 VDD.n814 4.6505
R3491 VDD.n788 VDD.n787 4.6505
R3492 VDD.n304 VDD.n303 4.6505
R3493 VDD.n302 VDD.n301 4.6505
R3494 VDD.n393 VDD.n392 4.6505
R3495 VDD.n391 VDD.n390 4.6505
R3496 VDD.n482 VDD.n481 4.6505
R3497 VDD.n480 VDD.n479 4.6505
R3498 VDD.n571 VDD.n570 4.6505
R3499 VDD.n569 VDD.n568 4.6505
R3500 VDD.n648 VDD.n76 4.6505
R3501 VDD.n70 VDD.n69 4.6505
R3502 VDD.n663 VDD.n68 4.6505
R3503 VDD.n675 VDD.n60 4.6505
R3504 VDD.n686 VDD.n54 4.6505
R3505 VDD.n48 VDD.n47 4.6505
R3506 VDD.n701 VDD.n46 4.6505
R3507 VDD.n713 VDD.n38 4.6505
R3508 VDD.n724 VDD.n32 4.6505
R3509 VDD.n729 VDD.n728 4.6505
R3510 VDD.n2760 VDD.n2759 4.6505
R3511 VDD.n2765 VDD.n2764 4.6505
R3512 VDD.n2596 VDD.n2595 4.6505
R3513 VDD.n2580 VDD.n2579 4.6505
R3514 VDD.n2472 VDD.n2471 4.6505
R3515 VDD.n2456 VDD.n2455 4.6505
R3516 VDD.n2348 VDD.n2347 4.6505
R3517 VDD.n2332 VDD.n2331 4.6505
R3518 VDD.n2275 VDD.n2274 4.6505
R3519 VDD.n2270 VDD.n2269 4.6505
R3520 VDD.n2748 VDD 4.55532
R3521 VDD.n2584 VDD 4.55532
R3522 VDD.n2460 VDD 4.55532
R3523 VDD.n2336 VDD 4.55532
R3524 VDD.n813 VDD.n774 4.5005
R3525 VDD.n793 VDD.n792 4.5005
R3526 VDD.n2753 VDD.n2752 4.46483
R3527 VDD.n2589 VDD.n2588 4.46483
R3528 VDD.n2465 VDD.n2464 4.46483
R3529 VDD.n2341 VDD.n2340 4.46483
R3530 VDD.n1305 VDD.n904 4.44959
R3531 VDD.n1385 VDD.n1384 4.44959
R3532 VDD.n1423 VDD.n842 4.43314
R3533 VDD.n1438 VDD.n1437 4.42059
R3534 VDD.n699 VDD.n698 4.1936
R3535 VDD.n635 VDD.n82 3.75222
R3536 VDD.n763 VDD 3.75222
R3537 VDD.n2310 VDD.n2309 3.75222
R3538 VDD.n2163 VDD 3.53153
R3539 VDD.n1698 VDD.n1651 3.53153
R3540 VDD.n1773 VDD.n1607 3.53153
R3541 VDD.n1851 VDD.n1570 3.53153
R3542 VDD.n1926 VDD.n1526 3.53153
R3543 VDD.n2004 VDD.n1489 3.53153
R3544 VDD.n1076 VDD.n1075 3.53153
R3545 VDD.n1155 VDD.n978 3.53153
R3546 VDD.n1234 VDD.n1233 3.53153
R3547 VDD.n1386 VDD.n863 3.53153
R3548 VDD.n754 VDD 3.53153
R3549 VDD.n545 VDD.n126 3.53153
R3550 VDD.n456 VDD.n161 3.53153
R3551 VDD.n367 VDD.n196 3.53153
R3552 VDD.n278 VDD.n231 3.53153
R3553 VDD.n2302 VDD.n2301 3.53153
R3554 VDD.n2308 VDD.n2304 3.52991
R3555 VDD.n1035 VDD.n1030 3.22029
R3556 VDD.n2678 VDD.n2672 3.22029
R3557 VDD.n800 VDD.n799 3.2005
R3558 VDD VDD.n2093 3.12394
R3559 VDD.n1667 VDD 3.12394
R3560 VDD.n247 VDD 3.12394
R3561 VDD.n289 VDD 3.10353
R3562 VDD.n378 VDD 3.10353
R3563 VDD.n467 VDD 3.10353
R3564 VDD.n556 VDD 3.10353
R3565 VDD.n2173 VDD.n2172 3.1005
R3566 VDD.n2166 VDD.n2165 3.1005
R3567 VDD.n2148 VDD.n2147 3.1005
R3568 VDD.n2090 VDD.n2089 3.1005
R3569 VDD.n2105 VDD.n2104 3.1005
R3570 VDD.n2106 VDD.n2086 3.1005
R3571 VDD.n2108 VDD.n2107 3.1005
R3572 VDD.n2083 VDD.n2082 3.1005
R3573 VDD.n2116 VDD.n2115 3.1005
R3574 VDD.n2117 VDD.n2081 3.1005
R3575 VDD.n2119 VDD.n2118 3.1005
R3576 VDD.n2127 VDD.n2126 3.1005
R3577 VDD.n2128 VDD.n2074 3.1005
R3578 VDD.n2130 VDD.n2129 3.1005
R3579 VDD.n2075 VDD.n2069 3.1005
R3580 VDD.n2138 VDD.n2137 3.1005
R3581 VDD.n2139 VDD.n2066 3.1005
R3582 VDD.n2141 VDD.n2140 3.1005
R3583 VDD.n2063 VDD.n2062 3.1005
R3584 VDD.n2154 VDD.n2153 3.1005
R3585 VDD.n2162 VDD.n2055 3.1005
R3586 VDD.n2164 VDD.n2163 3.1005
R3587 VDD.n2043 VDD.n2042 3.1005
R3588 VDD.n1671 VDD.n1662 3.1005
R3589 VDD.n1658 VDD.n1657 3.1005
R3590 VDD.n1682 VDD.n1681 3.1005
R3591 VDD.n1683 VDD.n1656 3.1005
R3592 VDD.n1684 VDD.n1653 3.1005
R3593 VDD.n1694 VDD.n1652 3.1005
R3594 VDD.n1696 VDD.n1695 3.1005
R3595 VDD.n1698 VDD.n1697 3.1005
R3596 VDD.n1646 VDD.n1645 3.1005
R3597 VDD.n1704 VDD.n1703 3.1005
R3598 VDD.n1705 VDD.n1644 3.1005
R3599 VDD.n1710 VDD.n1709 3.1005
R3600 VDD.n1717 VDD.n1639 3.1005
R3601 VDD.n1719 VDD.n1718 3.1005
R3602 VDD.n1721 VDD.n1720 3.1005
R3603 VDD.n1638 VDD.n1632 3.1005
R3604 VDD.n1728 VDD.n1727 3.1005
R3605 VDD.n1729 VDD.n1631 3.1005
R3606 VDD.n1731 VDD.n1730 3.1005
R3607 VDD.n1739 VDD.n1738 3.1005
R3608 VDD.n1740 VDD.n1623 3.1005
R3609 VDD.n1620 VDD.n1619 3.1005
R3610 VDD.n1754 VDD.n1618 3.1005
R3611 VDD.n1756 VDD.n1755 3.1005
R3612 VDD.n1615 VDD.n1613 3.1005
R3613 VDD.n1765 VDD.n1611 3.1005
R3614 VDD.n1767 VDD.n1766 3.1005
R3615 VDD.n1612 VDD.n1605 3.1005
R3616 VDD.n1774 VDD.n1773 3.1005
R3617 VDD.n1775 VDD.n1604 3.1005
R3618 VDD.n1777 VDD.n1776 3.1005
R3619 VDD.n1600 VDD.n1599 3.1005
R3620 VDD.n1784 VDD.n1783 3.1005
R3621 VDD.n1790 VDD.n1789 3.1005
R3622 VDD.n1788 VDD.n1598 3.1005
R3623 VDD.n1797 VDD.n1593 3.1005
R3624 VDD.n1799 VDD.n1798 3.1005
R3625 VDD.n1801 VDD.n1800 3.1005
R3626 VDD.n1588 VDD.n1587 3.1005
R3627 VDD.n1809 VDD.n1808 3.1005
R3628 VDD.n1815 VDD.n1814 3.1005
R3629 VDD.n1813 VDD.n1583 3.1005
R3630 VDD.n1824 VDD.n1581 3.1005
R3631 VDD.n1577 VDD.n1576 3.1005
R3632 VDD.n1835 VDD.n1834 3.1005
R3633 VDD.n1836 VDD.n1575 3.1005
R3634 VDD.n1837 VDD.n1572 3.1005
R3635 VDD.n1847 VDD.n1571 3.1005
R3636 VDD.n1849 VDD.n1848 3.1005
R3637 VDD.n1851 VDD.n1850 3.1005
R3638 VDD.n1565 VDD.n1564 3.1005
R3639 VDD.n1857 VDD.n1856 3.1005
R3640 VDD.n1858 VDD.n1563 3.1005
R3641 VDD.n1863 VDD.n1862 3.1005
R3642 VDD.n1870 VDD.n1558 3.1005
R3643 VDD.n1872 VDD.n1871 3.1005
R3644 VDD.n1874 VDD.n1873 3.1005
R3645 VDD.n1557 VDD.n1551 3.1005
R3646 VDD.n1881 VDD.n1880 3.1005
R3647 VDD.n1882 VDD.n1550 3.1005
R3648 VDD.n1884 VDD.n1883 3.1005
R3649 VDD.n1892 VDD.n1891 3.1005
R3650 VDD.n1893 VDD.n1542 3.1005
R3651 VDD.n1539 VDD.n1538 3.1005
R3652 VDD.n1907 VDD.n1537 3.1005
R3653 VDD.n1909 VDD.n1908 3.1005
R3654 VDD.n1534 VDD.n1532 3.1005
R3655 VDD.n1918 VDD.n1530 3.1005
R3656 VDD.n1920 VDD.n1919 3.1005
R3657 VDD.n1531 VDD.n1524 3.1005
R3658 VDD.n1927 VDD.n1926 3.1005
R3659 VDD.n1928 VDD.n1523 3.1005
R3660 VDD.n1930 VDD.n1929 3.1005
R3661 VDD.n1519 VDD.n1518 3.1005
R3662 VDD.n1937 VDD.n1936 3.1005
R3663 VDD.n1943 VDD.n1942 3.1005
R3664 VDD.n1941 VDD.n1517 3.1005
R3665 VDD.n1950 VDD.n1512 3.1005
R3666 VDD.n1952 VDD.n1951 3.1005
R3667 VDD.n1954 VDD.n1953 3.1005
R3668 VDD.n1507 VDD.n1506 3.1005
R3669 VDD.n1962 VDD.n1961 3.1005
R3670 VDD.n1968 VDD.n1967 3.1005
R3671 VDD.n1966 VDD.n1502 3.1005
R3672 VDD.n1977 VDD.n1500 3.1005
R3673 VDD.n1496 VDD.n1495 3.1005
R3674 VDD.n1988 VDD.n1987 3.1005
R3675 VDD.n1989 VDD.n1494 3.1005
R3676 VDD.n1990 VDD.n1491 3.1005
R3677 VDD.n2000 VDD.n1490 3.1005
R3678 VDD.n2002 VDD.n2001 3.1005
R3679 VDD.n2004 VDD.n2003 3.1005
R3680 VDD.n1484 VDD.n1483 3.1005
R3681 VDD.n2010 VDD.n2009 3.1005
R3682 VDD.n2011 VDD.n1482 3.1005
R3683 VDD.n2016 VDD.n2015 3.1005
R3684 VDD.n2023 VDD.n1477 3.1005
R3685 VDD.n2025 VDD.n2024 3.1005
R3686 VDD.n2027 VDD.n2026 3.1005
R3687 VDD.n1476 VDD.n1470 3.1005
R3688 VDD.n2034 VDD.n2033 3.1005
R3689 VDD.n2035 VDD.n1469 3.1005
R3690 VDD.n2037 VDD.n2036 3.1005
R3691 VDD.n1460 VDD.n1459 3.1005
R3692 VDD.n1042 VDD.n1041 3.1005
R3693 VDD.n1043 VDD.n1027 3.1005
R3694 VDD.n1045 VDD.n1044 3.1005
R3695 VDD.n1024 VDD.n1023 3.1005
R3696 VDD.n1054 VDD.n1053 3.1005
R3697 VDD.n1055 VDD.n1022 3.1005
R3698 VDD.n1057 VDD.n1056 3.1005
R3699 VDD.n1065 VDD.n1064 3.1005
R3700 VDD.n1066 VDD.n1015 3.1005
R3701 VDD.n1068 VDD.n1067 3.1005
R3702 VDD.n1012 VDD.n1011 3.1005
R3703 VDD.n1077 VDD.n1076 3.1005
R3704 VDD.n1078 VDD.n1010 3.1005
R3705 VDD.n1080 VDD.n1079 3.1005
R3706 VDD.n1007 VDD.n1005 3.1005
R3707 VDD.n1090 VDD.n1004 3.1005
R3708 VDD.n1092 VDD.n1091 3.1005
R3709 VDD.n1001 VDD.n1000 3.1005
R3710 VDD.n1102 VDD.n999 3.1005
R3711 VDD.n1103 VDD.n996 3.1005
R3712 VDD.n1115 VDD.n1114 3.1005
R3713 VDD.n1120 VDD.n1119 3.1005
R3714 VDD.n992 VDD.n991 3.1005
R3715 VDD.n1129 VDD.n1128 3.1005
R3716 VDD.n1130 VDD.n989 3.1005
R3717 VDD.n1132 VDD.n1131 3.1005
R3718 VDD.n985 VDD.n984 3.1005
R3719 VDD.n1140 VDD.n1139 3.1005
R3720 VDD.n1145 VDD.n1144 3.1005
R3721 VDD.n980 VDD.n979 3.1005
R3722 VDD.n1152 VDD.n1151 3.1005
R3723 VDD.n1153 VDD.n976 3.1005
R3724 VDD.n1155 VDD.n1154 3.1005
R3725 VDD.n973 VDD.n972 3.1005
R3726 VDD.n1163 VDD.n1162 3.1005
R3727 VDD.n1164 VDD.n971 3.1005
R3728 VDD.n968 VDD.n967 3.1005
R3729 VDD.n1176 VDD.n1175 3.1005
R3730 VDD.n1177 VDD.n966 3.1005
R3731 VDD.n963 VDD.n961 3.1005
R3732 VDD.n1190 VDD.n960 3.1005
R3733 VDD.n1192 VDD.n1191 3.1005
R3734 VDD.n1200 VDD.n1199 3.1005
R3735 VDD.n1201 VDD.n951 3.1005
R3736 VDD.n1203 VDD.n1202 3.1005
R3737 VDD.n948 VDD.n947 3.1005
R3738 VDD.n1212 VDD.n1211 3.1005
R3739 VDD.n1213 VDD.n946 3.1005
R3740 VDD.n1215 VDD.n1214 3.1005
R3741 VDD.n1223 VDD.n1222 3.1005
R3742 VDD.n1224 VDD.n939 3.1005
R3743 VDD.n1226 VDD.n1225 3.1005
R3744 VDD.n936 VDD.n935 3.1005
R3745 VDD.n1235 VDD.n1234 3.1005
R3746 VDD.n1236 VDD.n934 3.1005
R3747 VDD.n1238 VDD.n1237 3.1005
R3748 VDD.n931 VDD.n929 3.1005
R3749 VDD.n1248 VDD.n928 3.1005
R3750 VDD.n1250 VDD.n1249 3.1005
R3751 VDD.n925 VDD.n924 3.1005
R3752 VDD.n1260 VDD.n923 3.1005
R3753 VDD.n1261 VDD.n920 3.1005
R3754 VDD.n1273 VDD.n1272 3.1005
R3755 VDD.n1278 VDD.n1277 3.1005
R3756 VDD.n916 VDD.n915 3.1005
R3757 VDD.n1287 VDD.n1286 3.1005
R3758 VDD.n1288 VDD.n913 3.1005
R3759 VDD.n1290 VDD.n1289 3.1005
R3760 VDD.n908 VDD.n907 3.1005
R3761 VDD.n1302 VDD.n1301 3.1005
R3762 VDD.n1453 VDD.n1452 3.1005
R3763 VDD.n828 VDD.n823 3.1005
R3764 VDD.n306 VDD.n286 3.1005
R3765 VDD.n395 VDD.n375 3.1005
R3766 VDD.n484 VDD.n464 3.1005
R3767 VDD.n573 VDD.n553 3.1005
R3768 VDD.n764 VDD.n763 3.1005
R3769 VDD.n251 VDD.n242 3.1005
R3770 VDD.n238 VDD.n237 3.1005
R3771 VDD.n262 VDD.n261 3.1005
R3772 VDD.n263 VDD.n236 3.1005
R3773 VDD.n264 VDD.n233 3.1005
R3774 VDD.n274 VDD.n232 3.1005
R3775 VDD.n276 VDD.n275 3.1005
R3776 VDD.n278 VDD.n277 3.1005
R3777 VDD.n226 VDD.n225 3.1005
R3778 VDD.n284 VDD.n283 3.1005
R3779 VDD.n285 VDD.n224 3.1005
R3780 VDD.n300 VDD.n299 3.1005
R3781 VDD.n313 VDD.n219 3.1005
R3782 VDD.n315 VDD.n314 3.1005
R3783 VDD.n317 VDD.n316 3.1005
R3784 VDD.n214 VDD.n213 3.1005
R3785 VDD.n325 VDD.n324 3.1005
R3786 VDD.n331 VDD.n330 3.1005
R3787 VDD.n329 VDD.n209 3.1005
R3788 VDD.n340 VDD.n207 3.1005
R3789 VDD.n203 VDD.n202 3.1005
R3790 VDD.n351 VDD.n350 3.1005
R3791 VDD.n352 VDD.n201 3.1005
R3792 VDD.n353 VDD.n198 3.1005
R3793 VDD.n363 VDD.n197 3.1005
R3794 VDD.n365 VDD.n364 3.1005
R3795 VDD.n367 VDD.n366 3.1005
R3796 VDD.n191 VDD.n190 3.1005
R3797 VDD.n373 VDD.n372 3.1005
R3798 VDD.n374 VDD.n189 3.1005
R3799 VDD.n389 VDD.n388 3.1005
R3800 VDD.n402 VDD.n184 3.1005
R3801 VDD.n404 VDD.n403 3.1005
R3802 VDD.n406 VDD.n405 3.1005
R3803 VDD.n179 VDD.n178 3.1005
R3804 VDD.n414 VDD.n413 3.1005
R3805 VDD.n420 VDD.n419 3.1005
R3806 VDD.n418 VDD.n174 3.1005
R3807 VDD.n429 VDD.n172 3.1005
R3808 VDD.n168 VDD.n167 3.1005
R3809 VDD.n440 VDD.n439 3.1005
R3810 VDD.n441 VDD.n166 3.1005
R3811 VDD.n442 VDD.n163 3.1005
R3812 VDD.n452 VDD.n162 3.1005
R3813 VDD.n454 VDD.n453 3.1005
R3814 VDD.n456 VDD.n455 3.1005
R3815 VDD.n156 VDD.n155 3.1005
R3816 VDD.n462 VDD.n461 3.1005
R3817 VDD.n463 VDD.n154 3.1005
R3818 VDD.n478 VDD.n477 3.1005
R3819 VDD.n491 VDD.n149 3.1005
R3820 VDD.n493 VDD.n492 3.1005
R3821 VDD.n495 VDD.n494 3.1005
R3822 VDD.n144 VDD.n143 3.1005
R3823 VDD.n503 VDD.n502 3.1005
R3824 VDD.n509 VDD.n508 3.1005
R3825 VDD.n507 VDD.n139 3.1005
R3826 VDD.n518 VDD.n137 3.1005
R3827 VDD.n133 VDD.n132 3.1005
R3828 VDD.n529 VDD.n528 3.1005
R3829 VDD.n530 VDD.n131 3.1005
R3830 VDD.n531 VDD.n128 3.1005
R3831 VDD.n541 VDD.n127 3.1005
R3832 VDD.n543 VDD.n542 3.1005
R3833 VDD.n545 VDD.n544 3.1005
R3834 VDD.n121 VDD.n120 3.1005
R3835 VDD.n551 VDD.n550 3.1005
R3836 VDD.n552 VDD.n119 3.1005
R3837 VDD.n567 VDD.n566 3.1005
R3838 VDD.n580 VDD.n114 3.1005
R3839 VDD.n582 VDD.n581 3.1005
R3840 VDD.n585 VDD.n584 3.1005
R3841 VDD.n583 VDD.n109 3.1005
R3842 VDD.n592 VDD.n106 3.1005
R3843 VDD.n596 VDD.n104 3.1005
R3844 VDD.n598 VDD.n597 3.1005
R3845 VDD.n100 VDD.n99 3.1005
R3846 VDD.n608 VDD.n607 3.1005
R3847 VDD.n609 VDD.n96 3.1005
R3848 VDD.n611 VDD.n610 3.1005
R3849 VDD.n92 VDD.n91 3.1005
R3850 VDD.n622 VDD.n621 3.1005
R3851 VDD.n623 VDD.n90 3.1005
R3852 VDD.n625 VDD.n624 3.1005
R3853 VDD.n627 VDD.n83 3.1005
R3854 VDD.n637 VDD.n636 3.1005
R3855 VDD.n639 VDD.n638 3.1005
R3856 VDD.n741 VDD.n740 3.1005
R3857 VDD.n742 VDD.n23 3.1005
R3858 VDD.n745 VDD.n744 3.1005
R3859 VDD.n753 VDD.n18 3.1005
R3860 VDD.n755 VDD.n754 3.1005
R3861 VDD.n757 VDD.n756 3.1005
R3862 VDD.n2744 VDD.n2743 3.1005
R3863 VDD.n2601 VDD.n2600 3.1005
R3864 VDD.n2477 VDD.n2476 3.1005
R3865 VDD.n2353 VDD.n2352 3.1005
R3866 VDD.n2279 VDD.n2278 3.1005
R3867 VDD.n2177 VDD.n2175 3.1005
R3868 VDD.n2682 VDD.n2681 3.1005
R3869 VDD.n2686 VDD.n2685 3.1005
R3870 VDD.n2692 VDD.n2691 3.1005
R3871 VDD.n2696 VDD.n2695 3.1005
R3872 VDD.n2701 VDD.n2700 3.1005
R3873 VDD.n2705 VDD.n2704 3.1005
R3874 VDD.n2709 VDD.n2708 3.1005
R3875 VDD.n2719 VDD.n2718 3.1005
R3876 VDD.n2723 VDD.n2722 3.1005
R3877 VDD.n2726 VDD.n2725 3.1005
R3878 VDD.n2730 VDD.n2729 3.1005
R3879 VDD.n2734 VDD.n2733 3.1005
R3880 VDD.n2740 VDD.n2739 3.1005
R3881 VDD.n2769 VDD.n2768 3.1005
R3882 VDD.n2773 VDD.n2772 3.1005
R3883 VDD.n2777 VDD.n2776 3.1005
R3884 VDD.n2786 VDD.n2785 3.1005
R3885 VDD.n2787 VDD.n2670 3.1005
R3886 VDD.n2799 VDD.n2798 3.1005
R3887 VDD.n2663 VDD.n2662 3.1005
R3888 VDD.n2659 VDD.n2658 3.1005
R3889 VDD.n2655 VDD.n2654 3.1005
R3890 VDD.n2649 VDD.n2648 3.1005
R3891 VDD.n2645 VDD.n2644 3.1005
R3892 VDD.n2640 VDD.n2639 3.1005
R3893 VDD.n2636 VDD.n2635 3.1005
R3894 VDD.n2626 VDD.n2625 3.1005
R3895 VDD.n2622 VDD.n2621 3.1005
R3896 VDD.n2618 VDD.n2617 3.1005
R3897 VDD.n2615 VDD.n2614 3.1005
R3898 VDD.n2611 VDD.n2610 3.1005
R3899 VDD.n2607 VDD.n2606 3.1005
R3900 VDD.n2576 VDD.n2575 3.1005
R3901 VDD.n2572 VDD.n2571 3.1005
R3902 VDD.n2568 VDD.n2567 3.1005
R3903 VDD.n2559 VDD.n2558 3.1005
R3904 VDD.n2548 VDD.n0 3.1005
R3905 VDD.n2547 VDD.n2546 3.1005
R3906 VDD.n2539 VDD.n2538 3.1005
R3907 VDD.n2535 VDD.n2534 3.1005
R3908 VDD.n2531 VDD.n2530 3.1005
R3909 VDD.n2525 VDD.n2524 3.1005
R3910 VDD.n2521 VDD.n2520 3.1005
R3911 VDD.n2516 VDD.n2515 3.1005
R3912 VDD.n2512 VDD.n2511 3.1005
R3913 VDD.n2502 VDD.n2501 3.1005
R3914 VDD.n2498 VDD.n2497 3.1005
R3915 VDD.n2494 VDD.n2493 3.1005
R3916 VDD.n2491 VDD.n2490 3.1005
R3917 VDD.n2487 VDD.n2486 3.1005
R3918 VDD.n2483 VDD.n2482 3.1005
R3919 VDD.n2452 VDD.n2451 3.1005
R3920 VDD.n2448 VDD.n2447 3.1005
R3921 VDD.n2444 VDD.n2443 3.1005
R3922 VDD.n2435 VDD.n2434 3.1005
R3923 VDD.n2424 VDD.n4 3.1005
R3924 VDD.n2423 VDD.n2422 3.1005
R3925 VDD.n2415 VDD.n2414 3.1005
R3926 VDD.n2411 VDD.n2410 3.1005
R3927 VDD.n2407 VDD.n2406 3.1005
R3928 VDD.n2401 VDD.n2400 3.1005
R3929 VDD.n2397 VDD.n2396 3.1005
R3930 VDD.n2392 VDD.n2391 3.1005
R3931 VDD.n2388 VDD.n2387 3.1005
R3932 VDD.n2378 VDD.n2377 3.1005
R3933 VDD.n2374 VDD.n2373 3.1005
R3934 VDD.n2370 VDD.n2369 3.1005
R3935 VDD.n2367 VDD.n2366 3.1005
R3936 VDD.n2363 VDD.n2362 3.1005
R3937 VDD.n2359 VDD.n2358 3.1005
R3938 VDD.n2328 VDD.n2327 3.1005
R3939 VDD.n2324 VDD.n2323 3.1005
R3940 VDD.n2320 VDD.n2319 3.1005
R3941 VDD.n2311 VDD.n2310 3.1005
R3942 VDD.n2292 VDD.n8 3.1005
R3943 VDD.n2291 VDD.n2290 3.1005
R3944 VDD.n2283 VDD.n2282 3.1005
R3945 VDD.n2263 VDD.n2262 3.1005
R3946 VDD.n2258 VDD.n2257 3.1005
R3947 VDD.n2254 VDD.n2253 3.1005
R3948 VDD.n2244 VDD.n2243 3.1005
R3949 VDD.n2240 VDD.n2239 3.1005
R3950 VDD.n2236 VDD.n2235 3.1005
R3951 VDD.n2233 VDD.n2232 3.1005
R3952 VDD.n2229 VDD.n2228 3.1005
R3953 VDD.n2225 VDD.n2224 3.1005
R3954 VDD.n2219 VDD.n2218 3.1005
R3955 VDD.n2215 VDD.n2214 3.1005
R3956 VDD.n2205 VDD.n2204 3.1005
R3957 VDD.n2201 VDD.n2200 3.1005
R3958 VDD.n2197 VDD.n2196 3.1005
R3959 VDD.n2188 VDD.n2187 3.1005
R3960 VDD.n105 VDD.n100 3.09016
R3961 VDD.n626 VDD.n625 3.09016
R3962 VDD.n1721 VDD.n1637 3.05722
R3963 VDD.n1797 VDD.n1594 3.05722
R3964 VDD.n1874 VDD.n1556 3.05722
R3965 VDD.n1950 VDD.n1513 3.05722
R3966 VDD.n2027 VDD.n1475 3.05722
R3967 VDD.n1053 VDD.n1052 3.05722
R3968 VDD.n1132 VDD.n990 3.05722
R3969 VDD.n1211 VDD.n1210 3.05722
R3970 VDD.n1290 VDD.n914 3.05722
R3971 VDD.n580 VDD.n115 3.05722
R3972 VDD.n491 VDD.n150 3.05722
R3973 VDD.n402 VDD.n185 3.05722
R3974 VDD.n313 VDD.n220 3.05722
R3975 VDD.n2262 VDD.n2261 3.05722
R3976 VDD.n2396 VDD.n2395 3.05722
R3977 VDD.n2520 VDD.n2519 3.05722
R3978 VDD.n2644 VDD.n2643 3.05722
R3979 VDD.n2700 VDD.n2699 3.05722
R3980 VDD.n291 VDD 3.02729
R3981 VDD.n380 VDD 3.02729
R3982 VDD.n469 VDD 3.02729
R3983 VDD.n558 VDD 3.02729
R3984 VDD.n2749 VDD 3.02729
R3985 VDD.n2585 VDD 3.02729
R3986 VDD.n2461 VDD 3.02729
R3987 VDD.n2337 VDD 3.02729
R3988 VDD.n293 VDD.n292 2.92946
R3989 VDD.n382 VDD.n381 2.92946
R3990 VDD.n471 VDD.n470 2.92946
R3991 VDD.n560 VDD.n559 2.92946
R3992 VDD.n2753 VDD 2.89456
R3993 VDD.n2589 VDD 2.89456
R3994 VDD.n2465 VDD 2.89456
R3995 VDD.n2341 VDD 2.89456
R3996 VDD.n1306 VDD.n903 2.86947
R3997 VDD.n1439 VDD.n1438 2.7891
R3998 VDD.n572 VDD.n564 2.64878
R3999 VDD.n483 VDD.n475 2.64878
R4000 VDD.n394 VDD.n386 2.64878
R4001 VDD.n305 VDD.n297 2.64878
R4002 VDD.n1735 VDD 2.63939
R4003 VDD VDD.n1818 2.63939
R4004 VDD.n1888 VDD 2.63939
R4005 VDD VDD.n1971 2.63939
R4006 VDD.n2795 VDD 2.63208
R4007 VDD VDD.n2550 2.63208
R4008 VDD VDD.n2426 2.63208
R4009 VDD.n2307 VDD.n2306 2.63208
R4010 VDD VDD.n2294 2.63208
R4011 VDD VDD.n2179 2.63208
R4012 VDD.n1424 VDD.n1423 2.63101
R4013 VDD VDD.n334 2.60324
R4014 VDD VDD.n423 2.60324
R4015 VDD VDD.n512 2.60324
R4016 VDD.n1110 VDD 2.58202
R4017 VDD VDD.n1184 2.58202
R4018 VDD.n1268 VDD 2.58202
R4019 VDD.t47 VDD.n1312 2.58202
R4020 VDD.n1687 VDD.n1685 2.55931
R4021 VDD.n1708 VDD.n1707 2.55931
R4022 VDD.n1764 VDD.n1763 2.55931
R4023 VDD.n1787 VDD.n1786 2.55931
R4024 VDD.n1840 VDD.n1838 2.55931
R4025 VDD.n1861 VDD.n1860 2.55931
R4026 VDD.n1917 VDD.n1916 2.55931
R4027 VDD.n1940 VDD.n1939 2.55931
R4028 VDD.n1993 VDD.n1991 2.55931
R4029 VDD.n2014 VDD.n2013 2.55931
R4030 VDD.n1018 VDD.n1016 2.55931
R4031 VDD.n1089 VDD.n1088 2.55931
R4032 VDD.n1143 VDD.n1142 2.55931
R4033 VDD.n1167 VDD.n1165 2.55931
R4034 VDD.n942 VDD.n940 2.55931
R4035 VDD.n1247 VDD.n1246 2.55931
R4036 VDD.n267 VDD.n265 2.55931
R4037 VDD.n356 VDD.n354 2.55931
R4038 VDD.n445 VDD.n443 2.55931
R4039 VDD.n534 VDD.n532 2.55931
R4040 VDD.n2715 VDD.n2714 2.55931
R4041 VDD.n2632 VDD.n2631 2.55931
R4042 VDD.n2508 VDD.n2507 2.55931
R4043 VDD.n2384 VDD.n2383 2.55931
R4044 VDD.n2250 VDD.n2249 2.55931
R4045 VDD.n2211 VDD.n2210 2.55931
R4046 VDD.n294 VDD.n287 2.52171
R4047 VDD.n383 VDD.n376 2.52171
R4048 VDD.n472 VDD.n465 2.52171
R4049 VDD.n561 VDD.n554 2.52171
R4050 VDD.n2755 VDD.n2754 2.52171
R4051 VDD.n2591 VDD.n2590 2.52171
R4052 VDD.n2467 VDD.n2466 2.52171
R4053 VDD.n2343 VDD.n2342 2.52171
R4054 VDD.n1673 VDD.n1672 2.5203
R4055 VDD.n1753 VDD.n1752 2.5203
R4056 VDD.n1826 VDD.n1825 2.5203
R4057 VDD.n1906 VDD.n1905 2.5203
R4058 VDD.n1979 VDD.n1978 2.5203
R4059 VDD.n1101 VDD.n1100 2.5203
R4060 VDD.n1179 VDD.n1178 2.5203
R4061 VDD.n1259 VDD.n1258 2.5203
R4062 VDD.n253 VDD.n252 2.5203
R4063 VDD.n342 VDD.n341 2.5203
R4064 VDD.n431 VDD.n430 2.5203
R4065 VDD.n520 VDD.n519 2.5203
R4066 VDD.n2782 VDD.n2781 2.5203
R4067 VDD.n2564 VDD.n2563 2.5203
R4068 VDD.n2440 VDD.n2439 2.5203
R4069 VDD.n2316 VDD.n2315 2.5203
R4070 VDD.n2193 VDD.n2192 2.5203
R4071 VDD.n2077 VDD.n2076 2.51325
R4072 VDD.n2096 VDD.n2094 2.49102
R4073 VDD.n2152 VDD.n2061 2.49102
R4074 VDD.n2051 VDD.n2049 2.49102
R4075 VDD.n1670 VDD.n1669 2.49102
R4076 VDD.n1743 VDD.n1741 2.49102
R4077 VDD.n1823 VDD.n1822 2.49102
R4078 VDD.n1896 VDD.n1894 2.49102
R4079 VDD.n1976 VDD.n1975 2.49102
R4080 VDD.n1106 VDD.n1104 2.49102
R4081 VDD.n1189 VDD.n1188 2.49102
R4082 VDD.n1264 VDD.n1262 2.49102
R4083 VDD.n250 VDD.n249 2.49102
R4084 VDD.n339 VDD.n338 2.49102
R4085 VDD.n428 VDD.n427 2.49102
R4086 VDD.n517 VDD.n516 2.49102
R4087 VDD.n743 VDD.n25 2.49102
R4088 VDD.n14 VDD.n12 2.49102
R4089 VDD.n2790 VDD.n2788 2.49102
R4090 VDD.n2555 VDD.n2554 2.49102
R4091 VDD.n2431 VDD.n2430 2.49102
R4092 VDD.n2299 VDD.n2298 2.49102
R4093 VDD.n2184 VDD.n2183 2.49102
R4094 VDD.n792 VDD.n791 2.44756
R4095 VDD.n1626 VDD.n1624 2.43201
R4096 VDD.n1812 VDD.n1811 2.43201
R4097 VDD.n1545 VDD.n1543 2.43201
R4098 VDD.n1965 VDD.n1964 2.43201
R4099 VDD.n1464 VDD.n1462 2.43201
R4100 VDD.n1032 VDD.n1030 2.43201
R4101 VDD.n1118 VDD.n1117 2.43201
R4102 VDD.n956 VDD.n954 2.43201
R4103 VDD.n1276 VDD.n1275 2.43201
R4104 VDD.n328 VDD.n327 2.43201
R4105 VDD.n417 VDD.n416 2.43201
R4106 VDD.n506 VDD.n505 2.43201
R4107 VDD.n595 VDD.n594 2.43201
R4108 VDD.n2678 VDD.n2677 2.43201
R4109 VDD.n2669 VDD.n2668 2.43201
R4110 VDD.n2545 VDD.n2544 2.43201
R4111 VDD.n2421 VDD.n2420 2.43201
R4112 VDD.n2289 VDD.n2288 2.43201
R4113 VDD.n1306 VDD.n1305 2.42487
R4114 VDD.n1386 VDD.n1385 2.42487
R4115 VDD.n1388 VDD.n1387 2.35689
R4116 VDD.n1294 VDD.n906 2.35689
R4117 VDD.n1418 VDD.n844 2.35366
R4118 VDD.n1441 VDD.n1440 2.35119
R4119 VDD.n795 VDD.n780 2.28739
R4120 VDD.n811 VDD.n770 2.28739
R4121 VDD.n768 VDD.n766 2.27014
R4122 VDD.n796 VDD.n767 2.25996
R4123 VDD.n1695 VDD.n1651 2.2074
R4124 VDD.n1612 VDD.n1607 2.2074
R4125 VDD.n1848 VDD.n1570 2.2074
R4126 VDD.n1531 VDD.n1526 2.2074
R4127 VDD.n2001 VDD.n1489 2.2074
R4128 VDD.n1075 VDD.n1010 2.2074
R4129 VDD.n978 VDD.n973 2.2074
R4130 VDD.n1233 VDD.n934 2.2074
R4131 VDD.n1310 VDD.n1309 2.2074
R4132 VDD.n1321 VDD.n895 2.2074
R4133 VDD.n1329 VDD.n1328 2.2074
R4134 VDD.n1340 VDD.n885 2.2074
R4135 VDD.n1347 VDD.n1346 2.2074
R4136 VDD.n1369 VDD.n871 2.2074
R4137 VDD.n1377 VDD.n1376 2.2074
R4138 VDD.n1395 VDD.n1394 2.2074
R4139 VDD.n1406 VDD.n853 2.2074
R4140 VDD.n1414 VDD.n1413 2.2074
R4141 VDD.n1430 VDD.n1429 2.2074
R4142 VDD.n1448 VDD.n1447 2.2074
R4143 VDD.n639 VDD.n82 2.2074
R4144 VDD.n648 VDD.n647 2.2074
R4145 VDD.n653 VDD.n652 2.2074
R4146 VDD.n652 VDD.n70 2.2074
R4147 VDD.n665 VDD.n66 2.2074
R4148 VDD.n665 VDD.n68 2.2074
R4149 VDD.n673 VDD.n672 2.2074
R4150 VDD.n673 VDD.n60 2.2074
R4151 VDD.n685 VDD.n55 2.2074
R4152 VDD.n686 VDD.n685 2.2074
R4153 VDD.n691 VDD.n690 2.2074
R4154 VDD.n690 VDD.n48 2.2074
R4155 VDD.n703 VDD.n44 2.2074
R4156 VDD.n703 VDD.n46 2.2074
R4157 VDD.n711 VDD.n710 2.2074
R4158 VDD.n711 VDD.n38 2.2074
R4159 VDD.n723 VDD.n33 2.2074
R4160 VDD.n724 VDD.n723 2.2074
R4161 VDD.n732 VDD.n731 2.2074
R4162 VDD.n542 VDD.n126 2.2074
R4163 VDD.n453 VDD.n161 2.2074
R4164 VDD.n364 VDD.n196 2.2074
R4165 VDD.n275 VDD.n231 2.2074
R4166 VDD.n2224 VDD.n2221 2.2074
R4167 VDD.n2358 VDD.n2355 2.2074
R4168 VDD.n2347 VDD.n2334 2.2074
R4169 VDD.n2482 VDD.n2479 2.2074
R4170 VDD.n2471 VDD.n2458 2.2074
R4171 VDD.n2606 VDD.n2603 2.2074
R4172 VDD.n2595 VDD.n2582 2.2074
R4173 VDD.n2739 VDD.n2736 2.2074
R4174 VDD.n2759 VDD.n2746 2.2074
R4175 VDD.n815 VDD.n773 2.07109
R4176 VDD.n572 VDD.n571 2.02155
R4177 VDD.n483 VDD.n482 2.02155
R4178 VDD.n394 VDD.n393 2.02155
R4179 VDD.n305 VDD.n304 2.02155
R4180 VDD.n2331 VDD.n2329 2.02155
R4181 VDD.n2455 VDD.n2453 2.02155
R4182 VDD.n2579 VDD.n2577 2.02155
R4183 VDD.n2764 VDD.n2762 2.02155
R4184 VDD.n1309 VDD.n899 1.98671
R4185 VDD.n1321 VDD.n897 1.98671
R4186 VDD.n1329 VDD.n889 1.98671
R4187 VDD.n1341 VDD.n1340 1.98671
R4188 VDD.n1346 VDD.n883 1.98671
R4189 VDD.n1358 VDD.n875 1.98671
R4190 VDD.n1370 VDD.n1369 1.98671
R4191 VDD.n1376 VDD.n869 1.98671
R4192 VDD.n1395 VDD.n857 1.98671
R4193 VDD.n1407 VDD.n1406 1.98671
R4194 VDD.n1413 VDD.n851 1.98671
R4195 VDD.n1429 VDD.n841 1.98671
R4196 VDD.n1449 VDD.n1448 1.98671
R4197 VDD VDD.n290 1.91393
R4198 VDD VDD.n379 1.91393
R4199 VDD VDD.n468 1.91393
R4200 VDD VDD.n557 1.91393
R4201 VDD VDD.n2748 1.85046
R4202 VDD VDD.n2584 1.85046
R4203 VDD VDD.n2460 1.85046
R4204 VDD VDD.n2336 1.85046
R4205 VDD.n1317 VDD.n899 1.76602
R4206 VDD.n897 VDD.n896 1.76602
R4207 VDD.n1333 VDD.n889 1.76602
R4208 VDD.n1342 VDD.n1341 1.76602
R4209 VDD.n883 VDD.n877 1.76602
R4210 VDD.n1357 VDD.n877 1.76602
R4211 VDD.n1362 VDD.n875 1.76602
R4212 VDD.n1371 VDD.n1370 1.76602
R4213 VDD.n869 VDD.n863 1.76602
R4214 VDD.n1399 VDD.n857 1.76602
R4215 VDD.n1408 VDD.n1407 1.76602
R4216 VDD.n851 VDD.n843 1.76602
R4217 VDD.n841 VDD.n834 1.76602
R4218 VDD.n1449 VDD.n827 1.76602
R4219 VDD.n647 VDD.n78 1.76602
R4220 VDD.n1627 VDD.n1626 1.72554
R4221 VDD.n1811 VDD.n1586 1.72554
R4222 VDD.n1546 VDD.n1545 1.72554
R4223 VDD.n1964 VDD.n1505 1.72554
R4224 VDD.n1465 VDD.n1464 1.72554
R4225 VDD.n1033 VDD.n1032 1.72554
R4226 VDD.n1117 VDD.n995 1.72554
R4227 VDD.n957 VDD.n956 1.72554
R4228 VDD.n1275 VDD.n919 1.72554
R4229 VDD.n327 VDD.n212 1.72554
R4230 VDD.n416 VDD.n177 1.72554
R4231 VDD.n505 VDD.n142 1.72554
R4232 VDD.n594 VDD.n593 1.72554
R4233 VDD.n2677 VDD.n2676 1.72554
R4234 VDD.n2668 VDD.n2667 1.72554
R4235 VDD.n2544 VDD.n2543 1.72554
R4236 VDD.n2420 VDD.n2419 1.72554
R4237 VDD.n2288 VDD.n2287 1.72554
R4238 VDD.n2097 VDD.n2096 1.57241
R4239 VDD.n2155 VDD.n2061 1.57241
R4240 VDD.n2052 VDD.n2051 1.57241
R4241 VDD.n1669 VDD.n1668 1.57241
R4242 VDD.n1744 VDD.n1743 1.57241
R4243 VDD.n1822 VDD.n1821 1.57241
R4244 VDD.n1897 VDD.n1896 1.57241
R4245 VDD.n1975 VDD.n1974 1.57241
R4246 VDD.n1107 VDD.n1106 1.57241
R4247 VDD.n1188 VDD.n1187 1.57241
R4248 VDD.n1265 VDD.n1264 1.57241
R4249 VDD.n249 VDD.n248 1.57241
R4250 VDD.n338 VDD.n337 1.57241
R4251 VDD.n427 VDD.n426 1.57241
R4252 VDD.n516 VDD.n515 1.57241
R4253 VDD.n746 VDD.n25 1.57241
R4254 VDD.n15 VDD.n14 1.57241
R4255 VDD.n2791 VDD.n2790 1.57241
R4256 VDD.n2554 VDD.n2553 1.57241
R4257 VDD.n2430 VDD.n2429 1.57241
R4258 VDD.n2298 VDD.n2297 1.57241
R4259 VDD.n2183 VDD.n2182 1.57241
R4260 VDD.n1310 VDD.n903 1.54533
R4261 VDD.n1316 VDD.n895 1.54533
R4262 VDD.n1328 VDD.n891 1.54533
R4263 VDD.n1334 VDD.n885 1.54533
R4264 VDD.n1347 VDD.n882 1.54533
R4265 VDD.n1363 VDD.n871 1.54533
R4266 VDD.n1377 VDD.n868 1.54533
R4267 VDD.n1394 VDD.n859 1.54533
R4268 VDD.n1400 VDD.n853 1.54533
R4269 VDD.n1414 VDD.n850 1.54533
R4270 VDD.n1430 VDD.n840 1.54533
R4271 VDD.n1447 VDD.n830 1.54533
R4272 VDD.n641 VDD.n640 1.54533
R4273 VDD.n649 VDD.n648 1.54533
R4274 VDD.n653 VDD.n75 1.54533
R4275 VDD.n661 VDD.n70 1.54533
R4276 VDD.n660 VDD.n659 1.54533
R4277 VDD.n659 VDD.n66 1.54533
R4278 VDD.n68 VDD.n67 1.54533
R4279 VDD.n672 VDD.n62 1.54533
R4280 VDD.n677 VDD.n60 1.54533
R4281 VDD.n679 VDD.n55 1.54533
R4282 VDD.n687 VDD.n686 1.54533
R4283 VDD.n691 VDD.n53 1.54533
R4284 VDD.n699 VDD.n48 1.54533
R4285 VDD.n697 VDD.n44 1.54533
R4286 VDD.n46 VDD.n45 1.54533
R4287 VDD.n710 VDD.n40 1.54533
R4288 VDD.n715 VDD.n38 1.54533
R4289 VDD.n717 VDD.n33 1.54533
R4290 VDD.n725 VDD.n724 1.54533
R4291 VDD.n732 VDD.n30 1.54533
R4292 VDD.n728 VDD.n26 1.54533
R4293 VDD.n2347 VDD.n2346 1.54533
R4294 VDD.n2471 VDD.n2470 1.54533
R4295 VDD.n2595 VDD.n2594 1.54533
R4296 VDD.n2759 VDD.n2758 1.54533
R4297 VDD.n2078 VDD.n2077 1.5148
R4298 VDD.n1674 VDD.n1673 1.49652
R4299 VDD.n1752 VDD.n1751 1.49652
R4300 VDD.n1827 VDD.n1826 1.49652
R4301 VDD.n1905 VDD.n1904 1.49652
R4302 VDD.n1980 VDD.n1979 1.49652
R4303 VDD.n1100 VDD.n1099 1.49652
R4304 VDD.n1180 VDD.n1179 1.49652
R4305 VDD.n1258 VDD.n1257 1.49652
R4306 VDD.n254 VDD.n253 1.49652
R4307 VDD.n343 VDD.n342 1.49652
R4308 VDD.n432 VDD.n431 1.49652
R4309 VDD.n521 VDD.n520 1.49652
R4310 VDD.n2781 VDD.n2780 1.49652
R4311 VDD.n2563 VDD.n2562 1.49652
R4312 VDD.n2439 VDD.n2438 1.49652
R4313 VDD.n2315 VDD.n2314 1.49652
R4314 VDD.n2192 VDD.n2191 1.49652
R4315 VDD.n2269 VDD.n2267 1.43334
R4316 VDD.n1688 VDD.n1687 1.39551
R4317 VDD.n1707 VDD.n1640 1.39551
R4318 VDD.n1763 VDD.n1762 1.39551
R4319 VDD.n1786 VDD.n1597 1.39551
R4320 VDD.n1841 VDD.n1840 1.39551
R4321 VDD.n1860 VDD.n1559 1.39551
R4322 VDD.n1916 VDD.n1915 1.39551
R4323 VDD.n1939 VDD.n1516 1.39551
R4324 VDD.n1994 VDD.n1993 1.39551
R4325 VDD.n2013 VDD.n1478 1.39551
R4326 VDD.n1019 VDD.n1018 1.39551
R4327 VDD.n1088 VDD.n1087 1.39551
R4328 VDD.n1142 VDD.n983 1.39551
R4329 VDD.n1168 VDD.n1167 1.39551
R4330 VDD.n943 VDD.n942 1.39551
R4331 VDD.n1246 VDD.n1245 1.39551
R4332 VDD.n268 VDD.n267 1.39551
R4333 VDD.n357 VDD.n356 1.39551
R4334 VDD.n446 VDD.n445 1.39551
R4335 VDD.n535 VDD.n534 1.39551
R4336 VDD.n2714 VDD.n2713 1.39551
R4337 VDD.n2631 VDD.n2630 1.39551
R4338 VDD.n2507 VDD.n2506 1.39551
R4339 VDD.n2383 VDD.n2382 1.39551
R4340 VDD.n2249 VDD.n2248 1.39551
R4341 VDD.n2210 VDD.n2209 1.39551
R4342 VDD.n728 VDD.n31 1.32464
R4343 VDD.n815 VDD.n774 1.12991
R4344 VDD.n2137 VDD.n2071 1.10395
R4345 VDD.n2162 VDD.n2057 1.10395
R4346 VDD.n753 VDD.n20 1.10395
R4347 VDD.n807 VDD.n777 0.941676
R4348 VDD.n731 VDD.n31 0.883259
R4349 VDD.n293 VDD.n287 0.776258
R4350 VDD.n382 VDD.n376 0.776258
R4351 VDD.n471 VDD.n465 0.776258
R4352 VDD.n560 VDD.n554 0.776258
R4353 VDD.n791 VDD.n790 0.753441
R4354 VDD.n290 VDD.n289 0.750619
R4355 VDD.n379 VDD.n378 0.750619
R4356 VDD.n468 VDD.n467 0.750619
R4357 VDD.n557 VDD.n556 0.750619
R4358 VDD.n2141 VDD.n2068 0.662569
R4359 VDD.n1306 VDD.n905 0.662569
R4360 VDD.n716 VDD.n715 0.662569
R4361 VDD.n2150 VDD 0.622896
R4362 VDD.n1727 VDD.n1634 0.478112
R4363 VDD.n1801 VDD.n1592 0.478112
R4364 VDD.n1880 VDD.n1553 0.478112
R4365 VDD.n1954 VDD.n1511 0.478112
R4366 VDD.n2033 VDD.n1472 0.478112
R4367 VDD.n1045 VDD.n1029 0.478112
R4368 VDD.n1128 VDD.n1127 0.478112
R4369 VDD.n1203 VDD.n953 0.478112
R4370 VDD.n1286 VDD.n1285 0.478112
R4371 VDD.n585 VDD.n113 0.478112
R4372 VDD.n495 VDD.n148 0.478112
R4373 VDD.n406 VDD.n183 0.478112
R4374 VDD.n317 VDD.n218 0.478112
R4375 VDD.n2274 VDD.n2273 0.478112
R4376 VDD.n2406 VDD.n2405 0.478112
R4377 VDD.n2530 VDD.n2529 0.478112
R4378 VDD.n2654 VDD.n2653 0.478112
R4379 VDD.n2691 VDD.n2690 0.478112
R4380 VDD.n636 VDD.n85 0.441879
R4381 VDD.n640 VDD.n78 0.441879
R4382 VDD.n632 VDD.n87 0.426767
R4383 VDD.n87 VDD.n82 0.426767
R4384 VDD.n2754 VDD.n2753 0.373349
R4385 VDD.n2590 VDD.n2589 0.373349
R4386 VDD.n2466 VDD.n2465 0.373349
R4387 VDD.n2342 VDD.n2341 0.373349
R4388 VDD.n2346 VDD.n2345 0.332764
R4389 VDD.n2470 VDD.n2469 0.332063
R4390 VDD.n2594 VDD.n2593 0.332063
R4391 VDD.n2758 VDD.n2757 0.331371
R4392 VDD.n1461 VDD 0.282678
R4393 VDD.n291 VDD 0.259429
R4394 VDD.n380 VDD 0.259429
R4395 VDD.n469 VDD 0.259429
R4396 VDD.n558 VDD 0.259429
R4397 VDD.n2749 VDD 0.259429
R4398 VDD.n2585 VDD 0.259429
R4399 VDD.n2461 VDD 0.259429
R4400 VDD.n2337 VDD 0.259429
R4401 VDD.n2267 VDD.n2266 0.225571
R4402 VDD.n1358 VDD.n1357 0.22119
R4403 VDD.n740 VDD.n739 0.22119
R4404 VDD.n2310 VDD.n2302 0.22119
R4405 VDD.n788 VDD.n765 0.213502
R4406 VDD.n1461 VDD.n765 0.20861
R4407 VDD.n2269 VDD.n2268 0.191545
R4408 VDD.n800 VDD.n780 0.188735
R4409 VDD.n798 VDD.n782 0.188735
R4410 VDD.n2048 VDD 0.151171
R4411 VDD.n2094 VDD.n2089 0.120292
R4412 VDD.n2105 VDD.n2089 0.120292
R4413 VDD.n2106 VDD.n2105 0.120292
R4414 VDD.n2107 VDD.n2106 0.120292
R4415 VDD.n2107 VDD.n2082 0.120292
R4416 VDD.n2116 VDD.n2082 0.120292
R4417 VDD.n2117 VDD.n2116 0.120292
R4418 VDD.n2118 VDD.n2117 0.120292
R4419 VDD.n2118 VDD.n2076 0.120292
R4420 VDD.n2127 VDD.n2076 0.120292
R4421 VDD.n2128 VDD.n2127 0.120292
R4422 VDD.n2129 VDD.n2128 0.120292
R4423 VDD.n2129 VDD.n2069 0.120292
R4424 VDD.n2138 VDD.n2069 0.120292
R4425 VDD.n2139 VDD.n2138 0.120292
R4426 VDD.n2140 VDD.n2139 0.120292
R4427 VDD.n2140 VDD.n2062 0.120292
R4428 VDD.n2148 VDD.n2062 0.120292
R4429 VDD.n2151 VDD.n2150 0.120292
R4430 VDD.n2152 VDD.n2151 0.120292
R4431 VDD.n2153 VDD.n2152 0.120292
R4432 VDD.n2153 VDD.n2055 0.120292
R4433 VDD.n2164 VDD.n2055 0.120292
R4434 VDD.n2165 VDD.n2049 0.120292
R4435 VDD.n2173 VDD.n2049 0.120292
R4436 VDD.n1671 VDD.n1670 0.120292
R4437 VDD.n1672 VDD.n1671 0.120292
R4438 VDD.n1672 VDD.n1657 0.120292
R4439 VDD.n1682 VDD.n1657 0.120292
R4440 VDD.n1683 VDD.n1682 0.120292
R4441 VDD.n1685 VDD.n1683 0.120292
R4442 VDD.n1685 VDD.n1684 0.120292
R4443 VDD.n1684 VDD.n1652 0.120292
R4444 VDD.n1696 VDD.n1652 0.120292
R4445 VDD.n1697 VDD.n1696 0.120292
R4446 VDD.n1697 VDD.n1645 0.120292
R4447 VDD.n1704 VDD.n1645 0.120292
R4448 VDD.n1705 VDD.n1704 0.120292
R4449 VDD.n1709 VDD.n1705 0.120292
R4450 VDD.n1709 VDD.n1708 0.120292
R4451 VDD.n1708 VDD.n1639 0.120292
R4452 VDD.n1719 VDD.n1639 0.120292
R4453 VDD.n1720 VDD.n1719 0.120292
R4454 VDD.n1720 VDD.n1632 0.120292
R4455 VDD.n1728 VDD.n1632 0.120292
R4456 VDD.n1729 VDD.n1728 0.120292
R4457 VDD.n1730 VDD.n1729 0.120292
R4458 VDD.n1730 VDD.n1624 0.120292
R4459 VDD.n1739 VDD.n1624 0.120292
R4460 VDD.n1741 VDD.n1619 0.120292
R4461 VDD.n1753 VDD.n1619 0.120292
R4462 VDD.n1754 VDD.n1753 0.120292
R4463 VDD.n1755 VDD.n1754 0.120292
R4464 VDD.n1755 VDD.n1613 0.120292
R4465 VDD.n1764 VDD.n1613 0.120292
R4466 VDD.n1765 VDD.n1764 0.120292
R4467 VDD.n1766 VDD.n1765 0.120292
R4468 VDD.n1766 VDD.n1605 0.120292
R4469 VDD.n1774 VDD.n1605 0.120292
R4470 VDD.n1775 VDD.n1774 0.120292
R4471 VDD.n1776 VDD.n1775 0.120292
R4472 VDD.n1776 VDD.n1599 0.120292
R4473 VDD.n1784 VDD.n1599 0.120292
R4474 VDD.n1787 VDD.n1784 0.120292
R4475 VDD.n1789 VDD.n1787 0.120292
R4476 VDD.n1789 VDD.n1788 0.120292
R4477 VDD.n1788 VDD.n1593 0.120292
R4478 VDD.n1799 VDD.n1593 0.120292
R4479 VDD.n1800 VDD.n1799 0.120292
R4480 VDD.n1800 VDD.n1587 0.120292
R4481 VDD.n1809 VDD.n1587 0.120292
R4482 VDD.n1812 VDD.n1809 0.120292
R4483 VDD.n1814 VDD.n1812 0.120292
R4484 VDD.n1824 VDD.n1823 0.120292
R4485 VDD.n1825 VDD.n1824 0.120292
R4486 VDD.n1825 VDD.n1576 0.120292
R4487 VDD.n1835 VDD.n1576 0.120292
R4488 VDD.n1836 VDD.n1835 0.120292
R4489 VDD.n1838 VDD.n1836 0.120292
R4490 VDD.n1838 VDD.n1837 0.120292
R4491 VDD.n1837 VDD.n1571 0.120292
R4492 VDD.n1849 VDD.n1571 0.120292
R4493 VDD.n1850 VDD.n1849 0.120292
R4494 VDD.n1850 VDD.n1564 0.120292
R4495 VDD.n1857 VDD.n1564 0.120292
R4496 VDD.n1858 VDD.n1857 0.120292
R4497 VDD.n1862 VDD.n1858 0.120292
R4498 VDD.n1862 VDD.n1861 0.120292
R4499 VDD.n1861 VDD.n1558 0.120292
R4500 VDD.n1872 VDD.n1558 0.120292
R4501 VDD.n1873 VDD.n1872 0.120292
R4502 VDD.n1873 VDD.n1551 0.120292
R4503 VDD.n1881 VDD.n1551 0.120292
R4504 VDD.n1882 VDD.n1881 0.120292
R4505 VDD.n1883 VDD.n1882 0.120292
R4506 VDD.n1883 VDD.n1543 0.120292
R4507 VDD.n1892 VDD.n1543 0.120292
R4508 VDD.n1894 VDD.n1538 0.120292
R4509 VDD.n1906 VDD.n1538 0.120292
R4510 VDD.n1907 VDD.n1906 0.120292
R4511 VDD.n1908 VDD.n1907 0.120292
R4512 VDD.n1908 VDD.n1532 0.120292
R4513 VDD.n1917 VDD.n1532 0.120292
R4514 VDD.n1918 VDD.n1917 0.120292
R4515 VDD.n1919 VDD.n1918 0.120292
R4516 VDD.n1919 VDD.n1524 0.120292
R4517 VDD.n1927 VDD.n1524 0.120292
R4518 VDD.n1928 VDD.n1927 0.120292
R4519 VDD.n1929 VDD.n1928 0.120292
R4520 VDD.n1929 VDD.n1518 0.120292
R4521 VDD.n1937 VDD.n1518 0.120292
R4522 VDD.n1940 VDD.n1937 0.120292
R4523 VDD.n1942 VDD.n1940 0.120292
R4524 VDD.n1942 VDD.n1941 0.120292
R4525 VDD.n1941 VDD.n1512 0.120292
R4526 VDD.n1952 VDD.n1512 0.120292
R4527 VDD.n1953 VDD.n1952 0.120292
R4528 VDD.n1953 VDD.n1506 0.120292
R4529 VDD.n1962 VDD.n1506 0.120292
R4530 VDD.n1965 VDD.n1962 0.120292
R4531 VDD.n1967 VDD.n1965 0.120292
R4532 VDD.n1977 VDD.n1976 0.120292
R4533 VDD.n1978 VDD.n1977 0.120292
R4534 VDD.n1978 VDD.n1495 0.120292
R4535 VDD.n1988 VDD.n1495 0.120292
R4536 VDD.n1989 VDD.n1988 0.120292
R4537 VDD.n1991 VDD.n1989 0.120292
R4538 VDD.n1991 VDD.n1990 0.120292
R4539 VDD.n1990 VDD.n1490 0.120292
R4540 VDD.n2002 VDD.n1490 0.120292
R4541 VDD.n2003 VDD.n2002 0.120292
R4542 VDD.n2003 VDD.n1483 0.120292
R4543 VDD.n2010 VDD.n1483 0.120292
R4544 VDD.n2011 VDD.n2010 0.120292
R4545 VDD.n2015 VDD.n2011 0.120292
R4546 VDD.n2015 VDD.n2014 0.120292
R4547 VDD.n2014 VDD.n1477 0.120292
R4548 VDD.n2025 VDD.n1477 0.120292
R4549 VDD.n2026 VDD.n2025 0.120292
R4550 VDD.n2026 VDD.n1470 0.120292
R4551 VDD.n2034 VDD.n1470 0.120292
R4552 VDD.n2035 VDD.n2034 0.120292
R4553 VDD.n2036 VDD.n2035 0.120292
R4554 VDD.n2036 VDD.n1462 0.120292
R4555 VDD.n2043 VDD.n1462 0.120292
R4556 VDD.n1042 VDD.n1030 0.120292
R4557 VDD.n1043 VDD.n1042 0.120292
R4558 VDD.n1044 VDD.n1043 0.120292
R4559 VDD.n1044 VDD.n1023 0.120292
R4560 VDD.n1054 VDD.n1023 0.120292
R4561 VDD.n1055 VDD.n1054 0.120292
R4562 VDD.n1056 VDD.n1055 0.120292
R4563 VDD.n1056 VDD.n1016 0.120292
R4564 VDD.n1065 VDD.n1016 0.120292
R4565 VDD.n1066 VDD.n1065 0.120292
R4566 VDD.n1067 VDD.n1066 0.120292
R4567 VDD.n1067 VDD.n1011 0.120292
R4568 VDD.n1077 VDD.n1011 0.120292
R4569 VDD.n1078 VDD.n1077 0.120292
R4570 VDD.n1079 VDD.n1078 0.120292
R4571 VDD.n1079 VDD.n1005 0.120292
R4572 VDD.n1089 VDD.n1005 0.120292
R4573 VDD.n1090 VDD.n1089 0.120292
R4574 VDD.n1091 VDD.n1090 0.120292
R4575 VDD.n1091 VDD.n1000 0.120292
R4576 VDD.n1101 VDD.n1000 0.120292
R4577 VDD.n1102 VDD.n1101 0.120292
R4578 VDD.n1104 VDD.n1102 0.120292
R4579 VDD.n1104 VDD.n1103 0.120292
R4580 VDD.n1118 VDD.n1115 0.120292
R4581 VDD.n1119 VDD.n1118 0.120292
R4582 VDD.n1119 VDD.n991 0.120292
R4583 VDD.n1129 VDD.n991 0.120292
R4584 VDD.n1130 VDD.n1129 0.120292
R4585 VDD.n1131 VDD.n1130 0.120292
R4586 VDD.n1131 VDD.n984 0.120292
R4587 VDD.n1140 VDD.n984 0.120292
R4588 VDD.n1143 VDD.n1140 0.120292
R4589 VDD.n1144 VDD.n1143 0.120292
R4590 VDD.n1144 VDD.n979 0.120292
R4591 VDD.n1152 VDD.n979 0.120292
R4592 VDD.n1153 VDD.n1152 0.120292
R4593 VDD.n1154 VDD.n1153 0.120292
R4594 VDD.n1154 VDD.n972 0.120292
R4595 VDD.n1163 VDD.n972 0.120292
R4596 VDD.n1164 VDD.n1163 0.120292
R4597 VDD.n1165 VDD.n1164 0.120292
R4598 VDD.n1165 VDD.n967 0.120292
R4599 VDD.n1176 VDD.n967 0.120292
R4600 VDD.n1177 VDD.n1176 0.120292
R4601 VDD.n1178 VDD.n1177 0.120292
R4602 VDD.n1178 VDD.n961 0.120292
R4603 VDD.n1189 VDD.n961 0.120292
R4604 VDD.n1190 VDD.n1189 0.120292
R4605 VDD.n1191 VDD.n954 0.120292
R4606 VDD.n1200 VDD.n954 0.120292
R4607 VDD.n1201 VDD.n1200 0.120292
R4608 VDD.n1202 VDD.n1201 0.120292
R4609 VDD.n1202 VDD.n947 0.120292
R4610 VDD.n1212 VDD.n947 0.120292
R4611 VDD.n1213 VDD.n1212 0.120292
R4612 VDD.n1214 VDD.n1213 0.120292
R4613 VDD.n1214 VDD.n940 0.120292
R4614 VDD.n1223 VDD.n940 0.120292
R4615 VDD.n1224 VDD.n1223 0.120292
R4616 VDD.n1225 VDD.n1224 0.120292
R4617 VDD.n1225 VDD.n935 0.120292
R4618 VDD.n1235 VDD.n935 0.120292
R4619 VDD.n1236 VDD.n1235 0.120292
R4620 VDD.n1237 VDD.n1236 0.120292
R4621 VDD.n1237 VDD.n929 0.120292
R4622 VDD.n1247 VDD.n929 0.120292
R4623 VDD.n1248 VDD.n1247 0.120292
R4624 VDD.n1249 VDD.n1248 0.120292
R4625 VDD.n1249 VDD.n924 0.120292
R4626 VDD.n1259 VDD.n924 0.120292
R4627 VDD.n1260 VDD.n1259 0.120292
R4628 VDD.n1262 VDD.n1260 0.120292
R4629 VDD.n1262 VDD.n1261 0.120292
R4630 VDD.n1276 VDD.n1273 0.120292
R4631 VDD.n1277 VDD.n1276 0.120292
R4632 VDD.n1277 VDD.n915 0.120292
R4633 VDD.n1287 VDD.n915 0.120292
R4634 VDD.n1288 VDD.n1287 0.120292
R4635 VDD.n1289 VDD.n1288 0.120292
R4636 VDD.n1289 VDD.n907 0.120292
R4637 VDD.n1302 VDD.n907 0.120292
R4638 VDD.n1452 VDD.n823 0.120292
R4639 VDD.n1460 VDD.n823 0.120292
R4640 VDD.n251 VDD.n250 0.120292
R4641 VDD.n252 VDD.n251 0.120292
R4642 VDD.n252 VDD.n237 0.120292
R4643 VDD.n262 VDD.n237 0.120292
R4644 VDD.n263 VDD.n262 0.120292
R4645 VDD.n265 VDD.n263 0.120292
R4646 VDD.n265 VDD.n264 0.120292
R4647 VDD.n264 VDD.n232 0.120292
R4648 VDD.n276 VDD.n232 0.120292
R4649 VDD.n277 VDD.n276 0.120292
R4650 VDD.n277 VDD.n225 0.120292
R4651 VDD.n284 VDD.n225 0.120292
R4652 VDD.n285 VDD.n284 0.120292
R4653 VDD.n286 VDD.n285 0.120292
R4654 VDD.n303 VDD.n286 0.120292
R4655 VDD.n303 VDD.n302 0.120292
R4656 VDD.n302 VDD.n299 0.120292
R4657 VDD.n299 VDD.n219 0.120292
R4658 VDD.n315 VDD.n219 0.120292
R4659 VDD.n316 VDD.n315 0.120292
R4660 VDD.n316 VDD.n213 0.120292
R4661 VDD.n325 VDD.n213 0.120292
R4662 VDD.n328 VDD.n325 0.120292
R4663 VDD.n330 VDD.n328 0.120292
R4664 VDD.n340 VDD.n339 0.120292
R4665 VDD.n341 VDD.n340 0.120292
R4666 VDD.n341 VDD.n202 0.120292
R4667 VDD.n351 VDD.n202 0.120292
R4668 VDD.n352 VDD.n351 0.120292
R4669 VDD.n354 VDD.n352 0.120292
R4670 VDD.n354 VDD.n353 0.120292
R4671 VDD.n353 VDD.n197 0.120292
R4672 VDD.n365 VDD.n197 0.120292
R4673 VDD.n366 VDD.n365 0.120292
R4674 VDD.n366 VDD.n190 0.120292
R4675 VDD.n373 VDD.n190 0.120292
R4676 VDD.n374 VDD.n373 0.120292
R4677 VDD.n375 VDD.n374 0.120292
R4678 VDD.n392 VDD.n375 0.120292
R4679 VDD.n392 VDD.n391 0.120292
R4680 VDD.n391 VDD.n388 0.120292
R4681 VDD.n388 VDD.n184 0.120292
R4682 VDD.n404 VDD.n184 0.120292
R4683 VDD.n405 VDD.n404 0.120292
R4684 VDD.n405 VDD.n178 0.120292
R4685 VDD.n414 VDD.n178 0.120292
R4686 VDD.n417 VDD.n414 0.120292
R4687 VDD.n419 VDD.n417 0.120292
R4688 VDD.n429 VDD.n428 0.120292
R4689 VDD.n430 VDD.n429 0.120292
R4690 VDD.n430 VDD.n167 0.120292
R4691 VDD.n440 VDD.n167 0.120292
R4692 VDD.n441 VDD.n440 0.120292
R4693 VDD.n443 VDD.n441 0.120292
R4694 VDD.n443 VDD.n442 0.120292
R4695 VDD.n442 VDD.n162 0.120292
R4696 VDD.n454 VDD.n162 0.120292
R4697 VDD.n455 VDD.n454 0.120292
R4698 VDD.n455 VDD.n155 0.120292
R4699 VDD.n462 VDD.n155 0.120292
R4700 VDD.n463 VDD.n462 0.120292
R4701 VDD.n464 VDD.n463 0.120292
R4702 VDD.n481 VDD.n464 0.120292
R4703 VDD.n481 VDD.n480 0.120292
R4704 VDD.n480 VDD.n477 0.120292
R4705 VDD.n477 VDD.n149 0.120292
R4706 VDD.n493 VDD.n149 0.120292
R4707 VDD.n494 VDD.n493 0.120292
R4708 VDD.n494 VDD.n143 0.120292
R4709 VDD.n503 VDD.n143 0.120292
R4710 VDD.n506 VDD.n503 0.120292
R4711 VDD.n508 VDD.n506 0.120292
R4712 VDD.n518 VDD.n517 0.120292
R4713 VDD.n519 VDD.n518 0.120292
R4714 VDD.n519 VDD.n132 0.120292
R4715 VDD.n529 VDD.n132 0.120292
R4716 VDD.n530 VDD.n529 0.120292
R4717 VDD.n532 VDD.n530 0.120292
R4718 VDD.n532 VDD.n531 0.120292
R4719 VDD.n531 VDD.n127 0.120292
R4720 VDD.n543 VDD.n127 0.120292
R4721 VDD.n544 VDD.n543 0.120292
R4722 VDD.n544 VDD.n120 0.120292
R4723 VDD.n551 VDD.n120 0.120292
R4724 VDD.n552 VDD.n551 0.120292
R4725 VDD.n553 VDD.n552 0.120292
R4726 VDD.n570 VDD.n553 0.120292
R4727 VDD.n570 VDD.n569 0.120292
R4728 VDD.n569 VDD.n566 0.120292
R4729 VDD.n566 VDD.n114 0.120292
R4730 VDD.n582 VDD.n114 0.120292
R4731 VDD.n584 VDD.n582 0.120292
R4732 VDD.n584 VDD.n583 0.120292
R4733 VDD.n583 VDD.n106 0.120292
R4734 VDD.n595 VDD.n106 0.120292
R4735 VDD.n596 VDD.n595 0.120292
R4736 VDD.n597 VDD.n99 0.120292
R4737 VDD.n608 VDD.n99 0.120292
R4738 VDD.n609 VDD.n608 0.120292
R4739 VDD.n610 VDD.n609 0.120292
R4740 VDD.n610 VDD.n91 0.120292
R4741 VDD.n622 VDD.n91 0.120292
R4742 VDD.n623 VDD.n622 0.120292
R4743 VDD.n624 VDD.n623 0.120292
R4744 VDD.n624 VDD.n83 0.120292
R4745 VDD.n637 VDD.n83 0.120292
R4746 VDD.n638 VDD.n637 0.120292
R4747 VDD.n742 VDD.n741 0.120292
R4748 VDD.n743 VDD.n742 0.120292
R4749 VDD.n744 VDD.n743 0.120292
R4750 VDD.n744 VDD.n18 0.120292
R4751 VDD.n755 VDD.n18 0.120292
R4752 VDD.n756 VDD.n12 0.120292
R4753 VDD.n764 VDD.n12 0.120292
R4754 VDD.n2682 VDD.n2678 0.120292
R4755 VDD.n2686 VDD.n2682 0.120292
R4756 VDD.n2692 VDD.n2686 0.120292
R4757 VDD.n2696 VDD.n2692 0.120292
R4758 VDD.n2701 VDD.n2696 0.120292
R4759 VDD.n2705 VDD.n2701 0.120292
R4760 VDD.n2709 VDD.n2705 0.120292
R4761 VDD.n2715 VDD.n2709 0.120292
R4762 VDD.n2719 VDD.n2715 0.120292
R4763 VDD.n2723 VDD.n2719 0.120292
R4764 VDD.n2726 VDD.n2723 0.120292
R4765 VDD.n2730 VDD.n2726 0.120292
R4766 VDD.n2734 VDD.n2730 0.120292
R4767 VDD.n2740 VDD.n2734 0.120292
R4768 VDD.n2744 VDD.n2740 0.120292
R4769 VDD.n2769 VDD.n2765 0.120292
R4770 VDD.n2773 VDD.n2769 0.120292
R4771 VDD.n2777 VDD.n2773 0.120292
R4772 VDD.n2782 VDD.n2777 0.120292
R4773 VDD.n2786 VDD.n2782 0.120292
R4774 VDD.n2788 VDD.n2786 0.120292
R4775 VDD.n2788 VDD.n2787 0.120292
R4776 VDD.n2799 VDD.n2669 0.120292
R4777 VDD.n2669 VDD.n2663 0.120292
R4778 VDD.n2663 VDD.n2659 0.120292
R4779 VDD.n2659 VDD.n2655 0.120292
R4780 VDD.n2655 VDD.n2649 0.120292
R4781 VDD.n2649 VDD.n2645 0.120292
R4782 VDD.n2645 VDD.n2640 0.120292
R4783 VDD.n2640 VDD.n2636 0.120292
R4784 VDD.n2636 VDD.n2632 0.120292
R4785 VDD.n2632 VDD.n2626 0.120292
R4786 VDD.n2626 VDD.n2622 0.120292
R4787 VDD.n2622 VDD.n2618 0.120292
R4788 VDD.n2618 VDD.n2615 0.120292
R4789 VDD.n2615 VDD.n2611 0.120292
R4790 VDD.n2611 VDD.n2607 0.120292
R4791 VDD.n2607 VDD.n2601 0.120292
R4792 VDD.n2580 VDD.n2576 0.120292
R4793 VDD.n2576 VDD.n2572 0.120292
R4794 VDD.n2572 VDD.n2568 0.120292
R4795 VDD.n2568 VDD.n2564 0.120292
R4796 VDD.n2564 VDD.n2559 0.120292
R4797 VDD.n2559 VDD.n2555 0.120292
R4798 VDD.n2555 VDD.n0 0.120292
R4799 VDD.n2546 VDD.n2545 0.120292
R4800 VDD.n2545 VDD.n2539 0.120292
R4801 VDD.n2539 VDD.n2535 0.120292
R4802 VDD.n2535 VDD.n2531 0.120292
R4803 VDD.n2531 VDD.n2525 0.120292
R4804 VDD.n2525 VDD.n2521 0.120292
R4805 VDD.n2521 VDD.n2516 0.120292
R4806 VDD.n2516 VDD.n2512 0.120292
R4807 VDD.n2512 VDD.n2508 0.120292
R4808 VDD.n2508 VDD.n2502 0.120292
R4809 VDD.n2502 VDD.n2498 0.120292
R4810 VDD.n2498 VDD.n2494 0.120292
R4811 VDD.n2494 VDD.n2491 0.120292
R4812 VDD.n2491 VDD.n2487 0.120292
R4813 VDD.n2487 VDD.n2483 0.120292
R4814 VDD.n2483 VDD.n2477 0.120292
R4815 VDD.n2456 VDD.n2452 0.120292
R4816 VDD.n2452 VDD.n2448 0.120292
R4817 VDD.n2448 VDD.n2444 0.120292
R4818 VDD.n2444 VDD.n2440 0.120292
R4819 VDD.n2440 VDD.n2435 0.120292
R4820 VDD.n2435 VDD.n2431 0.120292
R4821 VDD.n2431 VDD.n4 0.120292
R4822 VDD.n2422 VDD.n2421 0.120292
R4823 VDD.n2421 VDD.n2415 0.120292
R4824 VDD.n2415 VDD.n2411 0.120292
R4825 VDD.n2411 VDD.n2407 0.120292
R4826 VDD.n2407 VDD.n2401 0.120292
R4827 VDD.n2401 VDD.n2397 0.120292
R4828 VDD.n2397 VDD.n2392 0.120292
R4829 VDD.n2392 VDD.n2388 0.120292
R4830 VDD.n2388 VDD.n2384 0.120292
R4831 VDD.n2384 VDD.n2378 0.120292
R4832 VDD.n2378 VDD.n2374 0.120292
R4833 VDD.n2374 VDD.n2370 0.120292
R4834 VDD.n2370 VDD.n2367 0.120292
R4835 VDD.n2367 VDD.n2363 0.120292
R4836 VDD.n2363 VDD.n2359 0.120292
R4837 VDD.n2359 VDD.n2353 0.120292
R4838 VDD.n2332 VDD.n2328 0.120292
R4839 VDD.n2328 VDD.n2324 0.120292
R4840 VDD.n2324 VDD.n2320 0.120292
R4841 VDD.n2320 VDD.n2316 0.120292
R4842 VDD.n2316 VDD.n2311 0.120292
R4843 VDD.n2299 VDD.n8 0.120292
R4844 VDD.n2290 VDD.n2289 0.120292
R4845 VDD.n2289 VDD.n2283 0.120292
R4846 VDD.n2283 VDD.n2279 0.120292
R4847 VDD.n2279 VDD.n2275 0.120292
R4848 VDD.n2263 VDD.n2258 0.120292
R4849 VDD.n2258 VDD.n2254 0.120292
R4850 VDD.n2254 VDD.n2250 0.120292
R4851 VDD.n2250 VDD.n2244 0.120292
R4852 VDD.n2244 VDD.n2240 0.120292
R4853 VDD.n2240 VDD.n2236 0.120292
R4854 VDD.n2236 VDD.n2233 0.120292
R4855 VDD.n2233 VDD.n2229 0.120292
R4856 VDD.n2229 VDD.n2225 0.120292
R4857 VDD.n2225 VDD.n2219 0.120292
R4858 VDD.n2219 VDD.n2215 0.120292
R4859 VDD.n2215 VDD.n2211 0.120292
R4860 VDD.n2211 VDD.n2205 0.120292
R4861 VDD.n2205 VDD.n2201 0.120292
R4862 VDD.n2201 VDD.n2197 0.120292
R4863 VDD.n2197 VDD.n2193 0.120292
R4864 VDD.n2193 VDD.n2188 0.120292
R4865 VDD.n2188 VDD.n2184 0.120292
R4866 VDD.n2184 VDD.n2175 0.120292
R4867 VDD VDD.n2174 0.119505
R4868 VDD.n2044 VDD 0.119303
R4869 VDD.n2264 VDD.n2263 0.117688
R4870 VDD.n2765 VDD.n2761 0.111177
R4871 VDD.n2581 VDD.n2580 0.111177
R4872 VDD.n2457 VDD.n2456 0.111177
R4873 VDD.n2333 VDD.n2332 0.111177
R4874 VDD.n1303 VDD.n1302 0.108573
R4875 VDD.n638 VDD.n79 0.107271
R4876 VDD.n2745 VDD.n2744 0.107271
R4877 VDD.n2601 VDD.n2597 0.107271
R4878 VDD.n2477 VDD.n2473 0.107271
R4879 VDD.n2353 VDD.n2349 0.107271
R4880 VDD.n2045 VDD 0.104922
R4881 VDD.n2275 VDD.n2271 0.10076
R4882 VDD.n1308 VDD.n1307 0.0981562
R4883 VDD.n1320 VDD.n1318 0.0981562
R4884 VDD.n1330 VDD.n890 0.0981562
R4885 VDD.n1332 VDD.n886 0.0981562
R4886 VDD.n1345 VDD.n1343 0.0981562
R4887 VDD.n1359 VDD.n876 0.0981562
R4888 VDD.n1361 VDD.n872 0.0981562
R4889 VDD.n1375 VDD.n1372 0.0981562
R4890 VDD.n1373 VDD.n864 0.0981562
R4891 VDD.n1396 VDD.n858 0.0981562
R4892 VDD.n1398 VDD.n854 0.0981562
R4893 VDD.n1412 VDD.n1409 0.0981562
R4894 VDD.n1410 VDD.n845 0.0981562
R4895 VDD.n1428 VDD.n1425 0.0981562
R4896 VDD.n1426 VDD.n836 0.0981562
R4897 VDD.n835 VDD.n829 0.0981562
R4898 VDD.n651 VDD.n650 0.0981562
R4899 VDD.n664 VDD.n662 0.0981562
R4900 VDD.n674 VDD.n61 0.0981562
R4901 VDD.n676 VDD.n56 0.0981562
R4902 VDD.n689 VDD.n688 0.0981562
R4903 VDD.n702 VDD.n700 0.0981562
R4904 VDD.n712 VDD.n39 0.0981562
R4905 VDD.n714 VDD.n34 0.0981562
R4906 VDD.n730 VDD.n726 0.0981562
R4907 VDD.n2300 VDD.n2299 0.0981562
R4908 VDD.n2094 VDD 0.0968542
R4909 VDD.n1670 VDD 0.0968542
R4910 VDD.n1741 VDD 0.0968542
R4911 VDD.n1823 VDD 0.0968542
R4912 VDD.n1894 VDD 0.0968542
R4913 VDD.n1976 VDD 0.0968542
R4914 VDD.n250 VDD 0.0968542
R4915 VDD.n339 VDD 0.0968542
R4916 VDD.n428 VDD 0.0968542
R4917 VDD.n517 VDD 0.0968542
R4918 VDD.n292 VDD 0.0821977
R4919 VDD.n381 VDD 0.0821977
R4920 VDD.n470 VDD 0.0821977
R4921 VDD.n559 VDD 0.0821977
R4922 VDD.n292 VDD.n291 0.0783056
R4923 VDD.n381 VDD.n380 0.0783056
R4924 VDD.n470 VDD.n469 0.0783056
R4925 VDD.n559 VDD.n558 0.0783056
R4926 VDD.n2750 VDD.n2749 0.076587
R4927 VDD.n2586 VDD.n2585 0.076587
R4928 VDD.n2462 VDD.n2461 0.076587
R4929 VDD.n2338 VDD.n2337 0.076587
R4930 VDD VDD.n2148 0.0603958
R4931 VDD VDD.n2164 0.0603958
R4932 VDD.n2165 VDD 0.0603958
R4933 VDD VDD.n1739 0.0603958
R4934 VDD.n1740 VDD 0.0603958
R4935 VDD.n1814 VDD 0.0603958
R4936 VDD VDD.n1813 0.0603958
R4937 VDD VDD.n1892 0.0603958
R4938 VDD.n1893 VDD 0.0603958
R4939 VDD.n1967 VDD 0.0603958
R4940 VDD VDD.n1966 0.0603958
R4941 VDD VDD.n2043 0.0603958
R4942 VDD.n1115 VDD 0.0603958
R4943 VDD.n1191 VDD 0.0603958
R4944 VDD.n1273 VDD 0.0603958
R4945 VDD.n330 VDD 0.0603958
R4946 VDD VDD.n329 0.0603958
R4947 VDD.n419 VDD 0.0603958
R4948 VDD VDD.n418 0.0603958
R4949 VDD.n508 VDD 0.0603958
R4950 VDD VDD.n507 0.0603958
R4951 VDD VDD.n596 0.0603958
R4952 VDD.n597 VDD 0.0603958
R4953 VDD VDD.n755 0.0603958
R4954 VDD.n756 VDD 0.0603958
R4955 VDD VDD.n764 0.0603958
R4956 VDD VDD.n2799 0.0603958
R4957 VDD.n2546 VDD 0.0603958
R4958 VDD.n2422 VDD 0.0603958
R4959 VDD.n2290 VDD 0.0603958
R4960 VDD.n797 VDD.n775 0.0505
R4961 VDD.n809 VDD.n775 0.0505
R4962 VDD.n789 VDD.n788 0.0483261
R4963 VDD.n2752 VDD.n2751 0.0439783
R4964 VDD.n2588 VDD.n2587 0.0439783
R4965 VDD.n2464 VDD.n2463 0.0439783
R4966 VDD.n2340 VDD.n2339 0.0439783
R4967 VDD.n822 VDD.n768 0.0414968
R4968 VDD.n794 VDD.n793 0.0396302
R4969 VDD.n797 VDD.n796 0.0395981
R4970 VDD.n813 VDD.n812 0.0359398
R4971 VDD.n2751 VDD 0.0358261
R4972 VDD.n2587 VDD 0.0358261
R4973 VDD.n2463 VDD 0.0358261
R4974 VDD.n2339 VDD 0.0358261
R4975 VDD.n1452 VDD 0.0356562
R4976 VDD.n741 VDD 0.0343542
R4977 VDD VDD.n1740 0.0239375
R4978 VDD.n1813 VDD 0.0239375
R4979 VDD VDD.n1893 0.0239375
R4980 VDD.n1966 VDD 0.0239375
R4981 VDD.n329 VDD 0.0239375
R4982 VDD.n418 VDD 0.0239375
R4983 VDD.n507 VDD 0.0239375
R4984 VDD VDD.n2173 0.0226354
R4985 VDD VDD.n1460 0.0226354
R4986 VDD.n2311 VDD.n2300 0.0226354
R4987 VDD.n1103 VDD 0.0213333
R4988 VDD VDD.n1190 0.0213333
R4989 VDD.n1261 VDD 0.0213333
R4990 VDD.n2787 VDD 0.0213333
R4991 VDD VDD.n0 0.0213333
R4992 VDD VDD.n4 0.0213333
R4993 VDD VDD.n8 0.0213333
R4994 VDD.n2175 VDD 0.0213333
R4995 VDD.n2271 VDD.n2270 0.0200312
R4996 VDD.n810 VDD 0.0195217
R4997 VDD.n79 VDD.n76 0.0135208
R4998 VDD.n651 VDD.n69 0.0135208
R4999 VDD.n664 VDD.n663 0.0135208
R5000 VDD.n675 VDD.n674 0.0135208
R5001 VDD.n56 VDD.n54 0.0135208
R5002 VDD.n689 VDD.n47 0.0135208
R5003 VDD.n702 VDD.n701 0.0135208
R5004 VDD.n713 VDD.n712 0.0135208
R5005 VDD.n34 VDD.n32 0.0135208
R5006 VDD.n730 VDD.n729 0.0135208
R5007 VDD.n2760 VDD.n2745 0.0135208
R5008 VDD.n2597 VDD.n2596 0.0135208
R5009 VDD.n2473 VDD.n2472 0.0135208
R5010 VDD.n2349 VDD.n2348 0.0135208
R5011 VDD.n812 VDD.n811 0.0135
R5012 VDD.n796 VDD.n795 0.0123444
R5013 VDD.n1303 VDD.n904 0.0122188
R5014 VDD.n1308 VDD.n898 0.0122188
R5015 VDD.n1320 VDD.n1319 0.0122188
R5016 VDD.n1331 VDD.n1330 0.0122188
R5017 VDD.n886 VDD.n884 0.0122188
R5018 VDD.n1345 VDD.n1344 0.0122188
R5019 VDD.n1360 VDD.n1359 0.0122188
R5020 VDD.n872 VDD.n870 0.0122188
R5021 VDD.n1375 VDD.n1374 0.0122188
R5022 VDD.n1384 VDD.n864 0.0122188
R5023 VDD.n1397 VDD.n1396 0.0122188
R5024 VDD.n854 VDD.n852 0.0122188
R5025 VDD.n1412 VDD.n1411 0.0122188
R5026 VDD.n845 VDD.n842 0.0122188
R5027 VDD.n1428 VDD.n1427 0.0122188
R5028 VDD.n1437 VDD.n836 0.0122188
R5029 VDD.n1450 VDD.n829 0.0122188
R5030 VDD.n727 VDD 0.0122188
R5031 VDD.n2048 VDD.n2047 0.0114224
R5032 VDD.n1307 VDD.n904 0.0109167
R5033 VDD.n1318 VDD.n898 0.0109167
R5034 VDD.n1319 VDD.n890 0.0109167
R5035 VDD.n1332 VDD.n1331 0.0109167
R5036 VDD.n1343 VDD.n884 0.0109167
R5037 VDD.n1344 VDD.n876 0.0109167
R5038 VDD.n1361 VDD.n1360 0.0109167
R5039 VDD.n1372 VDD.n870 0.0109167
R5040 VDD.n1374 VDD.n1373 0.0109167
R5041 VDD.n1384 VDD.n858 0.0109167
R5042 VDD.n1398 VDD.n1397 0.0109167
R5043 VDD.n1409 VDD.n852 0.0109167
R5044 VDD.n1411 VDD.n1410 0.0109167
R5045 VDD.n1425 VDD.n842 0.0109167
R5046 VDD.n1427 VDD.n1426 0.0109167
R5047 VDD.n1437 VDD.n835 0.0109167
R5048 VDD.n1451 VDD.n1450 0.0109167
R5049 VDD VDD.n1451 0.0109167
R5050 VDD.n811 VDD.n768 0.0104632
R5051 VDD VDD.n822 0.00973913
R5052 VDD.n650 VDD.n76 0.00961458
R5053 VDD.n662 VDD.n69 0.00961458
R5054 VDD.n663 VDD.n61 0.00961458
R5055 VDD.n676 VDD.n675 0.00961458
R5056 VDD.n688 VDD.n54 0.00961458
R5057 VDD.n700 VDD.n47 0.00961458
R5058 VDD.n701 VDD.n39 0.00961458
R5059 VDD.n714 VDD.n713 0.00961458
R5060 VDD.n726 VDD.n32 0.00961458
R5061 VDD.n729 VDD.n727 0.00961458
R5062 VDD.n2761 VDD.n2760 0.00961458
R5063 VDD.n2596 VDD.n2581 0.00961458
R5064 VDD.n2472 VDD.n2457 0.00961458
R5065 VDD.n2348 VDD.n2333 0.00961458
R5066 VDD.n2174 VDD.n2048 0.0093414
R5067 VDD VDD.n809 0.00919565
R5068 VDD.n793 VDD.n783 0.00756522
R5069 VDD.n814 VDD.n810 0.00647826
R5070 VDD.n795 VDD.n794 0.00589131
R5071 VDD.n814 VDD.n813 0.00376087
R5072 VDD.n2752 VDD.n2750 0.00321739
R5073 VDD.n2588 VDD.n2586 0.00321739
R5074 VDD.n2464 VDD.n2462 0.00321739
R5075 VDD.n2340 VDD.n2338 0.00321739
R5076 VDD.n2270 VDD.n2264 0.00310417
R5077 VDD.n789 VDD.n783 0.00267391
R5078 VDD.n2174 VDD 0.00195147
R5079 VDD.n812 VDD.n766 0.0010004
R5080 VDD.n794 VDD.n767 0.0010004
R5081 VDD.n2047 VDD.n765 0.001
R5082 VDD.n2045 VDD.n2044 0.000604271
R5083 VDD.n2047 VDD.n2046 0.000552135
R5084 VDD.n2046 VDD.n2045 0.000552135
R5085 VDD.n2044 VDD.n1461 0.000501704
R5086 VDD.n2046 VDD.n767 0.000501351
R5087 VDD.n2046 VDD.n766 0.000501351
R5088 check[1].n3 check[1].t5 331.51
R5089 check[1].n1 check[1].t2 280.899
R5090 check[1].n1 check[1].t3 216.238
R5091 check[1].n3 check[1].t4 209.403
R5092 check[1].n0 check[1].t1 207.373
R5093 check[1].n4 check[1].n3 76.0005
R5094 check[1].n7 check[1].n6 50.467
R5095 check[1].n2 check[1].n1 35.7166
R5096 check[1].n8 check[1].t0 33.1309
R5097 check[1].n5 check[1].n2 32.9012
R5098 check[1].n7 check[1] 15.9389
R5099 check[1].n6 check[1] 12.062
R5100 check[1] check[1].n0 9.01934
R5101 check[1].n5 check[1] 8.68932
R5102 check[1] check[1].n4 8.58587
R5103 check[1] check[1].n8 8.00801
R5104 check[1].n0 check[1] 7.45876
R5105 check[1].n6 check[1].n5 3.04357
R5106 check[1].n2 check[1] 2.56973
R5107 check[1].n4 check[1] 2.02977
R5108 check[1].n8 check[1].n7 1.94232
R5109 D[0].n8 D[0].t2 269.921
R5110 D[0].n8 D[0].t3 234.573
R5111 D[0].n7 D[0].t1 207.373
R5112 D[0].n9 D[0].n8 76.0005
R5113 D[0].n14 D[0].t0 33.3405
R5114 D[0].n12 D[0].n11 26.2261
R5115 D[0].n11 D[0] 19.418
R5116 D[0].n11 D[0].n10 14.9338
R5117 D[0] D[0].n14 9.32876
R5118 D[0] D[0].n7 9.01934
R5119 D[0].n7 D[0] 7.45876
R5120 D[0].n3 D[0] 6.42
R5121 D[0].n10 D[0] 5.9498
R5122 D[0].n9 D[0] 4.68782
R5123 D[0].n13 D[0].n12 3.50069
R5124 D[0].n12 D[0].n6 2.83165
R5125 D[0].n5 D[0].n1 2.26284
R5126 D[0].n4 D[0].n3 2.23869
R5127 D[0].n10 D[0].n9 1.62304
R5128 D[0].n14 D[0].n13 0.391757
R5129 D[0].n4 D[0].n2 0.0213333
R5130 D[0].n6 D[0].n0 0.0099697
R5131 D[0].n5 D[0].n4 0.00195195
R5132 D[0].n6 D[0].n5 0.00194159
R5133 eob.n10 eob.t11 331.51
R5134 eob.n4 eob 298.998
R5135 eob.n5 eob.n4 292.5
R5136 eob.n0 eob.t8 230.576
R5137 eob.n10 eob.t10 209.403
R5138 eob.n3 eob.n1 180.082
R5139 eob.n0 eob.t9 158.275
R5140 eob.n3 eob.n2 124.501
R5141 eob.n8 eob.n7 92.5005
R5142 eob eob.n0 82.6672
R5143 eob.n11 eob.n10 76.0005
R5144 eob.n6 eob.n3 36.0005
R5145 eob.n4 eob.t1 26.5955
R5146 eob.n4 eob.t3 26.5955
R5147 eob.n1 eob.t4 26.5955
R5148 eob.n1 eob.t2 26.5955
R5149 eob eob.n13 25.8571
R5150 eob.n7 eob.t0 24.9236
R5151 eob.n7 eob.t6 24.9236
R5152 eob.n2 eob.t7 24.9236
R5153 eob.n2 eob.t5 24.9236
R5154 eob.n12 eob.n9 11.9351
R5155 eob.n12 eob 11.6575
R5156 eob.n6 eob 10.2405
R5157 eob.n13 eob.n12 9.41338
R5158 eob eob.n11 8.58587
R5159 eob eob.n5 8.46819
R5160 eob eob.n8 8.07435
R5161 eob.n13 eob 7.22276
R5162 eob.n8 eob 5.31742
R5163 eob.n5 eob 4.92358
R5164 eob.n9 eob 2.95435
R5165 eob.n11 eob 2.02977
R5166 eob.n9 eob.n6 0.197423
R5167 VSS.n4169 VSS 52235.6
R5168 VSS.n3888 VSS.n3433 7556.59
R5169 VSS.n3433 VSS.n55 6484.98
R5170 VSS VSS.n3888 5751.89
R5171 VSS.n1994 VSS.n1991 2560.8
R5172 VSS.n1404 VSS.n1403 2487.33
R5173 VSS.n1482 VSS.n55 2302.75
R5174 VSS.n3433 VSS 1640.08
R5175 VSS.n4170 VSS.n4169 1234.15
R5176 VSS.n3888 VSS 1073.17
R5177 VSS.n4284 VSS 1019.51
R5178 VSS.n3544 VSS 1019.51
R5179 VSS.n3658 VSS 1019.51
R5180 VSS.n3772 VSS 1019.51
R5181 VSS.n3378 VSS.n3377 721.875
R5182 VSS.n3419 VSS 670.14
R5183 VSS.n3377 VSS.t658 653.125
R5184 VSS VSS.n3902 651.852
R5185 VSS VSS.t588 630.489
R5186 VSS VSS.t414 630.489
R5187 VSS VSS.t416 630.489
R5188 VSS VSS.t63 630.489
R5189 VSS.t642 VSS 630.489
R5190 VSS.n4259 VSS.t263 603.659
R5191 VSS.n3519 VSS.t652 603.659
R5192 VSS.n3633 VSS.t686 603.659
R5193 VSS.n3747 VSS.t277 603.659
R5194 VSS.n3861 VSS.t479 603.659
R5195 VSS.n4174 VSS.t436 590.245
R5196 VSS.n4267 VSS.t668 590.245
R5197 VSS.t588 VSS.n4280 590.245
R5198 VSS.n1 VSS.t220 590.245
R5199 VSS.n3527 VSS.t422 590.245
R5200 VSS.t414 VSS.n3542 590.245
R5201 VSS.n3548 VSS.t430 590.245
R5202 VSS.n3641 VSS.t77 590.245
R5203 VSS.t416 VSS.n3656 590.245
R5204 VSS.n3662 VSS.t666 590.245
R5205 VSS.n3755 VSS.t578 590.245
R5206 VSS.t63 VSS.n3770 590.245
R5207 VSS.n3776 VSS.t664 590.245
R5208 VSS.n3869 VSS.t396 590.245
R5209 VSS.n3878 VSS.t642 590.245
R5210 VSS.n74 VSS.t662 584.375
R5211 VSS VSS.n3333 574.659
R5212 VSS.n4180 VSS.t245 550
R5213 VSS.n3440 VSS.t308 550
R5214 VSS.n3554 VSS.t290 550
R5215 VSS.n3668 VSS.t109 550
R5216 VSS.n3782 VSS.t208 550
R5217 VSS.n4280 VSS.t265 536.586
R5218 VSS.n3542 VSS.t654 536.586
R5219 VSS.n3656 VSS.t684 536.586
R5220 VSS.n3770 VSS.t275 536.586
R5221 VSS.n3878 VSS.t481 536.586
R5222 VSS.n3420 VSS.n3417 533.059
R5223 VSS.n3904 VSS.n3901 533.059
R5224 VSS.n3376 VSS.n75 533.059
R5225 VSS.n3353 VSS.n3349 533.059
R5226 VSS.n3349 VSS.n3338 533.059
R5227 VSS.n3545 VSS.n3438 533.059
R5228 VSS.n3659 VSS.n3436 533.059
R5229 VSS.n3773 VSS.n3434 533.059
R5230 VSS.n4206 VSS.t52 509.757
R5231 VSS.n3466 VSS.t599 509.757
R5232 VSS.n3580 VSS.t598 509.757
R5233 VSS.n3694 VSS.t239 509.757
R5234 VSS.n3808 VSS.t624 509.757
R5235 VSS.n4188 VSS.t241 496.341
R5236 VSS.n3448 VSS.t310 496.341
R5237 VSS.n3562 VSS.t292 496.341
R5238 VSS.n3676 VSS.t111 496.341
R5239 VSS.n3790 VSS.t204 496.341
R5240 VSS.n3394 VSS 493.788
R5241 VSS.n285 VSS 488.889
R5242 VSS.n286 VSS.n281 475.118
R5243 VSS.n4194 VSS.t14 456.099
R5244 VSS.n3454 VSS.t117 456.099
R5245 VSS.n3568 VSS.t18 456.099
R5246 VSS.n3682 VSS.t271 456.099
R5247 VSS.n3796 VSS.t159 456.099
R5248 VSS.n917 VSS.n916 434.56
R5249 VSS.n599 VSS.n598 434.56
R5250 VSS VSS.n1219 428.851
R5251 VSS.n919 VSS 428.851
R5252 VSS.n601 VSS 428.851
R5253 VSS.n4255 VSS.t126 415.854
R5254 VSS.n3515 VSS.t462 415.854
R5255 VSS.n3629 VSS.t384 415.854
R5256 VSS.n3743 VSS.t478 415.854
R5257 VSS.n3857 VSS.t670 415.854
R5258 VSS.n4202 VSS.t446 402.44
R5259 VSS.n3462 VSS.t136 402.44
R5260 VSS.n3576 VSS.t513 402.44
R5261 VSS.n3690 VSS.t400 402.44
R5262 VSS.n3804 VSS.t506 402.44
R5263 VSS.n2014 VSS.t5 396
R5264 VSS.n2129 VSS.t321 396
R5265 VSS.n3411 VSS.t621 387.976
R5266 VSS.n3423 VSS.t192 387.976
R5267 VSS.n3423 VSS.t216 387.976
R5268 VSS.n1995 VSS.t65 387.2
R5269 VSS.n2005 VSS.t81 387.2
R5270 VSS.n2097 VSS.t8 387.2
R5271 VSS.n2110 VSS.t137 387.2
R5272 VSS.n2120 VSS.t87 387.2
R5273 VSS.n2271 VSS.t632 387.2
R5274 VSS.n2623 VSS.t371 387.2
R5275 VSS.n2975 VSS.t373 387.2
R5276 VSS VSS.n3351 383.486
R5277 VSS.n1221 VSS.n135 382.413
R5278 VSS.n3909 VSS.t523 377.389
R5279 VSS.n3893 VSS.t525 377.389
R5280 VSS.n3893 VSS.t0 377.389
R5281 VSS.n123 VSS.t602 377.389
R5282 VSS.n3984 VSS.t394 368.812
R5283 VSS.n3955 VSS.t388 368.812
R5284 VSS.n4251 VSS.t509 362.195
R5285 VSS.n3511 VSS.t452 362.195
R5286 VSS.n3625 VSS.t299 362.195
R5287 VSS.n3739 VSS.t547 362.195
R5288 VSS.n3853 VSS.t367 362.195
R5289 VSS.n2093 VSS.t438 360.8
R5290 VSS.n4013 VSS.t576 360.235
R5291 VSS.n3411 VSS.t563 352.705
R5292 VSS.n1995 VSS.t2 352
R5293 VSS.n2110 VSS.t319 352
R5294 VSS.n2243 VSS.t420 352
R5295 VSS.n2595 VSS.t120 352
R5296 VSS.n2947 VSS.t218 352
R5297 VSS.n1398 VSS.t251 351.658
R5298 VSS.n3358 VSS.t660 343.75
R5299 VSS.n3909 VSS.t180 343.08
R5300 VSS.n985 VSS.t647 343.08
R5301 VSS.n667 VSS.t255 343.08
R5302 VSS.n349 VSS.t323 343.08
R5303 VSS.n4027 VSS.t645 334.503
R5304 VSS.n2067 VSS.t240 334.401
R5305 VSS.n3063 VSS.t325 334.401
R5306 VSS.n262 VSS.t693 327.046
R5307 VSS.n1377 VSS.t253 325.926
R5308 VSS.n2083 VSS.t442 325.601
R5309 VSS.n128 VSS.t247 317.349
R5310 VSS.n1001 VSS.t426 308.772
R5311 VSS.n683 VSS.t472 308.772
R5312 VSS.n365 VSS.t83 308.772
R5313 VSS.n2079 VSS.t428 299.2
R5314 VSS.n3942 VSS.n3941 292.5
R5315 VSS.n3941 VSS.n3940 292.5
R5316 VSS.n3939 VSS.n3938 292.5
R5317 VSS.n3938 VSS.n3937 292.5
R5318 VSS.n3936 VSS.n3935 292.5
R5319 VSS.n3935 VSS.n3934 292.5
R5320 VSS.n3933 VSS.n3932 292.5
R5321 VSS.n3932 VSS.n3931 292.5
R5322 VSS.n3930 VSS.n3929 292.5
R5323 VSS.n3929 VSS.n3928 292.5
R5324 VSS.n3341 VSS.n3340 292.5
R5325 VSS.n3340 VSS.n3339 292.5
R5326 VSS.n3349 VSS.n3348 292.5
R5327 VSS.n3351 VSS.n3349 292.5
R5328 VSS.n3354 VSS.n3353 292.5
R5329 VSS.n3353 VSS.n3352 292.5
R5330 VSS.n3360 VSS.n3359 292.5
R5331 VSS.n3359 VSS.n3358 292.5
R5332 VSS.n3364 VSS.n3363 292.5
R5333 VSS.n3363 VSS.n3362 292.5
R5334 VSS.n3370 VSS.n3369 292.5
R5335 VSS.n3369 VSS.n3368 292.5
R5336 VSS.n3376 VSS.n3375 292.5
R5337 VSS.n3377 VSS.n3376 292.5
R5338 VSS.n1389 VSS.t269 291.618
R5339 VSS.n3405 VSS.t561 282.164
R5340 VSS.n3362 VSS.t656 275
R5341 VSS.n3913 VSS.t176 274.464
R5342 VSS.n2018 VSS.t475 272.8
R5343 VSS.n2133 VSS.t191 272.8
R5344 VSS.n1281 VSS.t493 265.887
R5345 VSS.t65 VSS 264
R5346 VSS.n2071 VSS.t261 264
R5347 VSS.t137 VSS 264
R5348 VSS.t596 VSS 264
R5349 VSS.t139 VSS 264
R5350 VSS.n3077 VSS.t337 264
R5351 VSS.n269 VSS.t692 260.281
R5352 VSS VSS.t381 257.31
R5353 VSS.n1381 VSS.t557 257.31
R5354 VSS.n2199 VSS.t24 246.4
R5355 VSS.n2296 VSS.t20 246.4
R5356 VSS.n2551 VSS.t410 246.4
R5357 VSS.n2648 VSS.t412 246.4
R5358 VSS.n2903 VSS.t519 246.4
R5359 VSS.n3000 VSS.t515 246.4
R5360 VSS.n3351 VSS.t569 242.202
R5361 VSS.n3352 VSS.t432 242.202
R5362 VSS.n4216 VSS.t243 241.464
R5363 VSS.n3476 VSS.t306 241.464
R5364 VSS.n3590 VSS.t288 241.464
R5365 VSS.n3704 VSS.t107 241.464
R5366 VSS.n3818 VSS.t206 241.464
R5367 VSS.n2024 VSS.t361 237.601
R5368 VSS.n2139 VSS.t258 237.601
R5369 VSS.n2241 VSS.t67 237.601
R5370 VSS.n2593 VSS.t623 237.601
R5371 VSS.n2945 VSS.t634 237.601
R5372 VSS.n1965 VSS.t280 237.126
R5373 VSS.n1864 VSS.t501 237.126
R5374 VSS.n1763 VSS.t298 237.126
R5375 VSS.n1662 VSS.t201 237.126
R5376 VSS.n1561 VSS.t502 237.126
R5377 VSS.t273 VSS.n1983 231.857
R5378 VSS.n1408 VSS.t608 231.857
R5379 VSS.n1417 VSS.t70 231.857
R5380 VSS.t194 VSS.n1882 231.857
R5381 VSS.n1423 VSS.t614 231.857
R5382 VSS.n1432 VSS.t202 231.857
R5383 VSS.t379 VSS.n1781 231.857
R5384 VSS.n1438 VSS.t616 231.857
R5385 VSS.n1447 VSS.t312 231.857
R5386 VSS.t386 VSS.n1680 231.857
R5387 VSS.n1453 VSS.t610 231.857
R5388 VSS.n1462 VSS.t690 231.857
R5389 VSS.t594 VSS.n1579 231.857
R5390 VSS.n1468 VSS.t604 231.857
R5391 VSS.n1477 VSS.t636 231.857
R5392 VSS.n1293 VSS.t316 231.579
R5393 VSS.n271 VSS.t541 229.315
R5394 VSS VSS.n3393 229.26
R5395 VSS.t569 VSS.n3350 222.018
R5396 VSS.n3350 VSS.t567 222.018
R5397 VSS.n2185 VSS.t318 220
R5398 VSS.n2368 VSS.t640 220
R5399 VSS.n2537 VSS.t638 220
R5400 VSS.n2720 VSS.t72 220
R5401 VSS.n2889 VSS.t74 220
R5402 VSS.n1891 VSS.t466 216.048
R5403 VSS.n1790 VSS.t674 216.048
R5404 VSS.n1689 VSS.t210 216.048
R5405 VSS.n1588 VSS.t41 216.048
R5406 VSS.n1487 VSS.t555 216.048
R5407 VSS VSS.n4283 214.635
R5408 VSS VSS.n3543 214.635
R5409 VSS VSS.n3657 214.635
R5410 VSS VSS.n3771 214.635
R5411 VSS VSS.n3887 214.635
R5412 VSS.n3399 VSS.t565 211.624
R5413 VSS.n2322 VSS.t22 211.201
R5414 VSS.n2674 VSS.t408 211.201
R5415 VSS.n3026 VSS.t517 211.201
R5416 VSS.n1983 VSS.t281 210.779
R5417 VSS.n1882 VSS.t499 210.779
R5418 VSS.n1781 VSS.t295 210.779
R5419 VSS.n1680 VSS.t198 210.779
R5420 VSS.n1579 VSS.t503 210.779
R5421 VSS.n3982 VSS.t390 205.849
R5422 VSS.n3953 VSS.t392 205.849
R5423 VSS.n3917 VSS.t182 205.849
R5424 VSS.n4220 VSS.t264 201.22
R5425 VSS.n3480 VSS.t653 201.22
R5426 VSS.n3594 VSS.t687 201.22
R5427 VSS.n3708 VSS.t278 201.22
R5428 VSS.n3822 VSS.t480 201.22
R5429 VSS.n1912 VSS.t458 200.24
R5430 VSS.n1811 VSS.t383 200.24
R5431 VSS.n1710 VSS.t370 200.24
R5432 VSS.n1609 VSS.t10 200.24
R5433 VSS.n1508 VSS.t575 200.24
R5434 VSS.n260 VSS.t544 198.691
R5435 VSS.n1412 VSS.t464 194.97
R5436 VSS.n1427 VSS.t678 194.97
R5437 VSS.n1442 VSS.t214 194.97
R5438 VSS.n1457 VSS.t45 194.97
R5439 VSS.n1472 VSS.t553 194.97
R5440 VSS.n2215 VSS.t171 193.601
R5441 VSS.n2567 VSS.t167 193.601
R5442 VSS.n2919 VSS.t155 193.601
R5443 VSS.n2040 VSS.t364 190.337
R5444 VSS.n2155 VSS.t257 190.337
R5445 VSS.n2498 VSS.t651 190.337
R5446 VSS.n2850 VSS.t484 190.337
R5447 VSS.n415 VSS.t86 190.337
R5448 VSS.n733 VSS.t471 190.337
R5449 VSS.n1051 VSS.t425 190.337
R5450 VSS.n1327 VSS.t315 190.337
R5451 VSS.n1938 VSS.t451 190.337
R5452 VSS.n1837 VSS.t37 190.337
R5453 VSS.n1736 VSS.t104 190.337
R5454 VSS.n1635 VSS.t124 190.337
R5455 VSS.n1534 VSS.t223 190.337
R5456 VSS.n4232 VSS.t512 190.337
R5457 VSS.n3492 VSS.t455 190.337
R5458 VSS.n3606 VSS.t302 190.337
R5459 VSS.n3720 VSS.t550 190.337
R5460 VSS.n3834 VSS.t366 190.337
R5461 VSS.n3058 VSS.t326 190.065
R5462 VSS.n136 VSS.t495 188.695
R5463 VSS.n912 VSS.t672 188.695
R5464 VSS.n594 VSS.t11 188.695
R5465 VSS.n282 VSS.t542 188.695
R5466 VSS.n2338 VSS.t95 184.8
R5467 VSS.n2394 VSS.t227 184.8
R5468 VSS.n2690 VSS.t48 184.8
R5469 VSS.n2746 VSS.t406 184.8
R5470 VSS.n95 VSS.t127 184.8
R5471 VSS.n4157 VSS.t491 180.118
R5472 VSS.n4041 VSS.t586 180.118
R5473 VSS.n1257 VSS.t235 180.118
R5474 VSS.n955 VSS.t59 180.118
R5475 VSS.n637 VSS.t573 180.118
R5476 VSS.n319 VSS.t378 180.118
R5477 VSS.n1900 VSS.t28 179.162
R5478 VSS.n1799 VSS.t402 179.162
R5479 VSS.n1698 VSS.t404 179.162
R5480 VSS.n1597 VSS.t50 179.162
R5481 VSS.n1496 VSS.t26 179.162
R5482 VSS.n3379 VSS.t535 172.049
R5483 VSS.n1961 VSS.t79 163.353
R5484 VSS.n1860 VSS.t303 163.353
R5485 VSS.n1759 VSS.t97 163.353
R5486 VSS.n1658 VSS.t185 163.353
R5487 VSS.n1557 VSS.t197 163.353
R5488 VSS.n4212 VSS.t161 160.976
R5489 VSS.n3472 VSS.t151 160.976
R5490 VSS.n3586 VSS.t143 160.976
R5491 VSS.n3700 VSS.t173 160.976
R5492 VSS.n3814 VSS.t434 160.976
R5493 VSS.n2057 VSS.t440 158.4
R5494 VSS.n2408 VSS.t639 158.4
R5495 VSS.n2760 VSS.t75 158.4
R5496 VSS VSS.t273 158.084
R5497 VSS.n1908 VSS.t189 158.084
R5498 VSS VSS.t194 158.084
R5499 VSS.n1807 VSS.t522 158.084
R5500 VSS VSS.t379 158.084
R5501 VSS.n1706 VSS.t187 158.084
R5502 VSS VSS.t386 158.084
R5503 VSS.n1605 VSS.t100 158.084
R5504 VSS VSS.t594 158.084
R5505 VSS.n1504 VSS.t460 158.084
R5506 VSS.n4138 VSS.t644 154.387
R5507 VSS.n1367 VSS.t249 154.387
R5508 VSS.n1248 VSS.t612 154.387
R5509 VSS.n142 VSS.t625 154.387
R5510 VSS.n1043 VSS.t285 154.387
R5511 VSS.n1015 VSS.t489 154.387
R5512 VSS.n151 VSS.t606 154.387
R5513 VSS.n179 VSS.t444 154.387
R5514 VSS.n725 VSS.t585 154.387
R5515 VSS.n697 VSS.t233 154.387
R5516 VSS.n196 VSS.t618 154.387
R5517 VSS.n224 VSS.t68 154.387
R5518 VSS.n407 VSS.t601 154.387
R5519 VSS.n379 VSS.t630 154.387
R5520 VSS.n241 VSS.t545 154.387
R5521 VSS.n2355 VSS.t596 149.601
R5522 VSS.n2707 VSS.t139 149.601
R5523 VSS.n1350 VSS.n1349 145.81
R5524 VSS.n1340 VSS.n1339 145.81
R5525 VSS.n1330 VSS.n1329 145.81
R5526 VSS.n1320 VSS.n1319 145.81
R5527 VSS.n1310 VSS.n1309 145.81
R5528 VSS.n1300 VSS.n1299 145.81
R5529 VSS.n1290 VSS.n1289 145.81
R5530 VSS.n1278 VSS.n1277 145.81
R5531 VSS.n1268 VSS.n1267 145.81
R5532 VSS.n1258 VSS.n1257 145.81
R5533 VSS.n1249 VSS.n1248 145.81
R5534 VSS.n1238 VSS.n1237 145.81
R5535 VSS.n1228 VSS.n1227 145.81
R5536 VSS.n139 VSS.n136 145.81
R5537 VSS.n1219 VSS.n1218 145.81
R5538 VSS.n143 VSS.n142 145.81
R5539 VSS.n1204 VSS.n1203 145.81
R5540 VSS.n1194 VSS.n1193 145.81
R5541 VSS.n1184 VSS.n1183 145.81
R5542 VSS.n1173 VSS.n1172 145.81
R5543 VSS.n1163 VSS.n1162 145.81
R5544 VSS.n1153 VSS.n1152 145.81
R5545 VSS.n3334 VSS 145.81
R5546 VSS.n40 VSS.t230 145.303
R5547 VSS.n2008 VSS.t82 145.203
R5548 VSS.n2123 VSS.t88 145.203
R5549 VSS.n1253 VSS.t613 145.203
R5550 VSS.n1411 VSS.t609 145.203
R5551 VSS.n1426 VSS.t615 145.203
R5552 VSS.n1441 VSS.t617 145.203
R5553 VSS.n1456 VSS.t611 145.203
R5554 VSS.n1471 VSS.t605 145.203
R5555 VSS.n4270 VSS.t669 145.203
R5556 VSS.n3530 VSS.t423 145.203
R5557 VSS.n3644 VSS.t78 145.203
R5558 VSS.n3758 VSS.t579 145.203
R5559 VSS.n3872 VSS.t397 145.203
R5560 VSS.n2386 VSS.t228 144.49
R5561 VSS.n2738 VSS.t407 144.49
R5562 VSS.n249 VSS.t546 144.49
R5563 VSS.n204 VSS.t619 144.49
R5564 VSS.n159 VSS.t607 144.49
R5565 VSS.n1957 VSS.t448 142.275
R5566 VSS.n1856 VSS.t38 142.275
R5567 VSS.n1755 VSS.t101 142.275
R5568 VSS.n1654 VSS.t121 142.275
R5569 VSS.n1553 VSS.t224 142.275
R5570 VSS.n57 VSS.t559 141.083
R5571 VSS VSS.n3418 141.083
R5572 VSS.t658 VSS.n74 137.5
R5573 VSS.n51 VSS.t178 137.232
R5574 VSS.n3903 VSS 137.232
R5575 VSS.n1220 VSS 137.232
R5576 VSS.n3214 VSS.t343 133.816
R5577 VSS VSS.n3432 132.266
R5578 VSS.n2053 VSS.t4 132
R5579 VSS.n3889 VSS 128.655
R5580 VSS.n1203 VSS.t34 128.655
R5581 VSS.n896 VSS.t131 128.655
R5582 VSS.n578 VSS.t55 128.655
R5583 VSS.n4237 VSS.t447 120.733
R5584 VSS.n4245 VSS.t163 120.733
R5585 VSS.n3497 VSS.t135 120.733
R5586 VSS.n3505 VSS.t165 120.733
R5587 VSS.n3611 VSS.t514 120.733
R5588 VSS.n3619 VSS.t149 120.733
R5589 VSS.n3725 VSS.t401 120.733
R5590 VSS.n3733 VSS.t141 120.733
R5591 VSS.n3839 VSS.t507 120.733
R5592 VSS.n3847 VSS.t89 120.733
R5593 VSS.n4167 VSS.n4166 120.079
R5594 VSS.n4159 VSS.n4158 120.079
R5595 VSS.n4140 VSS.n4139 120.079
R5596 VSS.n4126 VSS.n4125 120.079
R5597 VSS.n4110 VSS.n4109 120.079
R5598 VSS.n4098 VSS.n4097 120.079
R5599 VSS.n4084 VSS.n4083 120.079
R5600 VSS.n4070 VSS.n4069 120.079
R5601 VSS.n34 VSS.n33 120.079
R5602 VSS.n4053 VSS.n4052 120.079
R5603 VSS.n4041 VSS.n4040 120.079
R5604 VSS.n4027 VSS.n4026 120.079
R5605 VSS.n4013 VSS.n4012 120.079
R5606 VSS.n3998 VSS.n3997 120.079
R5607 VSS.n3984 VSS.n3983 120.079
R5608 VSS.n3969 VSS.n3968 120.079
R5609 VSS.n3955 VSS.n3954 120.079
R5610 VSS.n48 VSS.n47 120.079
R5611 VSS.n1227 VSS.t237 120.079
R5612 VSS.n1071 VSS.t424 120.079
R5613 VSS.n161 VSS.t61 120.079
R5614 VSS.n753 VSS.t470 120.079
R5615 VSS.n206 VSS.t571 120.079
R5616 VSS.n435 VSS.t85 120.079
R5617 VSS.n251 VSS.t376 120.079
R5618 VSS.n86 VSS.n85 116.219
R5619 VSS.n3321 VSS.n3320 116.219
R5620 VSS.n3291 VSS.n3290 116.219
R5621 VSS.n3262 VSS.n3261 116.219
R5622 VSS.n3232 VSS.n3222 116.219
R5623 VSS.n3195 VSS.n3192 116.219
R5624 VSS.n3163 VSS.n3162 116.219
R5625 VSS.n3156 VSS.n3155 116.219
R5626 VSS.n3126 VSS.n3125 116.219
R5627 VSS.n3096 VSS.n3095 116.219
R5628 VSS.n3390 VSS.t536 114.775
R5629 VSS.n4002 VSS.n4001 114.749
R5630 VSS.n2023 VSS.n2022 113.207
R5631 VSS.n2138 VSS.n2137 113.207
R5632 VSS.n2441 VSS.n2440 113.207
R5633 VSS.n2793 VSS.n2792 113.207
R5634 VSS.n358 VSS.n357 113.207
R5635 VSS.n676 VSS.n675 113.207
R5636 VSS.n994 VSS.n993 113.207
R5637 VSS.n1286 VSS.n1285 113.207
R5638 VSS.n1956 VSS.n1955 113.207
R5639 VSS.n1855 VSS.n1854 113.207
R5640 VSS.n1754 VSS.n1753 113.207
R5641 VSS.n1653 VSS.n1652 113.207
R5642 VSS.n1552 VSS.n1551 113.207
R5643 VSS.n4250 VSS.n4249 113.207
R5644 VSS.n3510 VSS.n3509 113.207
R5645 VSS.n3624 VSS.n3623 113.207
R5646 VSS.n3738 VSS.n3737 113.207
R5647 VSS.n3852 VSS.n3851 113.207
R5648 VSS.t381 VSS.n4168 111.501
R5649 VSS.n22 VSS.t283 111.501
R5650 VSS.n3410 VSS.n3409 109.3
R5651 VSS.n3908 VSS.n3907 109.3
R5652 VSS.n3357 VSS.n3356 109.3
R5653 VSS.n2101 VSS.n2100 109.231
R5654 VSS.n150 VSS.n149 109.231
R5655 VSS.n127 VSS.n126 109.231
R5656 VSS.n1421 VSS.n1420 109.231
R5657 VSS.n1436 VSS.n1435 109.231
R5658 VSS.n1451 VSS.n1450 109.231
R5659 VSS.n1466 VSS.n1465 109.231
R5660 VSS.n1481 VSS.n1480 109.231
R5661 VSS.n5 VSS.n4 109.231
R5662 VSS.n3552 VSS.n3551 109.231
R5663 VSS.n3666 VSS.n3665 109.231
R5664 VSS.n3780 VSS.n3779 109.231
R5665 VSS.n4178 VSS.n4177 109.231
R5666 VSS.n2330 VSS.n2320 108.416
R5667 VSS.n2682 VSS.n2672 108.416
R5668 VSS.n3034 VSS.n3024 108.416
R5669 VSS.n230 VSS.n229 108.416
R5670 VSS.n185 VSS.n184 108.416
R5671 VSS.n3200 VSS.t333 108.328
R5672 VSS.n3403 VSS.n3402 108.254
R5673 VSS.n3921 VSS.n3920 108.254
R5674 VSS.n1999 VSS.n1998 107.478
R5675 VSS.n2087 VSS.n2086 107.478
R5676 VSS.n2114 VSS.n2113 107.478
R5677 VSS.n3427 VSS.n3426 107.478
R5678 VSS.n3897 VSS.n3896 107.478
R5679 VSS.n1189 VSS.n1188 107.478
R5680 VSS.n1233 VSS.n1232 107.478
R5681 VSS.n132 VSS.n131 107.478
R5682 VSS.n1416 VSS.n1415 107.478
R5683 VSS.n1879 VSS.n1878 107.478
R5684 VSS.n1431 VSS.n1430 107.478
R5685 VSS.n1778 VSS.n1777 107.478
R5686 VSS.n1446 VSS.n1445 107.478
R5687 VSS.n1677 VSS.n1676 107.478
R5688 VSS.n1461 VSS.n1460 107.478
R5689 VSS.n1576 VSS.n1575 107.478
R5690 VSS.n1476 VSS.n1475 107.478
R5691 VSS.n1980 VSS.n1979 107.478
R5692 VSS.n4192 VSS.n4191 107.478
R5693 VSS.n4277 VSS.n7 107.478
R5694 VSS.n3452 VSS.n3451 107.478
R5695 VSS.n3539 VSS.n3439 107.478
R5696 VSS.n3566 VSS.n3565 107.478
R5697 VSS.n3653 VSS.n3437 107.478
R5698 VSS.n3680 VSS.n3679 107.478
R5699 VSS.n3767 VSS.n3435 107.478
R5700 VSS.n3794 VSS.n3793 107.478
R5701 VSS.n3882 VSS.n3881 107.478
R5702 VSS.n81 VSS.t399 107.195
R5703 VSS.n2288 VSS.n2279 106.731
R5704 VSS.n2360 VSS.n112 106.731
R5705 VSS.n2640 VSS.n2631 106.731
R5706 VSS.n2712 VSS.n101 106.731
R5707 VSS.n2992 VSS.n2983 106.731
R5708 VSS.n4154 VSS.n13 106.731
R5709 VSS.n27 VSS.n15 106.731
R5710 VSS.n259 VSS.n250 106.731
R5711 VSS.n240 VSS.n231 106.731
R5712 VSS.n214 VSS.n205 106.731
R5713 VSS.n195 VSS.n186 106.731
R5714 VSS.n169 VSS.n160 106.731
R5715 VSS.n2062 VSS.n2061 106.038
R5716 VSS.n2208 VSS.n2207 106.038
R5717 VSS.n2560 VSS.n2559 106.038
R5718 VSS.n2912 VSS.n2911 106.038
R5719 VSS.n495 VSS.n494 106.038
R5720 VSS.n813 VSS.n812 106.038
R5721 VSS.n1131 VSS.n1130 106.038
R5722 VSS.n1372 VSS.n1371 106.038
R5723 VSS.n1917 VSS.n1916 106.038
R5724 VSS.n1816 VSS.n1815 106.038
R5725 VSS.n1715 VSS.n1714 106.038
R5726 VSS.n1614 VSS.n1613 106.038
R5727 VSS.n1513 VSS.n1512 106.038
R5728 VSS.n4211 VSS.n4210 106.038
R5729 VSS.n3471 VSS.n3470 106.038
R5730 VSS.n3585 VSS.n3584 106.038
R5731 VSS.n3699 VSS.n3698 106.038
R5732 VSS.n3813 VSS.n3812 106.038
R5733 VSS.n60 VSS.t560 105.835
R5734 VSS.n54 VSS.t179 105.835
R5735 VSS.n2063 VSS.t153 105.6
R5736 VSS.n3367 VSS.n3366 104.719
R5737 VSS.n3944 VSS.t389 104.103
R5738 VSS.n3345 VSS.n3344 103.942
R5739 VSS.n1373 VSS.t93 102.924
R5740 VSS.n1141 VSS.t294 102.924
R5741 VSS.n823 VSS.t620 102.924
R5742 VSS.n505 VSS.t689 102.924
R5743 VSS.n76 VSS.t659 100.21
R5744 VSS.n1361 VSS.n1358 98.5005
R5745 VSS.n1351 VSS.n1348 98.5005
R5746 VSS.n1341 VSS.n1338 98.5005
R5747 VSS.n1331 VSS.n1328 98.5005
R5748 VSS.n1321 VSS.n1318 98.5005
R5749 VSS.n1311 VSS.n1308 98.5005
R5750 VSS.n1301 VSS.n1298 98.5005
R5751 VSS.n1291 VSS.n1288 98.5005
R5752 VSS.n1279 VSS.n1276 98.5005
R5753 VSS.n1269 VSS.n1266 98.5005
R5754 VSS.n1259 VSS.n1256 98.5005
R5755 VSS.n1250 VSS.n1247 98.5005
R5756 VSS.n1239 VSS.n1236 98.5005
R5757 VSS.n1229 VSS.n1226 98.5005
R5758 VSS.n138 VSS.n137 98.5005
R5759 VSS.n1217 VSS.n135 98.5005
R5760 VSS.n1205 VSS.n1202 98.5005
R5761 VSS.n1195 VSS.n1192 98.5005
R5762 VSS.n1185 VSS.n1182 98.5005
R5763 VSS.n1174 VSS.n1171 98.5005
R5764 VSS.n1164 VSS.n1161 98.5005
R5765 VSS.n1154 VSS.n1151 98.5005
R5766 VSS VSS.n2354 96.8005
R5767 VSS VSS.n2706 96.8005
R5768 VSS.n1922 VSS.t468 94.8508
R5769 VSS.n1821 VSS.t676 94.8508
R5770 VSS.n1720 VSS.t212 94.8508
R5771 VSS.n1619 VSS.t43 94.8508
R5772 VSS.n1518 VSS.t551 94.8508
R5773 VSS.t236 VSS.n1359 94.3475
R5774 VSS.n1183 VSS.t30 94.3475
R5775 VSS.n1085 VSS.t646 94.3475
R5776 VSS.n187 VSS.t133 94.3475
R5777 VSS.n767 VSS.t254 94.3475
R5778 VSS.n232 VSS.t57 94.3475
R5779 VSS.n449 VSS.t322 94.3475
R5780 VSS.n3393 VSS.n62 88.1769
R5781 VSS.n2171 VSS.n2170 88.0005
R5782 VSS.n2185 VSS.n2184 88.0005
R5783 VSS.n2199 VSS.n2198 88.0005
R5784 VSS.n2215 VSS.n2214 88.0005
R5785 VSS.n2229 VSS.n2228 88.0005
R5786 VSS.n2243 VSS.n2242 88.0005
R5787 VSS.n2257 VSS.n2256 88.0005
R5788 VSS.n2271 VSS.n2270 88.0005
R5789 VSS.n2285 VSS.n2284 88.0005
R5790 VSS.n2298 VSS.n2297 88.0005
R5791 VSS.n2312 VSS.n2311 88.0005
R5792 VSS.n2324 VSS.n2323 88.0005
R5793 VSS.n2340 VSS.n2339 88.0005
R5794 VSS.n2354 VSS.n117 88.0005
R5795 VSS.n2357 VSS.n2356 88.0005
R5796 VSS.n2370 VSS.n2369 88.0005
R5797 VSS.n2383 VSS.n2382 88.0005
R5798 VSS.n2396 VSS.n2395 88.0005
R5799 VSS.n2410 VSS.n2409 88.0005
R5800 VSS.n2424 VSS.n2423 88.0005
R5801 VSS.n2437 VSS.n2436 88.0005
R5802 VSS.n2453 VSS.n2452 88.0005
R5803 VSS.n2467 VSS.n2466 88.0005
R5804 VSS.n2481 VSS.n2480 88.0005
R5805 VSS.n2495 VSS.n2494 88.0005
R5806 VSS.n2509 VSS.n2508 88.0005
R5807 VSS.n2523 VSS.n2522 88.0005
R5808 VSS.n2537 VSS.n2536 88.0005
R5809 VSS.n2551 VSS.n2550 88.0005
R5810 VSS.n2567 VSS.n2566 88.0005
R5811 VSS.n2581 VSS.n2580 88.0005
R5812 VSS.n2595 VSS.n2594 88.0005
R5813 VSS.n2609 VSS.n2608 88.0005
R5814 VSS.n2623 VSS.n2622 88.0005
R5815 VSS.n2637 VSS.n2636 88.0005
R5816 VSS.n2650 VSS.n2649 88.0005
R5817 VSS.n2664 VSS.n2663 88.0005
R5818 VSS.n2676 VSS.n2675 88.0005
R5819 VSS.n2692 VSS.n2691 88.0005
R5820 VSS.n2706 VSS.n106 88.0005
R5821 VSS.n2709 VSS.n2708 88.0005
R5822 VSS.n2722 VSS.n2721 88.0005
R5823 VSS.n2735 VSS.n2734 88.0005
R5824 VSS.n2748 VSS.n2747 88.0005
R5825 VSS.n2762 VSS.n2761 88.0005
R5826 VSS.n2776 VSS.n2775 88.0005
R5827 VSS.n2789 VSS.n2788 88.0005
R5828 VSS.n2805 VSS.n2804 88.0005
R5829 VSS.n2819 VSS.n2818 88.0005
R5830 VSS.n2833 VSS.n2832 88.0005
R5831 VSS.n2847 VSS.n2846 88.0005
R5832 VSS.n2861 VSS.n2860 88.0005
R5833 VSS.n2875 VSS.n2874 88.0005
R5834 VSS.n2889 VSS.n2888 88.0005
R5835 VSS.n2903 VSS.n2902 88.0005
R5836 VSS.n2919 VSS.n2918 88.0005
R5837 VSS.n2933 VSS.n2932 88.0005
R5838 VSS.n2947 VSS.n2946 88.0005
R5839 VSS.n2961 VSS.n2960 88.0005
R5840 VSS.n2975 VSS.n2974 88.0005
R5841 VSS.n2989 VSS.n2988 88.0005
R5842 VSS.n3002 VSS.n3001 88.0005
R5843 VSS.n3016 VSS.n3015 88.0005
R5844 VSS.n3028 VSS.n3027 88.0005
R5845 VSS.n97 VSS.n96 88.0005
R5846 VSS.n3048 VSS.n3047 88.0005
R5847 VSS.n3063 VSS.n3062 88.0005
R5848 VSS.n3077 VSS.n3076 88.0005
R5849 VSS.n1143 VSS.n1142 85.7705
R5850 VSS.n1085 VSS.n1084 85.7705
R5851 VSS.n1071 VSS.n1070 85.7705
R5852 VSS.n1057 VSS.n1056 85.7705
R5853 VSS.n1043 VSS.n1042 85.7705
R5854 VSS.n1029 VSS.n1028 85.7705
R5855 VSS.n1029 VSS.t13 85.7705
R5856 VSS.n1015 VSS.n1014 85.7705
R5857 VSS.n1001 VSS.n1000 85.7705
R5858 VSS.n985 VSS.n984 85.7705
R5859 VSS.n971 VSS.n970 85.7705
R5860 VSS.n957 VSS.n956 85.7705
R5861 VSS.n153 VSS.n152 85.7705
R5862 VSS.n940 VSS.n939 85.7705
R5863 VSS.n163 VSS.n162 85.7705
R5864 VSS.n918 VSS.n913 85.7705
R5865 VSS.n921 VSS.n920 85.7705
R5866 VSS.n181 VSS.n180 85.7705
R5867 VSS.n898 VSS.n897 85.7705
R5868 VSS.n884 VSS.n883 85.7705
R5869 VSS.n189 VSS.n188 85.7705
R5870 VSS.n867 VSS.n866 85.7705
R5871 VSS.n853 VSS.n852 85.7705
R5872 VSS.n839 VSS.n838 85.7705
R5873 VSS.n825 VSS.n824 85.7705
R5874 VSS.n767 VSS.n766 85.7705
R5875 VSS.n753 VSS.n752 85.7705
R5876 VSS.n739 VSS.n738 85.7705
R5877 VSS.n725 VSS.n724 85.7705
R5878 VSS.n711 VSS.n710 85.7705
R5879 VSS.n711 VSS.t627 85.7705
R5880 VSS.n697 VSS.n696 85.7705
R5881 VSS.n683 VSS.n682 85.7705
R5882 VSS.n667 VSS.n666 85.7705
R5883 VSS.n653 VSS.n652 85.7705
R5884 VSS.n639 VSS.n638 85.7705
R5885 VSS.n198 VSS.n197 85.7705
R5886 VSS.n622 VSS.n621 85.7705
R5887 VSS.n208 VSS.n207 85.7705
R5888 VSS.n600 VSS.n595 85.7705
R5889 VSS.n603 VSS.n602 85.7705
R5890 VSS.n226 VSS.n225 85.7705
R5891 VSS.n580 VSS.n579 85.7705
R5892 VSS.n566 VSS.n565 85.7705
R5893 VSS.n234 VSS.n233 85.7705
R5894 VSS.n549 VSS.n548 85.7705
R5895 VSS.n535 VSS.n534 85.7705
R5896 VSS.n521 VSS.n520 85.7705
R5897 VSS.n507 VSS.n506 85.7705
R5898 VSS.n449 VSS.n448 85.7705
R5899 VSS.n435 VSS.n434 85.7705
R5900 VSS.n421 VSS.n420 85.7705
R5901 VSS.n407 VSS.n406 85.7705
R5902 VSS.n393 VSS.n392 85.7705
R5903 VSS.n393 VSS.t587 85.7705
R5904 VSS.n379 VSS.n378 85.7705
R5905 VSS.n365 VSS.n364 85.7705
R5906 VSS.n349 VSS.n348 85.7705
R5907 VSS.n335 VSS.n334 85.7705
R5908 VSS.n321 VSS.n320 85.7705
R5909 VSS.n243 VSS.n242 85.7705
R5910 VSS.n304 VSS.n303 85.7705
R5911 VSS.n253 VSS.n252 85.7705
R5912 VSS.n284 VSS.n283 85.7705
R5913 VSS.n145 VSS.n141 83.8127
R5914 VSS.n3184 VSS.t341 82.839
R5915 VSS.n4165 VSS.n10 81.1181
R5916 VSS.n4160 VSS.n4156 81.1181
R5917 VSS.n4141 VSS.n4137 81.1181
R5918 VSS.n4127 VSS.n4124 81.1181
R5919 VSS.n23 VSS.n19 81.1181
R5920 VSS.n4111 VSS.n4107 81.1181
R5921 VSS.n4099 VSS.n4095 81.1181
R5922 VSS.n4085 VSS.n4081 81.1181
R5923 VSS.n4071 VSS.n4067 81.1181
R5924 VSS.n35 VSS.n31 81.1181
R5925 VSS.n4054 VSS.n4050 81.1181
R5926 VSS.n4042 VSS.n4038 81.1181
R5927 VSS.n4028 VSS.n4024 81.1181
R5928 VSS.n4014 VSS.n4010 81.1181
R5929 VSS.n3999 VSS.n3995 81.1181
R5930 VSS.n3985 VSS.n3981 81.1181
R5931 VSS.n3970 VSS.n3966 81.1181
R5932 VSS.n3956 VSS.n3952 81.1181
R5933 VSS.n49 VSS.n45 81.1181
R5934 VSS.n3352 VSS 80.7344
R5935 VSS.n3212 VSS.t335 79.6529
R5936 VSS.n2028 VSS.t145 79.2005
R5937 VSS.n2036 VSS.t260 79.2005
R5938 VSS.n2143 VSS.t169 79.2005
R5939 VSS.n2151 VSS.t421 79.2005
R5940 VSS.n2467 VSS.t105 79.2005
R5941 VSS.n2819 VSS.t262 79.2005
R5942 VSS.n1926 VSS.t279 79.0424
R5943 VSS.n1825 VSS.t498 79.0424
R5944 VSS.n1724 VSS.t297 79.0424
R5945 VSS.n1623 VSS.t200 79.0424
R5946 VSS.n1522 VSS.t505 79.0424
R5947 VSS.n4084 VSS.t474 77.1935
R5948 VSS.n1323 VSS.t558 77.1935
R5949 VSS.n1303 VSS.t91 77.1935
R5950 VSS.n1113 VSS.t32 77.1935
R5951 VSS.n795 VSS.t129 77.1935
R5952 VSS.n477 VSS.t53 77.1935
R5953 VSS.n2022 VSS.t362 75.7148
R5954 VSS.n2137 VSS.t259 75.7148
R5955 VSS.n2440 VSS.t649 75.7148
R5956 VSS.n2792 VSS.t486 75.7148
R5957 VSS.n357 VSS.t84 75.7148
R5958 VSS.n675 VSS.t473 75.7148
R5959 VSS.n993 VSS.t427 75.7148
R5960 VSS.n1285 VSS.t317 75.7148
R5961 VSS.n1955 VSS.t449 75.7148
R5962 VSS.n1854 VSS.t39 75.7148
R5963 VSS.n1753 VSS.t102 75.7148
R5964 VSS.n1652 VSS.t122 75.7148
R5965 VSS.n1551 VSS.t225 75.7148
R5966 VSS.n4249 VSS.t510 75.7148
R5967 VSS.n3509 VSS.t453 75.7148
R5968 VSS.n3623 VSS.t300 75.7148
R5969 VSS.n3737 VSS.t548 75.7148
R5970 VSS.n3851 VSS.t368 75.7148
R5971 VSS VSS.n55 75.6886
R5972 VSS.n3339 VSS 70.6427
R5973 VSS.n2171 VSS.t190 70.4005
R5974 VSS.n2523 VSS.t456 70.4005
R5975 VSS.n2875 VSS.t419 70.4005
R5976 VSS.n3331 VSS.t355 70.0946
R5977 VSS VSS.n139 68.6165
R5978 VSS.n1172 VSS.t267 68.6165
R5979 VSS VSS.n918 68.6165
R5980 VSS.n865 VSS.t16 68.6165
R5981 VSS VSS.n600 68.6165
R5982 VSS.n547 VSS.t527 68.6165
R5983 VSS VSS.n284 68.6165
R5984 VSS.n4228 VSS.t511 67.0737
R5985 VSS.n3488 VSS.t454 67.0737
R5986 VSS.n3602 VSS.t301 67.0737
R5987 VSS.n3716 VSS.t549 67.0737
R5988 VSS.n3830 VSS.t365 67.0737
R5989 VSS.n3973 VSS.n3972 65.3332
R5990 VSS.n1918 VSS.t682 63.234
R5991 VSS.n1817 VSS.t582 63.234
R5992 VSS.n1716 VSS.t590 63.234
R5993 VSS.n1615 VSS.t359 63.234
R5994 VSS.n1514 VSS.t115 63.234
R5995 VSS.n4001 VSS.t577 62.3526
R5996 VSS.n62 VSS.n61 61.7239
R5997 VSS.n2170 VSS.n2169 61.6005
R5998 VSS.n2184 VSS.n2183 61.6005
R5999 VSS.n2198 VSS.n2197 61.6005
R6000 VSS.n2214 VSS.n2213 61.6005
R6001 VSS.n2228 VSS.n2227 61.6005
R6002 VSS.n2242 VSS.n2241 61.6005
R6003 VSS.n2256 VSS.n2255 61.6005
R6004 VSS.n2270 VSS.n2269 61.6005
R6005 VSS.n2284 VSS.n2283 61.6005
R6006 VSS.n2297 VSS.n2296 61.6005
R6007 VSS.n2311 VSS.n2310 61.6005
R6008 VSS.n2323 VSS.n2322 61.6005
R6009 VSS.n2339 VSS.n2338 61.6005
R6010 VSS.n117 VSS.n116 61.6005
R6011 VSS.n2356 VSS.n2355 61.6005
R6012 VSS.n2369 VSS.n2368 61.6005
R6013 VSS.n2382 VSS.n2381 61.6005
R6014 VSS.n2395 VSS.n2394 61.6005
R6015 VSS.n2409 VSS.n2408 61.6005
R6016 VSS.n2423 VSS.n2422 61.6005
R6017 VSS.n2436 VSS.t648 61.6005
R6018 VSS.n2452 VSS.n2451 61.6005
R6019 VSS.n2466 VSS.n2465 61.6005
R6020 VSS.n2480 VSS.n2479 61.6005
R6021 VSS.n2494 VSS.n2493 61.6005
R6022 VSS.n2508 VSS.n2507 61.6005
R6023 VSS.n2522 VSS.n2521 61.6005
R6024 VSS.n2536 VSS.n2535 61.6005
R6025 VSS.n2550 VSS.n2549 61.6005
R6026 VSS.n2566 VSS.n2565 61.6005
R6027 VSS.n2580 VSS.n2579 61.6005
R6028 VSS.n2594 VSS.n2593 61.6005
R6029 VSS.n2608 VSS.n2607 61.6005
R6030 VSS.n2622 VSS.n2621 61.6005
R6031 VSS.n2636 VSS.n2635 61.6005
R6032 VSS.n2649 VSS.n2648 61.6005
R6033 VSS.n2663 VSS.n2662 61.6005
R6034 VSS.n2675 VSS.n2674 61.6005
R6035 VSS.n2691 VSS.n2690 61.6005
R6036 VSS.n106 VSS.n105 61.6005
R6037 VSS.n2708 VSS.n2707 61.6005
R6038 VSS.n2721 VSS.n2720 61.6005
R6039 VSS.n2734 VSS.n2733 61.6005
R6040 VSS.n2747 VSS.n2746 61.6005
R6041 VSS.n2761 VSS.n2760 61.6005
R6042 VSS.n2775 VSS.n2774 61.6005
R6043 VSS.n2788 VSS.t485 61.6005
R6044 VSS.n2804 VSS.n2803 61.6005
R6045 VSS.n2818 VSS.n2817 61.6005
R6046 VSS.n2832 VSS.n2831 61.6005
R6047 VSS.n2846 VSS.n2845 61.6005
R6048 VSS.n2860 VSS.n2859 61.6005
R6049 VSS.n2874 VSS.n2873 61.6005
R6050 VSS.n2888 VSS.n2887 61.6005
R6051 VSS.n2902 VSS.n2901 61.6005
R6052 VSS.n2918 VSS.n2917 61.6005
R6053 VSS.n2932 VSS.n2931 61.6005
R6054 VSS.n2946 VSS.n2945 61.6005
R6055 VSS.n2960 VSS.n2959 61.6005
R6056 VSS.n2974 VSS.n2973 61.6005
R6057 VSS.n2988 VSS.n2987 61.6005
R6058 VSS.n3001 VSS.n3000 61.6005
R6059 VSS.n3015 VSS.n3014 61.6005
R6060 VSS.n3027 VSS.n3026 61.6005
R6061 VSS.n96 VSS.n95 61.6005
R6062 VSS.n3047 VSS.n3046 61.6005
R6063 VSS.n3062 VSS.n3061 61.6005
R6064 VSS.n3076 VSS.n3075 61.6005
R6065 VSS.n1142 VSS.n1141 60.0395
R6066 VSS.n1126 VSS.n1125 60.0395
R6067 VSS.t487 VSS.n1126 60.0395
R6068 VSS.n1112 VSS.n1111 60.0395
R6069 VSS.n1098 VSS.n1097 60.0395
R6070 VSS.n1084 VSS.n1083 60.0395
R6071 VSS.n1070 VSS.n1069 60.0395
R6072 VSS.n1056 VSS.n1055 60.0395
R6073 VSS.n1042 VSS.n1041 60.0395
R6074 VSS.n1028 VSS.n1027 60.0395
R6075 VSS.n1014 VSS.n1013 60.0395
R6076 VSS.n1000 VSS.n999 60.0395
R6077 VSS.n984 VSS.n983 60.0395
R6078 VSS.n970 VSS.n969 60.0395
R6079 VSS.n956 VSS.n955 60.0395
R6080 VSS.n152 VSS.n151 60.0395
R6081 VSS.n939 VSS.n938 60.0395
R6082 VSS.n162 VSS.n161 60.0395
R6083 VSS.n913 VSS.n912 60.0395
R6084 VSS.n920 VSS.n919 60.0395
R6085 VSS.n180 VSS.n179 60.0395
R6086 VSS.n897 VSS.n896 60.0395
R6087 VSS.n883 VSS.n882 60.0395
R6088 VSS.n188 VSS.n187 60.0395
R6089 VSS.n866 VSS.n865 60.0395
R6090 VSS.n852 VSS.n851 60.0395
R6091 VSS.n838 VSS.n837 60.0395
R6092 VSS.n824 VSS.n823 60.0395
R6093 VSS.n808 VSS.n807 60.0395
R6094 VSS.t231 VSS.n808 60.0395
R6095 VSS.n794 VSS.n793 60.0395
R6096 VSS.n780 VSS.n779 60.0395
R6097 VSS.n766 VSS.n765 60.0395
R6098 VSS.n752 VSS.n751 60.0395
R6099 VSS.n738 VSS.n737 60.0395
R6100 VSS.n724 VSS.n723 60.0395
R6101 VSS.n710 VSS.n709 60.0395
R6102 VSS.n696 VSS.n695 60.0395
R6103 VSS.n682 VSS.n681 60.0395
R6104 VSS.n666 VSS.n665 60.0395
R6105 VSS.n652 VSS.n651 60.0395
R6106 VSS.n638 VSS.n637 60.0395
R6107 VSS.n197 VSS.n196 60.0395
R6108 VSS.n621 VSS.n620 60.0395
R6109 VSS.n207 VSS.n206 60.0395
R6110 VSS.n595 VSS.n594 60.0395
R6111 VSS.n602 VSS.n601 60.0395
R6112 VSS.n225 VSS.n224 60.0395
R6113 VSS.n579 VSS.n578 60.0395
R6114 VSS.n565 VSS.n564 60.0395
R6115 VSS.n233 VSS.n232 60.0395
R6116 VSS.n548 VSS.n547 60.0395
R6117 VSS.n534 VSS.n533 60.0395
R6118 VSS.n520 VSS.n519 60.0395
R6119 VSS.n506 VSS.n505 60.0395
R6120 VSS.n490 VSS.n489 60.0395
R6121 VSS.t628 VSS.n490 60.0395
R6122 VSS.n476 VSS.n475 60.0395
R6123 VSS.n462 VSS.n461 60.0395
R6124 VSS.n448 VSS.n447 60.0395
R6125 VSS.n434 VSS.n433 60.0395
R6126 VSS.n420 VSS.n419 60.0395
R6127 VSS.n406 VSS.n405 60.0395
R6128 VSS.n392 VSS.n391 60.0395
R6129 VSS.n378 VSS.n377 60.0395
R6130 VSS.n364 VSS.n363 60.0395
R6131 VSS.n348 VSS.n347 60.0395
R6132 VSS.n334 VSS.n333 60.0395
R6133 VSS.n320 VSS.n319 60.0395
R6134 VSS.n242 VSS.n241 60.0395
R6135 VSS.n303 VSS.n302 60.0395
R6136 VSS.n252 VSS.n251 60.0395
R6137 VSS.n283 VSS.n282 60.0395
R6138 VSS.n1144 VSS.n1140 57.9417
R6139 VSS.n1128 VSS.n1124 57.9417
R6140 VSS.n1114 VSS.n1110 57.9417
R6141 VSS.n1100 VSS.n1096 57.9417
R6142 VSS.n1086 VSS.n1082 57.9417
R6143 VSS.n1072 VSS.n1068 57.9417
R6144 VSS.n1058 VSS.n1054 57.9417
R6145 VSS.n1044 VSS.n1040 57.9417
R6146 VSS.n1030 VSS.n1026 57.9417
R6147 VSS.n1016 VSS.n1012 57.9417
R6148 VSS.n1002 VSS.n998 57.9417
R6149 VSS.n986 VSS.n982 57.9417
R6150 VSS.n972 VSS.n968 57.9417
R6151 VSS.n958 VSS.n954 57.9417
R6152 VSS.n941 VSS.n937 57.9417
R6153 VSS.n917 VSS.n915 57.9417
R6154 VSS.n922 VSS.n911 57.9417
R6155 VSS.n182 VSS.n178 57.9417
R6156 VSS.n899 VSS.n895 57.9417
R6157 VSS.n885 VSS.n881 57.9417
R6158 VSS.n868 VSS.n864 57.9417
R6159 VSS.n854 VSS.n850 57.9417
R6160 VSS.n840 VSS.n836 57.9417
R6161 VSS.n826 VSS.n822 57.9417
R6162 VSS.n810 VSS.n806 57.9417
R6163 VSS.n796 VSS.n792 57.9417
R6164 VSS.n782 VSS.n778 57.9417
R6165 VSS.n768 VSS.n764 57.9417
R6166 VSS.n754 VSS.n750 57.9417
R6167 VSS.n740 VSS.n736 57.9417
R6168 VSS.n726 VSS.n722 57.9417
R6169 VSS.n712 VSS.n708 57.9417
R6170 VSS.n698 VSS.n694 57.9417
R6171 VSS.n684 VSS.n680 57.9417
R6172 VSS.n668 VSS.n664 57.9417
R6173 VSS.n654 VSS.n650 57.9417
R6174 VSS.n640 VSS.n636 57.9417
R6175 VSS.n623 VSS.n619 57.9417
R6176 VSS.n599 VSS.n597 57.9417
R6177 VSS.n604 VSS.n593 57.9417
R6178 VSS.n227 VSS.n223 57.9417
R6179 VSS.n581 VSS.n577 57.9417
R6180 VSS.n567 VSS.n563 57.9417
R6181 VSS.n550 VSS.n546 57.9417
R6182 VSS.n536 VSS.n532 57.9417
R6183 VSS.n522 VSS.n518 57.9417
R6184 VSS.n508 VSS.n504 57.9417
R6185 VSS.n492 VSS.n488 57.9417
R6186 VSS.n478 VSS.n474 57.9417
R6187 VSS.n464 VSS.n460 57.9417
R6188 VSS.n450 VSS.n446 57.9417
R6189 VSS.n436 VSS.n432 57.9417
R6190 VSS.n422 VSS.n418 57.9417
R6191 VSS.n408 VSS.n404 57.9417
R6192 VSS.n394 VSS.n390 57.9417
R6193 VSS.n380 VSS.n376 57.9417
R6194 VSS.n366 VSS.n362 57.9417
R6195 VSS.n350 VSS.n346 57.9417
R6196 VSS.n336 VSS.n332 57.9417
R6197 VSS.n322 VSS.n318 57.9417
R6198 VSS.n305 VSS.n301 57.9417
R6199 VSS.n281 VSS.n280 57.9417
R6200 VSS.n2172 VSS.n2168 57.9417
R6201 VSS.n2186 VSS.n2182 57.9417
R6202 VSS.n2200 VSS.n2196 57.9417
R6203 VSS.n2216 VSS.n2212 57.9417
R6204 VSS.n2230 VSS.n2226 57.9417
R6205 VSS.n2244 VSS.n2240 57.9417
R6206 VSS.n2258 VSS.n2254 57.9417
R6207 VSS.n2272 VSS.n2268 57.9417
R6208 VSS.n2286 VSS.n2282 57.9417
R6209 VSS.n2299 VSS.n2295 57.9417
R6210 VSS.n2313 VSS.n2309 57.9417
R6211 VSS.n2341 VSS.n2337 57.9417
R6212 VSS.n2353 VSS.n119 57.9417
R6213 VSS.n2358 VSS.n115 57.9417
R6214 VSS.n2371 VSS.n2367 57.9417
R6215 VSS.n2384 VSS.n2380 57.9417
R6216 VSS.n2397 VSS.n2393 57.9417
R6217 VSS.n2411 VSS.n2407 57.9417
R6218 VSS.n2425 VSS.n2421 57.9417
R6219 VSS.n2438 VSS.n2435 57.9417
R6220 VSS.n2454 VSS.n2450 57.9417
R6221 VSS.n2468 VSS.n2464 57.9417
R6222 VSS.n2482 VSS.n2478 57.9417
R6223 VSS.n2496 VSS.n2492 57.9417
R6224 VSS.n2510 VSS.n2506 57.9417
R6225 VSS.n2524 VSS.n2520 57.9417
R6226 VSS.n2538 VSS.n2534 57.9417
R6227 VSS.n2552 VSS.n2548 57.9417
R6228 VSS.n2568 VSS.n2564 57.9417
R6229 VSS.n2582 VSS.n2578 57.9417
R6230 VSS.n2596 VSS.n2592 57.9417
R6231 VSS.n2610 VSS.n2606 57.9417
R6232 VSS.n2624 VSS.n2620 57.9417
R6233 VSS.n2638 VSS.n2634 57.9417
R6234 VSS.n2651 VSS.n2647 57.9417
R6235 VSS.n2665 VSS.n2661 57.9417
R6236 VSS.n2693 VSS.n2689 57.9417
R6237 VSS.n2705 VSS.n108 57.9417
R6238 VSS.n2710 VSS.n104 57.9417
R6239 VSS.n2723 VSS.n2719 57.9417
R6240 VSS.n2736 VSS.n2732 57.9417
R6241 VSS.n2749 VSS.n2745 57.9417
R6242 VSS.n2763 VSS.n2759 57.9417
R6243 VSS.n2777 VSS.n2773 57.9417
R6244 VSS.n2790 VSS.n2787 57.9417
R6245 VSS.n2806 VSS.n2802 57.9417
R6246 VSS.n2820 VSS.n2816 57.9417
R6247 VSS.n2834 VSS.n2830 57.9417
R6248 VSS.n2848 VSS.n2844 57.9417
R6249 VSS.n2862 VSS.n2858 57.9417
R6250 VSS.n2876 VSS.n2872 57.9417
R6251 VSS.n2890 VSS.n2886 57.9417
R6252 VSS.n2904 VSS.n2900 57.9417
R6253 VSS.n2920 VSS.n2916 57.9417
R6254 VSS.n2934 VSS.n2930 57.9417
R6255 VSS.n2948 VSS.n2944 57.9417
R6256 VSS.n2962 VSS.n2958 57.9417
R6257 VSS.n2976 VSS.n2972 57.9417
R6258 VSS.n2990 VSS.n2986 57.9417
R6259 VSS.n3003 VSS.n2999 57.9417
R6260 VSS.n3017 VSS.n3013 57.9417
R6261 VSS.n98 VSS.n94 57.9417
R6262 VSS.n3049 VSS.n3045 57.9417
R6263 VSS.n3064 VSS.n3060 57.9417
R6264 VSS.n3078 VSS.n3074 57.9417
R6265 VSS.n3330 VSS.n84 57.9417
R6266 VSS.n3318 VSS.n3314 57.9417
R6267 VSS.n3304 VSS.n3300 57.9417
R6268 VSS.n3288 VSS.n3284 57.9417
R6269 VSS.n3274 VSS.n3271 57.9417
R6270 VSS.n3259 VSS.n3255 57.9417
R6271 VSS.n3245 VSS.n3241 57.9417
R6272 VSS.n3230 VSS.n3226 57.9417
R6273 VSS.n3215 VSS.n3211 57.9417
R6274 VSS.n3201 VSS.n3197 57.9417
R6275 VSS.n3185 VSS.n3181 57.9417
R6276 VSS.n3171 VSS.n3167 57.9417
R6277 VSS.n3153 VSS.n3149 57.9417
R6278 VSS.n3139 VSS.n3135 57.9417
R6279 VSS.n3123 VSS.n3119 57.9417
R6280 VSS.n3109 VSS.n3105 57.9417
R6281 VSS.n3093 VSS.n3089 57.9417
R6282 VSS.n3380 VSS.n71 57.9417
R6283 VSS.n3392 VSS.n64 57.9417
R6284 VSS.n3170 VSS.t329 57.3502
R6285 VSS.n15 VSS.t7 57.1434
R6286 VSS.n3024 VSS.t518 54.2862
R6287 VSS.n2086 VSS.t429 54.2862
R6288 VSS.n2100 VSS.t439 54.2862
R6289 VSS.n2279 VSS.t633 54.2862
R6290 VSS.n2320 VSS.t23 54.2862
R6291 VSS.n2631 VSS.t372 54.2862
R6292 VSS.n2672 VSS.t409 54.2862
R6293 VSS.n2983 VSS.t374 54.2862
R6294 VSS.n15 VSS.t284 54.2862
R6295 VSS.n231 VSS.t528 54.2862
R6296 VSS.n229 VSS.t56 54.2862
R6297 VSS.n186 VSS.t17 54.2862
R6298 VSS.n184 VSS.t132 54.2862
R6299 VSS.n1188 VSS.t268 54.2862
R6300 VSS.n149 VSS.t35 54.2862
R6301 VSS.n131 VSS.t270 54.2862
R6302 VSS.n126 VSS.t252 54.2862
R6303 VSS.n1415 VSS.t29 54.2862
R6304 VSS.n1420 VSS.t467 54.2862
R6305 VSS.n1430 VSS.t403 54.2862
R6306 VSS.n1435 VSS.t675 54.2862
R6307 VSS.n1445 VSS.t405 54.2862
R6308 VSS.n1450 VSS.t211 54.2862
R6309 VSS.n1460 VSS.t51 54.2862
R6310 VSS.n1465 VSS.t42 54.2862
R6311 VSS.n1475 VSS.t27 54.2862
R6312 VSS.n1480 VSS.t556 54.2862
R6313 VSS.n4191 VSS.t15 54.2862
R6314 VSS.n4 VSS.t309 54.2862
R6315 VSS.n3451 VSS.t118 54.2862
R6316 VSS.n3551 VSS.t291 54.2862
R6317 VSS.n3565 VSS.t19 54.2862
R6318 VSS.n3665 VSS.t110 54.2862
R6319 VSS.n3679 VSS.t272 54.2862
R6320 VSS.n3779 VSS.t209 54.2862
R6321 VSS.n3793 VSS.t160 54.2862
R6322 VSS.n4177 VSS.t246 54.2862
R6323 VSS.n3227 VSS.t347 54.1641
R6324 VSS.n4053 VSS.t229 51.4625
R6325 VSS.n1360 VSS.t236 51.4625
R6326 VSS.n1099 VSS.t60 51.4625
R6327 VSS.n781 VSS.t574 51.4625
R6328 VSS.n463 VSS.t375 51.4625
R6329 VSS.n1951 VSS.t680 47.4256
R6330 VSS.n1943 VSS.t188 47.4256
R6331 VSS.n1850 VSS.t580 47.4256
R6332 VSS.n1842 VSS.t521 47.4256
R6333 VSS.n1749 VSS.t592 47.4256
R6334 VSS.n1741 VSS.t186 47.4256
R6335 VSS.n1648 VSS.t357 47.4256
R6336 VSS.n1640 VSS.t99 47.4256
R6337 VSS.n1547 VSS.t113 47.4256
R6338 VSS.n1539 VSS.t461 47.4256
R6339 VSS.n2328 VSS.n2327 47.1979
R6340 VSS.n2680 VSS.n2679 47.1979
R6341 VSS.n3032 VSS.n3031 47.1979
R6342 VSS.n257 VSS.n256 47.1889
R6343 VSS.n238 VSS.n237 47.1889
R6344 VSS.n212 VSS.n211 47.1889
R6345 VSS.n193 VSS.n192 47.1889
R6346 VSS.n167 VSS.n166 47.1889
R6347 VSS.n247 VSS.n246 47.1845
R6348 VSS.n202 VSS.n201 47.1845
R6349 VSS.n157 VSS.n156 47.1845
R6350 VSS.n3317 VSS.t345 44.6059
R6351 VSS.n2045 VSS.t363 44.0005
R6352 VSS.n2160 VSS.t256 44.0005
R6353 VSS.n2509 VSS.t650 44.0005
R6354 VSS.n2861 VSS.t483 44.0005
R6355 VSS.n1343 VSS.t314 42.8855
R6356 VSS.n2061 VSS.t441 41.4291
R6357 VSS.n2207 VSS.t25 41.4291
R6358 VSS.n2559 VSS.t411 41.4291
R6359 VSS.n2911 VSS.t520 41.4291
R6360 VSS.n494 VSS.t54 41.4291
R6361 VSS.n812 VSS.t130 41.4291
R6362 VSS.n1130 VSS.t33 41.4291
R6363 VSS.n1371 VSS.t250 41.4291
R6364 VSS.n1916 VSS.t469 41.4291
R6365 VSS.n1815 VSS.t677 41.4291
R6366 VSS.n1714 VSS.t213 41.4291
R6367 VSS.n1613 VSS.t44 41.4291
R6368 VSS.n1512 VSS.t552 41.4291
R6369 VSS.n4210 VSS.t244 41.4291
R6370 VSS.n3470 VSS.t307 41.4291
R6371 VSS.n3584 VSS.t289 41.4291
R6372 VSS.n3698 VSS.t108 41.4291
R6373 VSS.n3812 VSS.t207 41.4291
R6374 VSS.n72 VSS.t529 41.4198
R6375 VSS.n1140 VSS.n1139 40.5593
R6376 VSS.n1124 VSS.n1123 40.5593
R6377 VSS.n1110 VSS.n1109 40.5593
R6378 VSS.n1096 VSS.n1095 40.5593
R6379 VSS.n1082 VSS.n1081 40.5593
R6380 VSS.n1068 VSS.n1067 40.5593
R6381 VSS.n1040 VSS.n1039 40.5593
R6382 VSS.n1026 VSS.n1025 40.5593
R6383 VSS.n1012 VSS.n1011 40.5593
R6384 VSS.n998 VSS.n997 40.5593
R6385 VSS.n982 VSS.n981 40.5593
R6386 VSS.n968 VSS.n967 40.5593
R6387 VSS.n954 VSS.n953 40.5593
R6388 VSS.n156 VSS.n155 40.5593
R6389 VSS.n937 VSS.n936 40.5593
R6390 VSS.n166 VSS.n165 40.5593
R6391 VSS.n915 VSS.n914 40.5593
R6392 VSS.n916 VSS.n911 40.5593
R6393 VSS.n895 VSS.n894 40.5593
R6394 VSS.n881 VSS.n880 40.5593
R6395 VSS.n192 VSS.n191 40.5593
R6396 VSS.n864 VSS.n863 40.5593
R6397 VSS.n850 VSS.n849 40.5593
R6398 VSS.n836 VSS.n835 40.5593
R6399 VSS.n822 VSS.n821 40.5593
R6400 VSS.n806 VSS.n805 40.5593
R6401 VSS.n792 VSS.n791 40.5593
R6402 VSS.n778 VSS.n777 40.5593
R6403 VSS.n764 VSS.n763 40.5593
R6404 VSS.n750 VSS.n749 40.5593
R6405 VSS.n722 VSS.n721 40.5593
R6406 VSS.n708 VSS.n707 40.5593
R6407 VSS.n694 VSS.n693 40.5593
R6408 VSS.n680 VSS.n679 40.5593
R6409 VSS.n664 VSS.n663 40.5593
R6410 VSS.n650 VSS.n649 40.5593
R6411 VSS.n636 VSS.n635 40.5593
R6412 VSS.n201 VSS.n200 40.5593
R6413 VSS.n619 VSS.n618 40.5593
R6414 VSS.n211 VSS.n210 40.5593
R6415 VSS.n597 VSS.n596 40.5593
R6416 VSS.n598 VSS.n593 40.5593
R6417 VSS.n577 VSS.n576 40.5593
R6418 VSS.n563 VSS.n562 40.5593
R6419 VSS.n237 VSS.n236 40.5593
R6420 VSS.n546 VSS.n545 40.5593
R6421 VSS.n532 VSS.n531 40.5593
R6422 VSS.n518 VSS.n517 40.5593
R6423 VSS.n504 VSS.n503 40.5593
R6424 VSS.n488 VSS.n487 40.5593
R6425 VSS.n474 VSS.n473 40.5593
R6426 VSS.n460 VSS.n459 40.5593
R6427 VSS.n446 VSS.n445 40.5593
R6428 VSS.n432 VSS.n431 40.5593
R6429 VSS.n404 VSS.n403 40.5593
R6430 VSS.n390 VSS.n389 40.5593
R6431 VSS.n376 VSS.n375 40.5593
R6432 VSS.n362 VSS.n361 40.5593
R6433 VSS.n346 VSS.n345 40.5593
R6434 VSS.n332 VSS.n331 40.5593
R6435 VSS.n318 VSS.n317 40.5593
R6436 VSS.n246 VSS.n245 40.5593
R6437 VSS.n301 VSS.n300 40.5593
R6438 VSS.n256 VSS.n255 40.5593
R6439 VSS.n280 VSS.n279 40.5593
R6440 VSS.n2168 VSS.n2167 40.5593
R6441 VSS.n2182 VSS.n2181 40.5593
R6442 VSS.n2196 VSS.n2195 40.5593
R6443 VSS.n2212 VSS.n2211 40.5593
R6444 VSS.n2226 VSS.n2225 40.5593
R6445 VSS.n2240 VSS.n2239 40.5593
R6446 VSS.n2254 VSS.n2253 40.5593
R6447 VSS.n2268 VSS.n2267 40.5593
R6448 VSS.n2295 VSS.n2294 40.5593
R6449 VSS.n2309 VSS.n2308 40.5593
R6450 VSS.n2327 VSS.n2326 40.5593
R6451 VSS.n2337 VSS.n2336 40.5593
R6452 VSS.n119 VSS.n118 40.5593
R6453 VSS.n2367 VSS.n2366 40.5593
R6454 VSS.n2393 VSS.n2392 40.5593
R6455 VSS.n2407 VSS.n2406 40.5593
R6456 VSS.n2421 VSS.n2420 40.5593
R6457 VSS.n2435 VSS.n2434 40.5593
R6458 VSS.n2450 VSS.n2449 40.5593
R6459 VSS.n2464 VSS.n2463 40.5593
R6460 VSS.n2478 VSS.n2477 40.5593
R6461 VSS.n2492 VSS.n2491 40.5593
R6462 VSS.n2520 VSS.n2519 40.5593
R6463 VSS.n2534 VSS.n2533 40.5593
R6464 VSS.n2548 VSS.n2547 40.5593
R6465 VSS.n2564 VSS.n2563 40.5593
R6466 VSS.n2578 VSS.n2577 40.5593
R6467 VSS.n2592 VSS.n2591 40.5593
R6468 VSS.n2606 VSS.n2605 40.5593
R6469 VSS.n2620 VSS.n2619 40.5593
R6470 VSS.n2647 VSS.n2646 40.5593
R6471 VSS.n2661 VSS.n2660 40.5593
R6472 VSS.n2679 VSS.n2678 40.5593
R6473 VSS.n2689 VSS.n2688 40.5593
R6474 VSS.n108 VSS.n107 40.5593
R6475 VSS.n2719 VSS.n2718 40.5593
R6476 VSS.n2745 VSS.n2744 40.5593
R6477 VSS.n2759 VSS.n2758 40.5593
R6478 VSS.n2773 VSS.n2772 40.5593
R6479 VSS.n2787 VSS.n2786 40.5593
R6480 VSS.n2802 VSS.n2801 40.5593
R6481 VSS.n2816 VSS.n2815 40.5593
R6482 VSS.n2830 VSS.n2829 40.5593
R6483 VSS.n2844 VSS.n2843 40.5593
R6484 VSS.n2872 VSS.n2871 40.5593
R6485 VSS.n2886 VSS.n2885 40.5593
R6486 VSS.n2900 VSS.n2899 40.5593
R6487 VSS.n2916 VSS.n2915 40.5593
R6488 VSS.n2930 VSS.n2929 40.5593
R6489 VSS.n2944 VSS.n2943 40.5593
R6490 VSS.n2958 VSS.n2957 40.5593
R6491 VSS.n2972 VSS.n2971 40.5593
R6492 VSS.n2999 VSS.n2998 40.5593
R6493 VSS.n3013 VSS.n3012 40.5593
R6494 VSS.n3031 VSS.n3030 40.5593
R6495 VSS.n94 VSS.n93 40.5593
R6496 VSS.n3045 VSS.n3044 40.5593
R6497 VSS.n3060 VSS.n3059 40.5593
R6498 VSS.n3074 VSS.n3073 40.5593
R6499 VSS.n84 VSS.n83 40.5593
R6500 VSS.n3314 VSS.n3313 40.5593
R6501 VSS.n3300 VSS.n3299 40.5593
R6502 VSS.n3284 VSS.n3283 40.5593
R6503 VSS.n3271 VSS.n3270 40.5593
R6504 VSS.n3255 VSS.n3254 40.5593
R6505 VSS.n3241 VSS.n3240 40.5593
R6506 VSS.n3226 VSS.n3225 40.5593
R6507 VSS.n3211 VSS.n3210 40.5593
R6508 VSS.n3197 VSS.n3196 40.5593
R6509 VSS.n3181 VSS.n3180 40.5593
R6510 VSS.n3167 VSS.n3166 40.5593
R6511 VSS.n3149 VSS.n3148 40.5593
R6512 VSS.n3135 VSS.n3134 40.5593
R6513 VSS.n3119 VSS.n3118 40.5593
R6514 VSS.n3105 VSS.n3104 40.5593
R6515 VSS.n3089 VSS.n3088 40.5593
R6516 VSS.n71 VSS.n70 40.5593
R6517 VSS.n64 VSS.n63 40.5593
R6518 VSS.n3972 VSS.t395 39.6928
R6519 VSS.n1998 VSS.t66 38.5719
R6520 VSS.n1998 VSS.t3 38.5719
R6521 VSS.n2022 VSS.t146 38.5719
R6522 VSS.n2061 VSS.t154 38.5719
R6523 VSS.n2113 VSS.t138 38.5719
R6524 VSS.n2113 VSS.t320 38.5719
R6525 VSS.n2137 VSS.t170 38.5719
R6526 VSS.n2207 VSS.t172 38.5719
R6527 VSS.n112 VSS.t597 38.5719
R6528 VSS.n112 VSS.t641 38.5719
R6529 VSS.n2440 VSS.t158 38.5719
R6530 VSS.n2559 VSS.t168 38.5719
R6531 VSS.n101 VSS.t140 38.5719
R6532 VSS.n101 VSS.t73 38.5719
R6533 VSS.n2792 VSS.t148 38.5719
R6534 VSS.n2911 VSS.t156 38.5719
R6535 VSS.n13 VSS.t382 38.5719
R6536 VSS.n13 VSS.t492 38.5719
R6537 VSS.n250 VSS.t377 38.5719
R6538 VSS.n250 VSS.t543 38.5719
R6539 VSS.n357 VSS.t631 38.5719
R6540 VSS.n494 VSS.t629 38.5719
R6541 VSS.n205 VSS.t572 38.5719
R6542 VSS.n205 VSS.t12 38.5719
R6543 VSS.n675 VSS.t234 38.5719
R6544 VSS.n812 VSS.t232 38.5719
R6545 VSS.n160 VSS.t62 38.5719
R6546 VSS.n160 VSS.t673 38.5719
R6547 VSS.n993 VSS.t490 38.5719
R6548 VSS.n1130 VSS.t488 38.5719
R6549 VSS.n1232 VSS.t238 38.5719
R6550 VSS.n1232 VSS.t496 38.5719
R6551 VSS.n1285 VSS.t92 38.5719
R6552 VSS.n1371 VSS.t94 38.5719
R6553 VSS.n1979 VSS.t274 38.5719
R6554 VSS.n1979 VSS.t282 38.5719
R6555 VSS.n1955 VSS.t681 38.5719
R6556 VSS.n1916 VSS.t683 38.5719
R6557 VSS.n1878 VSS.t195 38.5719
R6558 VSS.n1878 VSS.t500 38.5719
R6559 VSS.n1854 VSS.t581 38.5719
R6560 VSS.n1815 VSS.t583 38.5719
R6561 VSS.n1777 VSS.t380 38.5719
R6562 VSS.n1777 VSS.t296 38.5719
R6563 VSS.n1753 VSS.t593 38.5719
R6564 VSS.n1714 VSS.t591 38.5719
R6565 VSS.n1676 VSS.t387 38.5719
R6566 VSS.n1676 VSS.t199 38.5719
R6567 VSS.n1652 VSS.t358 38.5719
R6568 VSS.n1613 VSS.t360 38.5719
R6569 VSS.n1575 VSS.t595 38.5719
R6570 VSS.n1575 VSS.t504 38.5719
R6571 VSS.n1551 VSS.t114 38.5719
R6572 VSS.n1512 VSS.t116 38.5719
R6573 VSS.n4210 VSS.t162 38.5719
R6574 VSS.n4249 VSS.t164 38.5719
R6575 VSS.n7 VSS.t266 38.5719
R6576 VSS.n7 VSS.t589 38.5719
R6577 VSS.n3470 VSS.t152 38.5719
R6578 VSS.n3509 VSS.t166 38.5719
R6579 VSS.n3439 VSS.t655 38.5719
R6580 VSS.n3439 VSS.t415 38.5719
R6581 VSS.n3584 VSS.t144 38.5719
R6582 VSS.n3623 VSS.t150 38.5719
R6583 VSS.n3437 VSS.t685 38.5719
R6584 VSS.n3437 VSS.t417 38.5719
R6585 VSS.n3698 VSS.t174 38.5719
R6586 VSS.n3737 VSS.t142 38.5719
R6587 VSS.n3435 VSS.t276 38.5719
R6588 VSS.n3435 VSS.t64 38.5719
R6589 VSS.n3812 VSS.t435 38.5719
R6590 VSS.n3851 VSS.t90 38.5719
R6591 VSS.n3881 VSS.t482 38.5719
R6592 VSS.n3881 VSS.t643 38.5719
R6593 VSS.n2422 VSS.t457 35.2005
R6594 VSS.n2774 VSS.t418 35.2005
R6595 VSS.n1152 VSS.t286 34.3085
R6596 VSS.t60 VSS.n1098 34.3085
R6597 VSS.n837 VSS.t584 34.3085
R6598 VSS.t574 VSS.n780 34.3085
R6599 VSS.n519 VSS.t600 34.3085
R6600 VSS.t375 VSS.n462 34.3085
R6601 VSS.n3426 VSS.t193 33.462
R6602 VSS.n3426 VSS.t217 33.462
R6603 VSS.n3896 VSS.t526 33.462
R6604 VSS.n3896 VSS.t1 33.462
R6605 VSS.n3344 VSS.t570 33.462
R6606 VSS.n3344 VSS.t568 33.462
R6607 VSS.n3332 VSS.n3331 31.8615
R6608 VSS.n3317 VSS.n3316 31.8615
R6609 VSS.n3303 VSS.n3302 31.8615
R6610 VSS.n3273 VSS.t331 31.8615
R6611 VSS.n3258 VSS.n3257 31.8615
R6612 VSS.n3244 VSS.n3243 31.8615
R6613 VSS.n3229 VSS.n3228 31.8615
R6614 VSS.n3214 VSS.n3213 31.8615
R6615 VSS.n3200 VSS.n3199 31.8615
R6616 VSS.n3184 VSS.n3183 31.8615
R6617 VSS.n3170 VSS.n3169 31.8615
R6618 VSS.n3152 VSS.n3151 31.8615
R6619 VSS.n3152 VSS.t351 31.8615
R6620 VSS.n3138 VSS.n3137 31.8615
R6621 VSS.n3108 VSS.n3107 31.8615
R6622 VSS.n3092 VSS.n3091 31.8615
R6623 VSS.n3379 VSS.n73 31.8615
R6624 VSS.n3942 VSS.n3939 30.1954
R6625 VSS.n3939 VSS.n3936 30.1954
R6626 VSS.n3936 VSS.n3933 30.1954
R6627 VSS.n3933 VSS.n3930 30.1954
R6628 VSS.n3242 VSS.t327 28.6754
R6629 VSS.n4224 VSS.t125 26.8298
R6630 VSS.n3484 VSS.t463 26.8298
R6631 VSS.n3598 VSS.t385 26.8298
R6632 VSS.n3712 VSS.t477 26.8298
R6633 VSS.n3826 VSS.t671 26.8298
R6634 VSS.n1934 VSS.t450 26.3478
R6635 VSS.n1833 VSS.t36 26.3478
R6636 VSS.n1732 VSS.t103 26.3478
R6637 VSS.n1631 VSS.t123 26.3478
R6638 VSS.n1530 VSS.t222 26.3478
R6639 VSS.n3024 VSS.t128 25.9346
R6640 VSS.n2086 VSS.t443 25.9346
R6641 VSS.n2100 VSS.t9 25.9346
R6642 VSS.n2279 VSS.t21 25.9346
R6643 VSS.n2320 VSS.t96 25.9346
R6644 VSS.n2631 VSS.t413 25.9346
R6645 VSS.n2672 VSS.t49 25.9346
R6646 VSS.n2983 VSS.t516 25.9346
R6647 VSS.n231 VSS.t58 25.9346
R6648 VSS.n229 VSS.t69 25.9346
R6649 VSS.n186 VSS.t134 25.9346
R6650 VSS.n184 VSS.t445 25.9346
R6651 VSS.n1188 VSS.t31 25.9346
R6652 VSS.n149 VSS.t626 25.9346
R6653 VSS.n131 VSS.t248 25.9346
R6654 VSS.n126 VSS.t603 25.9346
R6655 VSS.n1415 VSS.t465 25.9346
R6656 VSS.n1420 VSS.t71 25.9346
R6657 VSS.n1430 VSS.t679 25.9346
R6658 VSS.n1435 VSS.t203 25.9346
R6659 VSS.n1445 VSS.t215 25.9346
R6660 VSS.n1450 VSS.t313 25.9346
R6661 VSS.n1460 VSS.t46 25.9346
R6662 VSS.n1465 VSS.t691 25.9346
R6663 VSS.n1475 VSS.t554 25.9346
R6664 VSS.n1480 VSS.t637 25.9346
R6665 VSS.n4191 VSS.t242 25.9346
R6666 VSS.n4 VSS.t221 25.9346
R6667 VSS.n3451 VSS.t311 25.9346
R6668 VSS.n3551 VSS.t431 25.9346
R6669 VSS.n3565 VSS.t293 25.9346
R6670 VSS.n3665 VSS.t667 25.9346
R6671 VSS.n3679 VSS.t112 25.9346
R6672 VSS.n3779 VSS.t665 25.9346
R6673 VSS.n3793 VSS.t205 25.9346
R6674 VSS.n4177 VSS.t437 25.9346
R6675 VSS.n2379 VSS.n2378 25.7776
R6676 VSS.n2731 VSS.n2730 25.7776
R6677 VSS.n1053 VSS.n1052 25.7735
R6678 VSS.n735 VSS.n734 25.7735
R6679 VSS.n417 VSS.n416 25.7735
R6680 VSS.n2505 VSS.n2504 25.7735
R6681 VSS.n2857 VSS.n2856 25.7735
R6682 VSS.n2281 VSS.n2280 25.7735
R6683 VSS.n114 VSS.n113 25.7735
R6684 VSS.n2633 VSS.n2632 25.7735
R6685 VSS.n103 VSS.n102 25.7735
R6686 VSS.n2985 VSS.n2984 25.7735
R6687 VSS.n177 VSS.n176 25.765
R6688 VSS.n222 VSS.n221 25.765
R6689 VSS.n4168 VSS.n4167 25.7315
R6690 VSS.n4158 VSS.n4157 25.7315
R6691 VSS.n4139 VSS.n4138 25.7315
R6692 VSS.n4125 VSS.t508 25.7315
R6693 VSS.n21 VSS.n20 25.7315
R6694 VSS.n4109 VSS.n4108 25.7315
R6695 VSS.n4110 VSS.t6 25.7315
R6696 VSS.n4097 VSS.n4096 25.7315
R6697 VSS.n4083 VSS.n4082 25.7315
R6698 VSS.n4069 VSS.n4068 25.7315
R6699 VSS.n33 VSS.n32 25.7315
R6700 VSS.n4052 VSS.n4051 25.7315
R6701 VSS.n4040 VSS.n4039 25.7315
R6702 VSS.n4026 VSS.n4025 25.7315
R6703 VSS.n4012 VSS.n4011 25.7315
R6704 VSS.n3997 VSS.n3996 25.7315
R6705 VSS.n3983 VSS.n3982 25.7315
R6706 VSS.n3968 VSS.n3967 25.7315
R6707 VSS.n3954 VSS.n3953 25.7315
R6708 VSS.n47 VSS.n46 25.7315
R6709 VSS.n1127 VSS.t487 25.7315
R6710 VSS.n809 VSS.t231 25.7315
R6711 VSS.n491 VSS.t628 25.7315
R6712 VSS.n77 VSS.t398 25.7315
R6713 VSS.t353 VSS.n3286 25.4893
R6714 VSS.n3930 VSS.n3927 25.2497
R6715 VSS.n4001 VSS.t391 24.9241
R6716 VSS.n3402 VSS.t566 24.9236
R6717 VSS.n3402 VSS.t562 24.9236
R6718 VSS.n3409 VSS.t564 24.9236
R6719 VSS.n3409 VSS.t622 24.9236
R6720 VSS.n85 VSS.t338 24.9236
R6721 VSS.n85 VSS.t356 24.9236
R6722 VSS.n3320 VSS.t346 24.9236
R6723 VSS.n3320 VSS.t340 24.9236
R6724 VSS.n3290 VSS.t354 24.9236
R6725 VSS.n3290 VSS.t332 24.9236
R6726 VSS.n3261 VSS.t350 24.9236
R6727 VSS.n3261 VSS.t328 24.9236
R6728 VSS.n3222 VSS.t348 24.9236
R6729 VSS.n3222 VSS.t336 24.9236
R6730 VSS.n3192 VSS.t344 24.9236
R6731 VSS.n3192 VSS.t334 24.9236
R6732 VSS.n3162 VSS.t342 24.9236
R6733 VSS.n3162 VSS.t330 24.9236
R6734 VSS.n3155 VSS.t352 24.9236
R6735 VSS.n3155 VSS.t534 24.9236
R6736 VSS.n3125 VSS.t540 24.9236
R6737 VSS.n3125 VSS.t532 24.9236
R6738 VSS.n3095 VSS.t538 24.9236
R6739 VSS.n3095 VSS.t530 24.9236
R6740 VSS.n3972 VSS.t393 24.9236
R6741 VSS.n3920 VSS.t183 24.9236
R6742 VSS.n3920 VSS.t177 24.9236
R6743 VSS.n3907 VSS.t181 24.9236
R6744 VSS.n3907 VSS.t524 24.9236
R6745 VSS.n3366 VSS.t663 24.9236
R6746 VSS.n3366 VSS.t657 24.9236
R6747 VSS.n3356 VSS.t661 24.9236
R6748 VSS.n3356 VSS.t433 24.9236
R6749 VSS.n3316 VSS.n3315 22.3032
R6750 VSS.n3302 VSS.n3301 22.3032
R6751 VSS.n3286 VSS.n3285 22.3032
R6752 VSS.t331 VSS.n3272 22.3032
R6753 VSS.n3257 VSS.n3256 22.3032
R6754 VSS.n3243 VSS.n3242 22.3032
R6755 VSS.n3228 VSS.n3227 22.3032
R6756 VSS.n3213 VSS.n3212 22.3032
R6757 VSS.n3199 VSS.n3198 22.3032
R6758 VSS.n3183 VSS.n3182 22.3032
R6759 VSS.n3169 VSS.n3168 22.3032
R6760 VSS.n3151 VSS.n3150 22.3032
R6761 VSS.n3137 VSS.n3136 22.3032
R6762 VSS.n3121 VSS.n3120 22.3032
R6763 VSS.n3091 VSS.n3090 22.3032
R6764 VSS.n73 VSS.n72 22.3032
R6765 VSS.n2107 VSS.n2106 20.3039
R6766 VSS.n1888 VSS.n1885 20.3039
R6767 VSS.n1787 VSS.n1784 20.3039
R6768 VSS.n1686 VSS.n1683 20.3039
R6769 VSS.n1585 VSS.n1582 20.3039
R6770 VSS.n3333 VSS.n3332 19.1171
R6771 VSS.n3303 VSS.t339 19.1171
R6772 VSS.n3122 VSS.t539 19.1171
R6773 VSS.n2049 VSS.t476 17.6005
R6774 VSS.n4156 VSS.n4155 17.3829
R6775 VSS.n4137 VSS.n4136 17.3829
R6776 VSS.n4124 VSS.n4123 17.3829
R6777 VSS.n19 VSS.n18 17.3829
R6778 VSS.n4107 VSS.n4106 17.3829
R6779 VSS.n4095 VSS.n4094 17.3829
R6780 VSS.n4081 VSS.n4080 17.3829
R6781 VSS.n4067 VSS.n4066 17.3829
R6782 VSS.n31 VSS.n30 17.3829
R6783 VSS.n4050 VSS.n4049 17.3829
R6784 VSS.n4038 VSS.n4037 17.3829
R6785 VSS.n4024 VSS.n4023 17.3829
R6786 VSS.n4010 VSS.n4009 17.3829
R6787 VSS.n3995 VSS.n3994 17.3829
R6788 VSS.n3981 VSS.n3980 17.3829
R6789 VSS.n3966 VSS.n3965 17.3829
R6790 VSS.n3952 VSS.n3951 17.3829
R6791 VSS.n45 VSS.n44 17.3829
R6792 VSS.n4164 VSS.n12 17.2298
R6793 VSS.n4070 VSS.t226 17.1545
R6794 VSS.n1353 VSS.t494 17.1545
R6795 VSS.n3421 VSS 16.7729
R6796 VSS.n3900 VSS 16.7729
R6797 VSS.n4286 VSS 16.7729
R6798 VSS.n3546 VSS 16.7729
R6799 VSS.n3660 VSS 16.7729
R6800 VSS.n3774 VSS 16.7729
R6801 VSS.n3090 VSS.t537 15.931
R6802 VSS.n3943 VSS.n3942 15.3978
R6803 VSS.n3396 VSS.n56 14.3453
R6804 VSS.n3348 VSS 14.0991
R6805 VSS.n4241 VSS.t369 13.4151
R6806 VSS.n4283 VSS 13.4151
R6807 VSS.n3501 VSS.t324 13.4151
R6808 VSS.n3543 VSS 13.4151
R6809 VSS.n3615 VSS.t635 13.4151
R6810 VSS.n3657 VSS 13.4151
R6811 VSS.n3729 VSS.t47 13.4151
R6812 VSS.n3771 VSS 13.4151
R6813 VSS.n3843 VSS.t106 13.4151
R6814 VSS.n3887 VSS 13.4151
R6815 VSS.n178 VSS.n177 13.0096
R6816 VSS.n223 VSS.n222 13.0096
R6817 VSS.n2282 VSS.n2281 13.0005
R6818 VSS.n115 VSS.n114 13.0005
R6819 VSS.n2634 VSS.n2633 13.0005
R6820 VSS.n104 VSS.n103 13.0005
R6821 VSS.n2986 VSS.n2985 13.0005
R6822 VSS.n2506 VSS.n2505 13.0005
R6823 VSS.n2858 VSS.n2857 13.0005
R6824 VSS.n418 VSS.n417 13.0005
R6825 VSS.n736 VSS.n735 13.0005
R6826 VSS.n1054 VSS.n1053 13.0005
R6827 VSS.n2380 VSS.n2379 12.9961
R6828 VSS.n2732 VSS.n2731 12.9961
R6829 VSS.n2344 VSS.n2343 12.8005
R6830 VSS.n2696 VSS.n2695 12.8005
R6831 VSS.n3042 VSS.n3041 12.8005
R6832 VSS.n3052 VSS.n3051 12.8005
R6833 VSS.t539 VSS.n3121 12.7449
R6834 VSS.n3107 VSS.t531 12.7449
R6835 VSS VSS.n287 12.5798
R6836 VSS.n1885 VSS.n1880 12.5798
R6837 VSS.n1784 VSS.n1779 12.5798
R6838 VSS.n1683 VSS.n1678 12.5798
R6839 VSS.n1582 VSS.n1577 12.5798
R6840 VSS.n1986 VSS.n1981 12.5798
R6841 VSS.n12 VSS.n11 12.0275
R6842 VSS VSS.n607 11.035
R6843 VSS VSS.n925 11.035
R6844 VSS.n140 VSS 11.035
R6845 VSS.n261 VSS.n260 10.7116
R6846 VSS.n1930 VSS.t80 10.5394
R6847 VSS.n1829 VSS.t304 10.5394
R6848 VSS.n1728 VSS.t98 10.5394
R6849 VSS.n1627 VSS.t184 10.5394
R6850 VSS.n1526 VSS.t196 10.5394
R6851 VSS.n270 VSS.n269 9.6405
R6852 VSS.t531 VSS.n3106 9.55879
R6853 VSS.t535 VSS.n3378 9.3622
R6854 VSS.n50 VSS.n49 9.3005
R6855 VSS.n49 VSS.n48 9.3005
R6856 VSS.n3957 VSS.n3956 9.3005
R6857 VSS.n3956 VSS.n3955 9.3005
R6858 VSS.n3971 VSS.n3970 9.3005
R6859 VSS.n3970 VSS.n3969 9.3005
R6860 VSS.n3986 VSS.n3985 9.3005
R6861 VSS.n3985 VSS.n3984 9.3005
R6862 VSS.n4000 VSS.n3999 9.3005
R6863 VSS.n3999 VSS.n3998 9.3005
R6864 VSS.n4015 VSS.n4014 9.3005
R6865 VSS.n4014 VSS.n4013 9.3005
R6866 VSS.n4029 VSS.n4028 9.3005
R6867 VSS.n4028 VSS.n4027 9.3005
R6868 VSS.n4043 VSS.n4042 9.3005
R6869 VSS.n4042 VSS.n4041 9.3005
R6870 VSS.n4055 VSS.n4054 9.3005
R6871 VSS.n4054 VSS.n4053 9.3005
R6872 VSS.n36 VSS.n35 9.3005
R6873 VSS.n35 VSS.n34 9.3005
R6874 VSS.n4072 VSS.n4071 9.3005
R6875 VSS.n4071 VSS.n4070 9.3005
R6876 VSS.n4086 VSS.n4085 9.3005
R6877 VSS.n4085 VSS.n4084 9.3005
R6878 VSS.n4100 VSS.n4099 9.3005
R6879 VSS.n4099 VSS.n4098 9.3005
R6880 VSS.n4112 VSS.n4111 9.3005
R6881 VSS.n4111 VSS.n4110 9.3005
R6882 VSS.n26 VSS.n23 9.3005
R6883 VSS.n23 VSS.n22 9.3005
R6884 VSS.n4128 VSS.n4127 9.3005
R6885 VSS.n4127 VSS.n4126 9.3005
R6886 VSS.n4142 VSS.n4141 9.3005
R6887 VSS.n4141 VSS.n4140 9.3005
R6888 VSS.n4161 VSS.n4160 9.3005
R6889 VSS.n4160 VSS.n4159 9.3005
R6890 VSS.n4165 VSS.n4164 9.3005
R6891 VSS.n4166 VSS.n4165 9.3005
R6892 VSS.n3392 VSS.n3391 9.3005
R6893 VSS.n3393 VSS.n3392 9.3005
R6894 VSS.n3330 VSS.n3329 9.3005
R6895 VSS.n3331 VSS.n3330 9.3005
R6896 VSS.n3319 VSS.n3318 9.3005
R6897 VSS.n3318 VSS.n3317 9.3005
R6898 VSS.n3305 VSS.n3304 9.3005
R6899 VSS.n3304 VSS.n3303 9.3005
R6900 VSS.n3289 VSS.n3288 9.3005
R6901 VSS.n3288 VSS.n3287 9.3005
R6902 VSS.n3275 VSS.n3274 9.3005
R6903 VSS.n3274 VSS.n3273 9.3005
R6904 VSS.n3260 VSS.n3259 9.3005
R6905 VSS.n3259 VSS.n3258 9.3005
R6906 VSS.n3246 VSS.n3245 9.3005
R6907 VSS.n3245 VSS.n3244 9.3005
R6908 VSS.n3231 VSS.n3230 9.3005
R6909 VSS.n3230 VSS.n3229 9.3005
R6910 VSS.n3216 VSS.n3215 9.3005
R6911 VSS.n3215 VSS.n3214 9.3005
R6912 VSS.n3202 VSS.n3201 9.3005
R6913 VSS.n3201 VSS.n3200 9.3005
R6914 VSS.n3186 VSS.n3185 9.3005
R6915 VSS.n3185 VSS.n3184 9.3005
R6916 VSS.n3172 VSS.n3171 9.3005
R6917 VSS.n3171 VSS.n3170 9.3005
R6918 VSS.n3154 VSS.n3153 9.3005
R6919 VSS.n3153 VSS.n3152 9.3005
R6920 VSS.n3140 VSS.n3139 9.3005
R6921 VSS.n3139 VSS.n3138 9.3005
R6922 VSS.n3124 VSS.n3123 9.3005
R6923 VSS.n3123 VSS.n3122 9.3005
R6924 VSS.n3110 VSS.n3109 9.3005
R6925 VSS.n3109 VSS.n3108 9.3005
R6926 VSS.n3094 VSS.n3093 9.3005
R6927 VSS.n3093 VSS.n3092 9.3005
R6928 VSS.n3381 VSS.n3380 9.3005
R6929 VSS.n3380 VSS.n3379 9.3005
R6930 VSS.n1365 VSS.n1364 9.3005
R6931 VSS.n1364 VSS.n1363 9.3005
R6932 VSS.n1355 VSS.n1354 9.3005
R6933 VSS.n1354 VSS.n1353 9.3005
R6934 VSS.n1335 VSS.n1334 9.3005
R6935 VSS.n1334 VSS.n1333 9.3005
R6936 VSS.n1325 VSS.n1324 9.3005
R6937 VSS.n1324 VSS.n1323 9.3005
R6938 VSS.n1315 VSS.n1314 9.3005
R6939 VSS.n1314 VSS.n1313 9.3005
R6940 VSS.n1295 VSS.n1294 9.3005
R6941 VSS.n1294 VSS.n1293 9.3005
R6942 VSS.n1283 VSS.n1282 9.3005
R6943 VSS.n1282 VSS.n1281 9.3005
R6944 VSS.n1273 VSS.n1272 9.3005
R6945 VSS.n1272 VSS.n1271 9.3005
R6946 VSS.n1246 VSS.n1245 9.3005
R6947 VSS.n1243 VSS.n1242 9.3005
R6948 VSS.n1242 VSS.n1241 9.3005
R6949 VSS.n1225 VSS.n1224 9.3005
R6950 VSS.n1215 VSS.n1214 9.3005
R6951 VSS.n1214 VSS.n1213 9.3005
R6952 VSS.n148 VSS.n147 9.3005
R6953 VSS.n147 VSS.n146 9.3005
R6954 VSS.n1209 VSS.n1208 9.3005
R6955 VSS.n1208 VSS.n1207 9.3005
R6956 VSS.n1181 VSS.n1180 9.3005
R6957 VSS.n1178 VSS.n1177 9.3005
R6958 VSS.n1177 VSS.n1176 9.3005
R6959 VSS.n1168 VSS.n1167 9.3005
R6960 VSS.n1167 VSS.n1166 9.3005
R6961 VSS.n1145 VSS.n1144 9.3005
R6962 VSS.n1144 VSS.n1143 9.3005
R6963 VSS.n1129 VSS.n1128 9.3005
R6964 VSS.n1128 VSS.n1127 9.3005
R6965 VSS.n1115 VSS.n1114 9.3005
R6966 VSS.n1114 VSS.n1113 9.3005
R6967 VSS.n1101 VSS.n1100 9.3005
R6968 VSS.n1100 VSS.n1099 9.3005
R6969 VSS.n1087 VSS.n1086 9.3005
R6970 VSS.n1086 VSS.n1085 9.3005
R6971 VSS.n1073 VSS.n1072 9.3005
R6972 VSS.n1072 VSS.n1071 9.3005
R6973 VSS.n1059 VSS.n1058 9.3005
R6974 VSS.n1058 VSS.n1057 9.3005
R6975 VSS.n1045 VSS.n1044 9.3005
R6976 VSS.n1044 VSS.n1043 9.3005
R6977 VSS.n1031 VSS.n1030 9.3005
R6978 VSS.n1030 VSS.n1029 9.3005
R6979 VSS.n1017 VSS.n1016 9.3005
R6980 VSS.n1016 VSS.n1015 9.3005
R6981 VSS.n1003 VSS.n1002 9.3005
R6982 VSS.n1002 VSS.n1001 9.3005
R6983 VSS.n987 VSS.n986 9.3005
R6984 VSS.n986 VSS.n985 9.3005
R6985 VSS.n973 VSS.n972 9.3005
R6986 VSS.n972 VSS.n971 9.3005
R6987 VSS.n959 VSS.n958 9.3005
R6988 VSS.n958 VSS.n957 9.3005
R6989 VSS.n154 VSS.n153 9.3005
R6990 VSS.n942 VSS.n941 9.3005
R6991 VSS.n941 VSS.n940 9.3005
R6992 VSS.n164 VSS.n163 9.3005
R6993 VSS.n917 VSS.n173 9.3005
R6994 VSS.n918 VSS.n917 9.3005
R6995 VSS.n923 VSS.n922 9.3005
R6996 VSS.n922 VSS.n921 9.3005
R6997 VSS.n183 VSS.n182 9.3005
R6998 VSS.n182 VSS.n181 9.3005
R6999 VSS.n900 VSS.n899 9.3005
R7000 VSS.n899 VSS.n898 9.3005
R7001 VSS.n886 VSS.n885 9.3005
R7002 VSS.n885 VSS.n884 9.3005
R7003 VSS.n190 VSS.n189 9.3005
R7004 VSS.n869 VSS.n868 9.3005
R7005 VSS.n868 VSS.n867 9.3005
R7006 VSS.n855 VSS.n854 9.3005
R7007 VSS.n854 VSS.n853 9.3005
R7008 VSS.n841 VSS.n840 9.3005
R7009 VSS.n840 VSS.n839 9.3005
R7010 VSS.n827 VSS.n826 9.3005
R7011 VSS.n826 VSS.n825 9.3005
R7012 VSS.n811 VSS.n810 9.3005
R7013 VSS.n810 VSS.n809 9.3005
R7014 VSS.n797 VSS.n796 9.3005
R7015 VSS.n796 VSS.n795 9.3005
R7016 VSS.n783 VSS.n782 9.3005
R7017 VSS.n782 VSS.n781 9.3005
R7018 VSS.n769 VSS.n768 9.3005
R7019 VSS.n768 VSS.n767 9.3005
R7020 VSS.n755 VSS.n754 9.3005
R7021 VSS.n754 VSS.n753 9.3005
R7022 VSS.n741 VSS.n740 9.3005
R7023 VSS.n740 VSS.n739 9.3005
R7024 VSS.n727 VSS.n726 9.3005
R7025 VSS.n726 VSS.n725 9.3005
R7026 VSS.n713 VSS.n712 9.3005
R7027 VSS.n712 VSS.n711 9.3005
R7028 VSS.n699 VSS.n698 9.3005
R7029 VSS.n698 VSS.n697 9.3005
R7030 VSS.n685 VSS.n684 9.3005
R7031 VSS.n684 VSS.n683 9.3005
R7032 VSS.n669 VSS.n668 9.3005
R7033 VSS.n668 VSS.n667 9.3005
R7034 VSS.n655 VSS.n654 9.3005
R7035 VSS.n654 VSS.n653 9.3005
R7036 VSS.n641 VSS.n640 9.3005
R7037 VSS.n640 VSS.n639 9.3005
R7038 VSS.n199 VSS.n198 9.3005
R7039 VSS.n624 VSS.n623 9.3005
R7040 VSS.n623 VSS.n622 9.3005
R7041 VSS.n209 VSS.n208 9.3005
R7042 VSS.n599 VSS.n218 9.3005
R7043 VSS.n600 VSS.n599 9.3005
R7044 VSS.n605 VSS.n604 9.3005
R7045 VSS.n604 VSS.n603 9.3005
R7046 VSS.n228 VSS.n227 9.3005
R7047 VSS.n227 VSS.n226 9.3005
R7048 VSS.n582 VSS.n581 9.3005
R7049 VSS.n581 VSS.n580 9.3005
R7050 VSS.n568 VSS.n567 9.3005
R7051 VSS.n567 VSS.n566 9.3005
R7052 VSS.n235 VSS.n234 9.3005
R7053 VSS.n551 VSS.n550 9.3005
R7054 VSS.n550 VSS.n549 9.3005
R7055 VSS.n537 VSS.n536 9.3005
R7056 VSS.n536 VSS.n535 9.3005
R7057 VSS.n523 VSS.n522 9.3005
R7058 VSS.n522 VSS.n521 9.3005
R7059 VSS.n509 VSS.n508 9.3005
R7060 VSS.n508 VSS.n507 9.3005
R7061 VSS.n493 VSS.n492 9.3005
R7062 VSS.n492 VSS.n491 9.3005
R7063 VSS.n479 VSS.n478 9.3005
R7064 VSS.n478 VSS.n477 9.3005
R7065 VSS.n465 VSS.n464 9.3005
R7066 VSS.n464 VSS.n463 9.3005
R7067 VSS.n451 VSS.n450 9.3005
R7068 VSS.n450 VSS.n449 9.3005
R7069 VSS.n437 VSS.n436 9.3005
R7070 VSS.n436 VSS.n435 9.3005
R7071 VSS.n423 VSS.n422 9.3005
R7072 VSS.n422 VSS.n421 9.3005
R7073 VSS.n409 VSS.n408 9.3005
R7074 VSS.n408 VSS.n407 9.3005
R7075 VSS.n395 VSS.n394 9.3005
R7076 VSS.n394 VSS.n393 9.3005
R7077 VSS.n381 VSS.n380 9.3005
R7078 VSS.n380 VSS.n379 9.3005
R7079 VSS.n367 VSS.n366 9.3005
R7080 VSS.n366 VSS.n365 9.3005
R7081 VSS.n351 VSS.n350 9.3005
R7082 VSS.n350 VSS.n349 9.3005
R7083 VSS.n337 VSS.n336 9.3005
R7084 VSS.n336 VSS.n335 9.3005
R7085 VSS.n323 VSS.n322 9.3005
R7086 VSS.n322 VSS.n321 9.3005
R7087 VSS.n244 VSS.n243 9.3005
R7088 VSS.n306 VSS.n305 9.3005
R7089 VSS.n305 VSS.n304 9.3005
R7090 VSS.n254 VSS.n253 9.3005
R7091 VSS.n281 VSS.n277 9.3005
R7092 VSS.n284 VSS.n281 9.3005
R7093 VSS.n1158 VSS.n1157 9.3005
R7094 VSS.n1157 VSS.n1156 9.3005
R7095 VSS.n1199 VSS.n1198 9.3005
R7096 VSS.n1198 VSS.n1197 9.3005
R7097 VSS.n1222 VSS.n1221 9.3005
R7098 VSS.n1221 VSS.n1220 9.3005
R7099 VSS.n1263 VSS.n1262 9.3005
R7100 VSS.n1262 VSS.n1261 9.3005
R7101 VSS.n1305 VSS.n1304 9.3005
R7102 VSS.n1304 VSS.n1303 9.3005
R7103 VSS.n1345 VSS.n1344 9.3005
R7104 VSS.n1344 VSS.n1343 9.3005
R7105 VSS.n2173 VSS.n2172 9.3005
R7106 VSS.n2172 VSS.n2171 9.3005
R7107 VSS.n2187 VSS.n2186 9.3005
R7108 VSS.n2186 VSS.n2185 9.3005
R7109 VSS.n2201 VSS.n2200 9.3005
R7110 VSS.n2200 VSS.n2199 9.3005
R7111 VSS.n2217 VSS.n2216 9.3005
R7112 VSS.n2216 VSS.n2215 9.3005
R7113 VSS.n2231 VSS.n2230 9.3005
R7114 VSS.n2230 VSS.n2229 9.3005
R7115 VSS.n2245 VSS.n2244 9.3005
R7116 VSS.n2244 VSS.n2243 9.3005
R7117 VSS.n2259 VSS.n2258 9.3005
R7118 VSS.n2258 VSS.n2257 9.3005
R7119 VSS.n2273 VSS.n2272 9.3005
R7120 VSS.n2272 VSS.n2271 9.3005
R7121 VSS.n2287 VSS.n2286 9.3005
R7122 VSS.n2286 VSS.n2285 9.3005
R7123 VSS.n2300 VSS.n2299 9.3005
R7124 VSS.n2299 VSS.n2298 9.3005
R7125 VSS.n2314 VSS.n2313 9.3005
R7126 VSS.n2313 VSS.n2312 9.3005
R7127 VSS.n2325 VSS.n2324 9.3005
R7128 VSS.n2342 VSS.n2341 9.3005
R7129 VSS.n2341 VSS.n2340 9.3005
R7130 VSS.n2353 VSS.n2352 9.3005
R7131 VSS.n2354 VSS.n2353 9.3005
R7132 VSS.n2359 VSS.n2358 9.3005
R7133 VSS.n2358 VSS.n2357 9.3005
R7134 VSS.n2372 VSS.n2371 9.3005
R7135 VSS.n2371 VSS.n2370 9.3005
R7136 VSS.n2385 VSS.n2384 9.3005
R7137 VSS.n2384 VSS.n2383 9.3005
R7138 VSS.n2398 VSS.n2397 9.3005
R7139 VSS.n2397 VSS.n2396 9.3005
R7140 VSS.n2412 VSS.n2411 9.3005
R7141 VSS.n2411 VSS.n2410 9.3005
R7142 VSS.n2426 VSS.n2425 9.3005
R7143 VSS.n2425 VSS.n2424 9.3005
R7144 VSS.n2439 VSS.n2438 9.3005
R7145 VSS.n2438 VSS.n2437 9.3005
R7146 VSS.n2455 VSS.n2454 9.3005
R7147 VSS.n2454 VSS.n2453 9.3005
R7148 VSS.n2469 VSS.n2468 9.3005
R7149 VSS.n2468 VSS.n2467 9.3005
R7150 VSS.n2483 VSS.n2482 9.3005
R7151 VSS.n2482 VSS.n2481 9.3005
R7152 VSS.n2497 VSS.n2496 9.3005
R7153 VSS.n2496 VSS.n2495 9.3005
R7154 VSS.n2511 VSS.n2510 9.3005
R7155 VSS.n2510 VSS.n2509 9.3005
R7156 VSS.n2525 VSS.n2524 9.3005
R7157 VSS.n2524 VSS.n2523 9.3005
R7158 VSS.n2539 VSS.n2538 9.3005
R7159 VSS.n2538 VSS.n2537 9.3005
R7160 VSS.n2553 VSS.n2552 9.3005
R7161 VSS.n2552 VSS.n2551 9.3005
R7162 VSS.n2569 VSS.n2568 9.3005
R7163 VSS.n2568 VSS.n2567 9.3005
R7164 VSS.n2583 VSS.n2582 9.3005
R7165 VSS.n2582 VSS.n2581 9.3005
R7166 VSS.n2597 VSS.n2596 9.3005
R7167 VSS.n2596 VSS.n2595 9.3005
R7168 VSS.n2611 VSS.n2610 9.3005
R7169 VSS.n2610 VSS.n2609 9.3005
R7170 VSS.n2625 VSS.n2624 9.3005
R7171 VSS.n2624 VSS.n2623 9.3005
R7172 VSS.n2639 VSS.n2638 9.3005
R7173 VSS.n2638 VSS.n2637 9.3005
R7174 VSS.n2652 VSS.n2651 9.3005
R7175 VSS.n2651 VSS.n2650 9.3005
R7176 VSS.n2666 VSS.n2665 9.3005
R7177 VSS.n2665 VSS.n2664 9.3005
R7178 VSS.n2677 VSS.n2676 9.3005
R7179 VSS.n2694 VSS.n2693 9.3005
R7180 VSS.n2693 VSS.n2692 9.3005
R7181 VSS.n2705 VSS.n2704 9.3005
R7182 VSS.n2706 VSS.n2705 9.3005
R7183 VSS.n2711 VSS.n2710 9.3005
R7184 VSS.n2710 VSS.n2709 9.3005
R7185 VSS.n2724 VSS.n2723 9.3005
R7186 VSS.n2723 VSS.n2722 9.3005
R7187 VSS.n2737 VSS.n2736 9.3005
R7188 VSS.n2736 VSS.n2735 9.3005
R7189 VSS.n2750 VSS.n2749 9.3005
R7190 VSS.n2749 VSS.n2748 9.3005
R7191 VSS.n2764 VSS.n2763 9.3005
R7192 VSS.n2763 VSS.n2762 9.3005
R7193 VSS.n2778 VSS.n2777 9.3005
R7194 VSS.n2777 VSS.n2776 9.3005
R7195 VSS.n2791 VSS.n2790 9.3005
R7196 VSS.n2790 VSS.n2789 9.3005
R7197 VSS.n2807 VSS.n2806 9.3005
R7198 VSS.n2806 VSS.n2805 9.3005
R7199 VSS.n2821 VSS.n2820 9.3005
R7200 VSS.n2820 VSS.n2819 9.3005
R7201 VSS.n2835 VSS.n2834 9.3005
R7202 VSS.n2834 VSS.n2833 9.3005
R7203 VSS.n2849 VSS.n2848 9.3005
R7204 VSS.n2848 VSS.n2847 9.3005
R7205 VSS.n2863 VSS.n2862 9.3005
R7206 VSS.n2862 VSS.n2861 9.3005
R7207 VSS.n2877 VSS.n2876 9.3005
R7208 VSS.n2876 VSS.n2875 9.3005
R7209 VSS.n2891 VSS.n2890 9.3005
R7210 VSS.n2890 VSS.n2889 9.3005
R7211 VSS.n2905 VSS.n2904 9.3005
R7212 VSS.n2904 VSS.n2903 9.3005
R7213 VSS.n2921 VSS.n2920 9.3005
R7214 VSS.n2920 VSS.n2919 9.3005
R7215 VSS.n2935 VSS.n2934 9.3005
R7216 VSS.n2934 VSS.n2933 9.3005
R7217 VSS.n2949 VSS.n2948 9.3005
R7218 VSS.n2948 VSS.n2947 9.3005
R7219 VSS.n2963 VSS.n2962 9.3005
R7220 VSS.n2962 VSS.n2961 9.3005
R7221 VSS.n2977 VSS.n2976 9.3005
R7222 VSS.n2976 VSS.n2975 9.3005
R7223 VSS.n2991 VSS.n2990 9.3005
R7224 VSS.n2990 VSS.n2989 9.3005
R7225 VSS.n3004 VSS.n3003 9.3005
R7226 VSS.n3003 VSS.n3002 9.3005
R7227 VSS.n3018 VSS.n3017 9.3005
R7228 VSS.n3017 VSS.n3016 9.3005
R7229 VSS.n3029 VSS.n3028 9.3005
R7230 VSS.n99 VSS.n98 9.3005
R7231 VSS.n98 VSS.n97 9.3005
R7232 VSS.n3050 VSS.n3049 9.3005
R7233 VSS.n3049 VSS.n3048 9.3005
R7234 VSS.n3065 VSS.n3064 9.3005
R7235 VSS.n3064 VSS.n3063 9.3005
R7236 VSS.n3079 VSS.n3078 9.3005
R7237 VSS.n3078 VSS.n3077 9.3005
R7238 VSS.n2026 VSS.n2023 9.04877
R7239 VSS.n2141 VSS.n2138 9.04877
R7240 VSS.n3336 VSS.n81 9.04877
R7241 VSS.n1959 VSS.n1956 9.04877
R7242 VSS.n1858 VSS.n1855 9.04877
R7243 VSS.n1757 VSS.n1754 9.04877
R7244 VSS.n1656 VSS.n1653 9.04877
R7245 VSS.n1555 VSS.n1552 9.04877
R7246 VSS.n4253 VSS.n4250 9.04877
R7247 VSS.n3513 VSS.n3510 9.04877
R7248 VSS.n3627 VSS.n3624 9.04877
R7249 VSS.n3741 VSS.n3738 9.04877
R7250 VSS.n3855 VSS.n3852 9.04877
R7251 VSS.n3 VSS.n2 9.01861
R7252 VSS.n3550 VSS.n3549 9.01861
R7253 VSS.n3664 VSS.n3663 9.01861
R7254 VSS.n3778 VSS.n3777 9.01861
R7255 VSS.n3919 VSS.n3918 9.01832
R7256 VSS.n4176 VSS.n4175 9.01761
R7257 VSS.n3895 VSS.n3894 9.01734
R7258 VSS.n4190 VSS.n4189 9.01732
R7259 VSS.n4279 VSS.n4278 9.01732
R7260 VSS.n3450 VSS.n3449 9.01732
R7261 VSS.n3541 VSS.n3540 9.01732
R7262 VSS.n3564 VSS.n3563 9.01732
R7263 VSS.n3655 VSS.n3654 9.01732
R7264 VSS.n3678 VSS.n3677 9.01732
R7265 VSS.n3769 VSS.n3768 9.01732
R7266 VSS.n3792 VSS.n3791 9.01732
R7267 VSS.n3880 VSS.n3879 9.01732
R7268 VSS.n4269 VSS.n4268 9.01719
R7269 VSS.n3529 VSS.n3528 9.01719
R7270 VSS.n3643 VSS.n3642 9.01719
R7271 VSS.n3757 VSS.n3756 9.01719
R7272 VSS.n3871 VSS.n3870 9.01719
R7273 VSS.n2099 VSS.n2098 9.01662
R7274 VSS.n125 VSS.n124 9.01662
R7275 VSS.n1419 VSS.n1418 9.01662
R7276 VSS.n1434 VSS.n1433 9.01662
R7277 VSS.n1449 VSS.n1448 9.01662
R7278 VSS.n1464 VSS.n1463 9.01662
R7279 VSS.n1479 VSS.n1478 9.01662
R7280 VSS.n1997 VSS.n1996 9.01634
R7281 VSS.n2085 VSS.n2084 9.01634
R7282 VSS.n2112 VSS.n2111 9.01634
R7283 VSS.n3401 VSS.n3400 9.01634
R7284 VSS.n3425 VSS.n3424 9.01634
R7285 VSS.n130 VSS.n129 9.01634
R7286 VSS.n1414 VSS.n1413 9.01634
R7287 VSS.n1881 VSS.n1880 9.01634
R7288 VSS.n1429 VSS.n1428 9.01634
R7289 VSS.n1780 VSS.n1779 9.01634
R7290 VSS.n1444 VSS.n1443 9.01634
R7291 VSS.n1679 VSS.n1678 9.01634
R7292 VSS.n1459 VSS.n1458 9.01634
R7293 VSS.n1578 VSS.n1577 9.01634
R7294 VSS.n1474 VSS.n1473 9.01634
R7295 VSS.n1982 VSS.n1981 9.01634
R7296 VSS.n2007 VSS.n2006 9.0162
R7297 VSS.n2122 VSS.n2121 9.0162
R7298 VSS.n1410 VSS.n1409 9.0162
R7299 VSS.n1425 VSS.n1424 9.0162
R7300 VSS.n1440 VSS.n1439 9.0162
R7301 VSS.n1455 VSS.n1454 9.0162
R7302 VSS.n1470 VSS.n1469 9.0162
R7303 VSS.n3894 VSS.n3893 9.01392
R7304 VSS.n3927 VSS.n3926 9.01392
R7305 VSS.n53 VSS.n52 9.01392
R7306 VSS.n3915 VSS.n3914 9.01392
R7307 VSS.n3911 VSS.n3910 9.01392
R7308 VSS.n3905 VSS.n3904 9.01392
R7309 VSS.n3901 VSS.n3900 9.01392
R7310 VSS.n1986 VSS.n1985 9.01392
R7311 VSS.n1985 VSS.n1984 9.01392
R7312 VSS.n1976 VSS.n1975 9.01392
R7313 VSS.n1971 VSS.n1970 9.01392
R7314 VSS.n1967 VSS.n1966 9.01392
R7315 VSS.n1963 VSS.n1962 9.01392
R7316 VSS.n1959 VSS.n1958 9.01392
R7317 VSS.n1953 VSS.n1952 9.01392
R7318 VSS.n1949 VSS.n1948 9.01392
R7319 VSS.n1945 VSS.n1944 9.01392
R7320 VSS.n1941 VSS.n1940 9.01392
R7321 VSS.n1936 VSS.n1935 9.01392
R7322 VSS.n1932 VSS.n1931 9.01392
R7323 VSS.n1928 VSS.n1927 9.01392
R7324 VSS.n1924 VSS.n1923 9.01392
R7325 VSS.n1920 VSS.n1919 9.01392
R7326 VSS.n1914 VSS.n1913 9.01392
R7327 VSS.n1910 VSS.n1909 9.01392
R7328 VSS.n1906 VSS.n1905 9.01392
R7329 VSS.n1902 VSS.n1901 9.01392
R7330 VSS.n1897 VSS.n1896 9.01392
R7331 VSS.n1893 VSS.n1892 9.01392
R7332 VSS.n1888 VSS.n1887 9.01392
R7333 VSS.n1885 VSS.n1884 9.01392
R7334 VSS.n1875 VSS.n1874 9.01392
R7335 VSS.n1870 VSS.n1869 9.01392
R7336 VSS.n1866 VSS.n1865 9.01392
R7337 VSS.n1862 VSS.n1861 9.01392
R7338 VSS.n1858 VSS.n1857 9.01392
R7339 VSS.n1852 VSS.n1851 9.01392
R7340 VSS.n1848 VSS.n1847 9.01392
R7341 VSS.n1844 VSS.n1843 9.01392
R7342 VSS.n1840 VSS.n1839 9.01392
R7343 VSS.n1835 VSS.n1834 9.01392
R7344 VSS.n1831 VSS.n1830 9.01392
R7345 VSS.n1827 VSS.n1826 9.01392
R7346 VSS.n1823 VSS.n1822 9.01392
R7347 VSS.n1819 VSS.n1818 9.01392
R7348 VSS.n1813 VSS.n1812 9.01392
R7349 VSS.n1809 VSS.n1808 9.01392
R7350 VSS.n1805 VSS.n1804 9.01392
R7351 VSS.n1801 VSS.n1800 9.01392
R7352 VSS.n1796 VSS.n1795 9.01392
R7353 VSS.n1792 VSS.n1791 9.01392
R7354 VSS.n1787 VSS.n1786 9.01392
R7355 VSS.n1784 VSS.n1783 9.01392
R7356 VSS.n1774 VSS.n1773 9.01392
R7357 VSS.n1769 VSS.n1768 9.01392
R7358 VSS.n1765 VSS.n1764 9.01392
R7359 VSS.n1761 VSS.n1760 9.01392
R7360 VSS.n1757 VSS.n1756 9.01392
R7361 VSS.n1751 VSS.n1750 9.01392
R7362 VSS.n1747 VSS.n1746 9.01392
R7363 VSS.n1743 VSS.n1742 9.01392
R7364 VSS.n1739 VSS.n1738 9.01392
R7365 VSS.n1734 VSS.n1733 9.01392
R7366 VSS.n1730 VSS.n1729 9.01392
R7367 VSS.n1726 VSS.n1725 9.01392
R7368 VSS.n1722 VSS.n1721 9.01392
R7369 VSS.n1718 VSS.n1717 9.01392
R7370 VSS.n1712 VSS.n1711 9.01392
R7371 VSS.n1708 VSS.n1707 9.01392
R7372 VSS.n1704 VSS.n1703 9.01392
R7373 VSS.n1700 VSS.n1699 9.01392
R7374 VSS.n1695 VSS.n1694 9.01392
R7375 VSS.n1691 VSS.n1690 9.01392
R7376 VSS.n1686 VSS.n1685 9.01392
R7377 VSS.n1683 VSS.n1682 9.01392
R7378 VSS.n1673 VSS.n1672 9.01392
R7379 VSS.n1668 VSS.n1667 9.01392
R7380 VSS.n1664 VSS.n1663 9.01392
R7381 VSS.n1660 VSS.n1659 9.01392
R7382 VSS.n1656 VSS.n1655 9.01392
R7383 VSS.n1650 VSS.n1649 9.01392
R7384 VSS.n1646 VSS.n1645 9.01392
R7385 VSS.n1642 VSS.n1641 9.01392
R7386 VSS.n1638 VSS.n1637 9.01392
R7387 VSS.n1633 VSS.n1632 9.01392
R7388 VSS.n1629 VSS.n1628 9.01392
R7389 VSS.n1625 VSS.n1624 9.01392
R7390 VSS.n1621 VSS.n1620 9.01392
R7391 VSS.n1617 VSS.n1616 9.01392
R7392 VSS.n1611 VSS.n1610 9.01392
R7393 VSS.n1607 VSS.n1606 9.01392
R7394 VSS.n1603 VSS.n1602 9.01392
R7395 VSS.n1599 VSS.n1598 9.01392
R7396 VSS.n1594 VSS.n1593 9.01392
R7397 VSS.n1590 VSS.n1589 9.01392
R7398 VSS.n1585 VSS.n1584 9.01392
R7399 VSS.n1582 VSS.n1581 9.01392
R7400 VSS.n1572 VSS.n1571 9.01392
R7401 VSS.n1567 VSS.n1566 9.01392
R7402 VSS.n1563 VSS.n1562 9.01392
R7403 VSS.n1559 VSS.n1558 9.01392
R7404 VSS.n1555 VSS.n1554 9.01392
R7405 VSS.n1549 VSS.n1548 9.01392
R7406 VSS.n1545 VSS.n1544 9.01392
R7407 VSS.n1541 VSS.n1540 9.01392
R7408 VSS.n1537 VSS.n1536 9.01392
R7409 VSS.n1532 VSS.n1531 9.01392
R7410 VSS.n1528 VSS.n1527 9.01392
R7411 VSS.n1524 VSS.n1523 9.01392
R7412 VSS.n1520 VSS.n1519 9.01392
R7413 VSS.n1516 VSS.n1515 9.01392
R7414 VSS.n1510 VSS.n1509 9.01392
R7415 VSS.n1506 VSS.n1505 9.01392
R7416 VSS.n1502 VSS.n1501 9.01392
R7417 VSS.n1498 VSS.n1497 9.01392
R7418 VSS.n1493 VSS.n1492 9.01392
R7419 VSS.n1489 VSS.n1488 9.01392
R7420 VSS.n59 VSS.n58 9.01392
R7421 VSS.n3407 VSS.n3406 9.01392
R7422 VSS.n3413 VSS.n3412 9.01392
R7423 VSS.n3417 VSS.n3416 9.01392
R7424 VSS.n3421 VSS.n3420 9.01392
R7425 VSS.n3396 VSS.n3395 9.01392
R7426 VSS.n1406 VSS.n1405 9.01392
R7427 VSS.n1405 VSS.n1404 9.01392
R7428 VSS.n79 VSS.n78 9.01392
R7429 VSS.n287 VSS.n286 9.01392
R7430 VSS.n1369 VSS.n1368 9.01392
R7431 VSS.n1379 VSS.n1378 9.01392
R7432 VSS.n1383 VSS.n1382 9.01392
R7433 VSS.n1391 VSS.n1390 9.01392
R7434 VSS.n1400 VSS.n1399 9.01392
R7435 VSS.n2003 VSS.n2002 9.01392
R7436 VSS.n2012 VSS.n2011 9.01392
R7437 VSS.n2016 VSS.n2015 9.01392
R7438 VSS.n2020 VSS.n2019 9.01392
R7439 VSS.n2026 VSS.n2025 9.01392
R7440 VSS.n2030 VSS.n2029 9.01392
R7441 VSS.n2034 VSS.n2033 9.01392
R7442 VSS.n2038 VSS.n2037 9.01392
R7443 VSS.n2043 VSS.n2042 9.01392
R7444 VSS.n2047 VSS.n2046 9.01392
R7445 VSS.n2051 VSS.n2050 9.01392
R7446 VSS.n2055 VSS.n2054 9.01392
R7447 VSS.n2059 VSS.n2058 9.01392
R7448 VSS.n2065 VSS.n2064 9.01392
R7449 VSS.n2069 VSS.n2068 9.01392
R7450 VSS.n2073 VSS.n2072 9.01392
R7451 VSS.n2077 VSS.n2076 9.01392
R7452 VSS.n2081 VSS.n2080 9.01392
R7453 VSS.n2091 VSS.n2090 9.01392
R7454 VSS.n2095 VSS.n2094 9.01392
R7455 VSS.n2106 VSS.n2105 9.01392
R7456 VSS.n2108 VSS.n2107 9.01392
R7457 VSS.n2118 VSS.n2117 9.01392
R7458 VSS.n2127 VSS.n2126 9.01392
R7459 VSS.n2131 VSS.n2130 9.01392
R7460 VSS.n2135 VSS.n2134 9.01392
R7461 VSS.n2141 VSS.n2140 9.01392
R7462 VSS.n2145 VSS.n2144 9.01392
R7463 VSS.n2149 VSS.n2148 9.01392
R7464 VSS.n2153 VSS.n2152 9.01392
R7465 VSS.n2158 VSS.n2157 9.01392
R7466 VSS.n2162 VSS.n2161 9.01392
R7467 VSS.n3886 VSS.n3885 9.01392
R7468 VSS.n3887 VSS.n3886 9.01392
R7469 VSS.n4175 VSS.n4174 9.01392
R7470 VSS.n4172 VSS.n4171 9.01392
R7471 VSS.n3902 VSS.n3901 9.01392
R7472 VSS.n3904 VSS.n3903 9.01392
R7473 VSS.n3910 VSS.n3909 9.01392
R7474 VSS.n3914 VSS.n3913 9.01392
R7475 VSS.n3918 VSS.n3917 9.01392
R7476 VSS.n52 VSS.n51 9.01392
R7477 VSS.n3926 VSS.n3925 9.01392
R7478 VSS.n3891 VSS.n3890 9.01392
R7479 VSS.n3890 VSS.n3889 9.01392
R7480 VSS.n1983 VSS.n1982 9.01392
R7481 VSS.n1975 VSS.n1974 9.01392
R7482 VSS.n1409 VSS.n1408 9.01392
R7483 VSS.n1970 VSS.n1969 9.01392
R7484 VSS.n1966 VSS.n1965 9.01392
R7485 VSS.n1962 VSS.n1961 9.01392
R7486 VSS.n1958 VSS.n1957 9.01392
R7487 VSS.n1952 VSS.n1951 9.01392
R7488 VSS.n1948 VSS.n1947 9.01392
R7489 VSS.n1944 VSS.n1943 9.01392
R7490 VSS.n1940 VSS.n1939 9.01392
R7491 VSS.n1935 VSS.n1934 9.01392
R7492 VSS.n1931 VSS.n1930 9.01392
R7493 VSS.n1927 VSS.n1926 9.01392
R7494 VSS.n1923 VSS.n1922 9.01392
R7495 VSS.n1919 VSS.n1918 9.01392
R7496 VSS.n1913 VSS.n1912 9.01392
R7497 VSS.n1909 VSS.n1908 9.01392
R7498 VSS.n1905 VSS.n1904 9.01392
R7499 VSS.n1901 VSS.n1900 9.01392
R7500 VSS.n1413 VSS.n1412 9.01392
R7501 VSS.n1896 VSS.n1895 9.01392
R7502 VSS.n1892 VSS.n1891 9.01392
R7503 VSS.n1418 VSS.n1417 9.01392
R7504 VSS.n1887 VSS.n1886 9.01392
R7505 VSS.n1884 VSS.n1883 9.01392
R7506 VSS.n1882 VSS.n1881 9.01392
R7507 VSS.n1874 VSS.n1873 9.01392
R7508 VSS.n1424 VSS.n1423 9.01392
R7509 VSS.n1869 VSS.n1868 9.01392
R7510 VSS.n1865 VSS.n1864 9.01392
R7511 VSS.n1861 VSS.n1860 9.01392
R7512 VSS.n1857 VSS.n1856 9.01392
R7513 VSS.n1851 VSS.n1850 9.01392
R7514 VSS.n1847 VSS.n1846 9.01392
R7515 VSS.n1843 VSS.n1842 9.01392
R7516 VSS.n1839 VSS.n1838 9.01392
R7517 VSS.n1834 VSS.n1833 9.01392
R7518 VSS.n1830 VSS.n1829 9.01392
R7519 VSS.n1826 VSS.n1825 9.01392
R7520 VSS.n1822 VSS.n1821 9.01392
R7521 VSS.n1818 VSS.n1817 9.01392
R7522 VSS.n1812 VSS.n1811 9.01392
R7523 VSS.n1808 VSS.n1807 9.01392
R7524 VSS.n1804 VSS.n1803 9.01392
R7525 VSS.n1800 VSS.n1799 9.01392
R7526 VSS.n1428 VSS.n1427 9.01392
R7527 VSS.n1795 VSS.n1794 9.01392
R7528 VSS.n1791 VSS.n1790 9.01392
R7529 VSS.n1433 VSS.n1432 9.01392
R7530 VSS.n1786 VSS.n1785 9.01392
R7531 VSS.n1783 VSS.n1782 9.01392
R7532 VSS.n1781 VSS.n1780 9.01392
R7533 VSS.n1773 VSS.n1772 9.01392
R7534 VSS.n1439 VSS.n1438 9.01392
R7535 VSS.n1768 VSS.n1767 9.01392
R7536 VSS.n1764 VSS.n1763 9.01392
R7537 VSS.n1760 VSS.n1759 9.01392
R7538 VSS.n1756 VSS.n1755 9.01392
R7539 VSS.n1750 VSS.n1749 9.01392
R7540 VSS.n1746 VSS.n1745 9.01392
R7541 VSS.n1742 VSS.n1741 9.01392
R7542 VSS.n1738 VSS.n1737 9.01392
R7543 VSS.n1733 VSS.n1732 9.01392
R7544 VSS.n1729 VSS.n1728 9.01392
R7545 VSS.n1725 VSS.n1724 9.01392
R7546 VSS.n1721 VSS.n1720 9.01392
R7547 VSS.n1717 VSS.n1716 9.01392
R7548 VSS.n1711 VSS.n1710 9.01392
R7549 VSS.n1707 VSS.n1706 9.01392
R7550 VSS.n1703 VSS.n1702 9.01392
R7551 VSS.n1699 VSS.n1698 9.01392
R7552 VSS.n1443 VSS.n1442 9.01392
R7553 VSS.n1694 VSS.n1693 9.01392
R7554 VSS.n1690 VSS.n1689 9.01392
R7555 VSS.n1448 VSS.n1447 9.01392
R7556 VSS.n1685 VSS.n1684 9.01392
R7557 VSS.n1682 VSS.n1681 9.01392
R7558 VSS.n1680 VSS.n1679 9.01392
R7559 VSS.n1672 VSS.n1671 9.01392
R7560 VSS.n1454 VSS.n1453 9.01392
R7561 VSS.n1667 VSS.n1666 9.01392
R7562 VSS.n1663 VSS.n1662 9.01392
R7563 VSS.n1659 VSS.n1658 9.01392
R7564 VSS.n1655 VSS.n1654 9.01392
R7565 VSS.n1649 VSS.n1648 9.01392
R7566 VSS.n1645 VSS.n1644 9.01392
R7567 VSS.n1641 VSS.n1640 9.01392
R7568 VSS.n1637 VSS.n1636 9.01392
R7569 VSS.n1632 VSS.n1631 9.01392
R7570 VSS.n1628 VSS.n1627 9.01392
R7571 VSS.n1624 VSS.n1623 9.01392
R7572 VSS.n1620 VSS.n1619 9.01392
R7573 VSS.n1616 VSS.n1615 9.01392
R7574 VSS.n1610 VSS.n1609 9.01392
R7575 VSS.n1606 VSS.n1605 9.01392
R7576 VSS.n1602 VSS.n1601 9.01392
R7577 VSS.n1598 VSS.n1597 9.01392
R7578 VSS.n1458 VSS.n1457 9.01392
R7579 VSS.n1593 VSS.n1592 9.01392
R7580 VSS.n1589 VSS.n1588 9.01392
R7581 VSS.n1463 VSS.n1462 9.01392
R7582 VSS.n1584 VSS.n1583 9.01392
R7583 VSS.n1581 VSS.n1580 9.01392
R7584 VSS.n1579 VSS.n1578 9.01392
R7585 VSS.n1571 VSS.n1570 9.01392
R7586 VSS.n1469 VSS.n1468 9.01392
R7587 VSS.n1566 VSS.n1565 9.01392
R7588 VSS.n1562 VSS.n1561 9.01392
R7589 VSS.n1558 VSS.n1557 9.01392
R7590 VSS.n1554 VSS.n1553 9.01392
R7591 VSS.n1548 VSS.n1547 9.01392
R7592 VSS.n1544 VSS.n1543 9.01392
R7593 VSS.n1540 VSS.n1539 9.01392
R7594 VSS.n1536 VSS.n1535 9.01392
R7595 VSS.n1531 VSS.n1530 9.01392
R7596 VSS.n1527 VSS.n1526 9.01392
R7597 VSS.n1523 VSS.n1522 9.01392
R7598 VSS.n1519 VSS.n1518 9.01392
R7599 VSS.n1515 VSS.n1514 9.01392
R7600 VSS.n1509 VSS.n1508 9.01392
R7601 VSS.n1505 VSS.n1504 9.01392
R7602 VSS.n1501 VSS.n1500 9.01392
R7603 VSS.n1497 VSS.n1496 9.01392
R7604 VSS.n1473 VSS.n1472 9.01392
R7605 VSS.n1492 VSS.n1491 9.01392
R7606 VSS.n1488 VSS.n1487 9.01392
R7607 VSS.n1478 VSS.n1477 9.01392
R7608 VSS.n1484 VSS.n1483 9.01392
R7609 VSS.n1483 VSS.n1482 9.01392
R7610 VSS.n3395 VSS.n3394 9.01392
R7611 VSS.n58 VSS.n57 9.01392
R7612 VSS.n3400 VSS.n3399 9.01392
R7613 VSS.n3406 VSS.n3405 9.01392
R7614 VSS.n3412 VSS.n3411 9.01392
R7615 VSS.n3418 VSS.n3417 9.01392
R7616 VSS.n3420 VSS.n3419 9.01392
R7617 VSS.n3424 VSS.n3423 9.01392
R7618 VSS.n3431 VSS.n3430 9.01392
R7619 VSS.n3432 VSS.n3431 9.01392
R7620 VSS.n124 VSS.n123 9.01392
R7621 VSS.n1399 VSS.n1398 9.01392
R7622 VSS.n129 VSS.n128 9.01392
R7623 VSS.n1390 VSS.n1389 9.01392
R7624 VSS.n1382 VSS.n1381 9.01392
R7625 VSS.n1378 VSS.n1377 9.01392
R7626 VSS.n1368 VSS.n1367 9.01392
R7627 VSS.n286 VSS.n285 9.01392
R7628 VSS.n78 VSS.n77 9.01392
R7629 VSS.n3336 VSS.n3335 9.01392
R7630 VSS.n3335 VSS.n3334 9.01392
R7631 VSS.n1375 VSS.n1374 9.01392
R7632 VSS.n1374 VSS.n1373 9.01392
R7633 VSS.n1387 VSS.n1386 9.01392
R7634 VSS.n1386 VSS.n1385 9.01392
R7635 VSS.n1396 VSS.n1395 9.01392
R7636 VSS.n1395 VSS.n1394 9.01392
R7637 VSS.n1996 VSS.n1995 9.01392
R7638 VSS.n2002 VSS.n2001 9.01392
R7639 VSS.n2006 VSS.n2005 9.01392
R7640 VSS.n2011 VSS.n2010 9.01392
R7641 VSS.n2015 VSS.n2014 9.01392
R7642 VSS.n2019 VSS.n2018 9.01392
R7643 VSS.n2025 VSS.n2024 9.01392
R7644 VSS.n2029 VSS.n2028 9.01392
R7645 VSS.n2033 VSS.n2032 9.01392
R7646 VSS.n2037 VSS.n2036 9.01392
R7647 VSS.n2042 VSS.n2041 9.01392
R7648 VSS.n2046 VSS.n2045 9.01392
R7649 VSS.n2050 VSS.n2049 9.01392
R7650 VSS.n2054 VSS.n2053 9.01392
R7651 VSS.n2058 VSS.n2057 9.01392
R7652 VSS.n2064 VSS.n2063 9.01392
R7653 VSS.n2068 VSS.n2067 9.01392
R7654 VSS.n2072 VSS.n2071 9.01392
R7655 VSS.n2076 VSS.n2075 9.01392
R7656 VSS.n2080 VSS.n2079 9.01392
R7657 VSS.n2084 VSS.n2083 9.01392
R7658 VSS.n2090 VSS.n2089 9.01392
R7659 VSS.n2094 VSS.n2093 9.01392
R7660 VSS.n2098 VSS.n2097 9.01392
R7661 VSS.n2105 VSS.n2104 9.01392
R7662 VSS.n2109 VSS.n2108 9.01392
R7663 VSS.n2111 VSS.n2110 9.01392
R7664 VSS.n2117 VSS.n2116 9.01392
R7665 VSS.n2121 VSS.n2120 9.01392
R7666 VSS.n2126 VSS.n2125 9.01392
R7667 VSS.n2130 VSS.n2129 9.01392
R7668 VSS.n2134 VSS.n2133 9.01392
R7669 VSS.n2140 VSS.n2139 9.01392
R7670 VSS.n2144 VSS.n2143 9.01392
R7671 VSS.n2148 VSS.n2147 9.01392
R7672 VSS.n2152 VSS.n2151 9.01392
R7673 VSS.n2157 VSS.n2156 9.01392
R7674 VSS.n2161 VSS.n2160 9.01392
R7675 VSS.n1993 VSS.n1992 9.01392
R7676 VSS.n1994 VSS.n1993 9.01392
R7677 VSS.n3879 VSS.n3878 9.01392
R7678 VSS.n3876 VSS.n3875 9.01392
R7679 VSS.n3875 VSS.n3874 9.01392
R7680 VSS.n3870 VSS.n3869 9.01392
R7681 VSS.n3867 VSS.n3866 9.01392
R7682 VSS.n3866 VSS.n3865 9.01392
R7683 VSS.n3863 VSS.n3862 9.01392
R7684 VSS.n3862 VSS.n3861 9.01392
R7685 VSS.n3859 VSS.n3858 9.01392
R7686 VSS.n3858 VSS.n3857 9.01392
R7687 VSS.n3855 VSS.n3854 9.01392
R7688 VSS.n3854 VSS.n3853 9.01392
R7689 VSS.n3849 VSS.n3848 9.01392
R7690 VSS.n3848 VSS.n3847 9.01392
R7691 VSS.n3845 VSS.n3844 9.01392
R7692 VSS.n3844 VSS.n3843 9.01392
R7693 VSS.n3841 VSS.n3840 9.01392
R7694 VSS.n3840 VSS.n3839 9.01392
R7695 VSS.n3837 VSS.n3836 9.01392
R7696 VSS.n3836 VSS.n3835 9.01392
R7697 VSS.n3832 VSS.n3831 9.01392
R7698 VSS.n3831 VSS.n3830 9.01392
R7699 VSS.n3828 VSS.n3827 9.01392
R7700 VSS.n3827 VSS.n3826 9.01392
R7701 VSS.n3824 VSS.n3823 9.01392
R7702 VSS.n3823 VSS.n3822 9.01392
R7703 VSS.n3820 VSS.n3819 9.01392
R7704 VSS.n3819 VSS.n3818 9.01392
R7705 VSS.n3816 VSS.n3815 9.01392
R7706 VSS.n3815 VSS.n3814 9.01392
R7707 VSS.n3810 VSS.n3809 9.01392
R7708 VSS.n3809 VSS.n3808 9.01392
R7709 VSS.n3806 VSS.n3805 9.01392
R7710 VSS.n3805 VSS.n3804 9.01392
R7711 VSS.n3802 VSS.n3801 9.01392
R7712 VSS.n3801 VSS.n3800 9.01392
R7713 VSS.n3798 VSS.n3797 9.01392
R7714 VSS.n3797 VSS.n3796 9.01392
R7715 VSS.n3791 VSS.n3790 9.01392
R7716 VSS.n3788 VSS.n3787 9.01392
R7717 VSS.n3787 VSS.n3786 9.01392
R7718 VSS.n3784 VSS.n3783 9.01392
R7719 VSS.n3783 VSS.n3782 9.01392
R7720 VSS.n3777 VSS.n3776 9.01392
R7721 VSS.n3774 VSS.n3773 9.01392
R7722 VSS.n3773 VSS.n3772 9.01392
R7723 VSS.n3764 VSS.n3434 9.01392
R7724 VSS.n3771 VSS.n3434 9.01392
R7725 VSS.n3770 VSS.n3769 9.01392
R7726 VSS.n3762 VSS.n3761 9.01392
R7727 VSS.n3761 VSS.n3760 9.01392
R7728 VSS.n3756 VSS.n3755 9.01392
R7729 VSS.n3753 VSS.n3752 9.01392
R7730 VSS.n3752 VSS.n3751 9.01392
R7731 VSS.n3749 VSS.n3748 9.01392
R7732 VSS.n3748 VSS.n3747 9.01392
R7733 VSS.n3745 VSS.n3744 9.01392
R7734 VSS.n3744 VSS.n3743 9.01392
R7735 VSS.n3741 VSS.n3740 9.01392
R7736 VSS.n3740 VSS.n3739 9.01392
R7737 VSS.n3735 VSS.n3734 9.01392
R7738 VSS.n3734 VSS.n3733 9.01392
R7739 VSS.n3731 VSS.n3730 9.01392
R7740 VSS.n3730 VSS.n3729 9.01392
R7741 VSS.n3727 VSS.n3726 9.01392
R7742 VSS.n3726 VSS.n3725 9.01392
R7743 VSS.n3723 VSS.n3722 9.01392
R7744 VSS.n3722 VSS.n3721 9.01392
R7745 VSS.n3718 VSS.n3717 9.01392
R7746 VSS.n3717 VSS.n3716 9.01392
R7747 VSS.n3714 VSS.n3713 9.01392
R7748 VSS.n3713 VSS.n3712 9.01392
R7749 VSS.n3710 VSS.n3709 9.01392
R7750 VSS.n3709 VSS.n3708 9.01392
R7751 VSS.n3706 VSS.n3705 9.01392
R7752 VSS.n3705 VSS.n3704 9.01392
R7753 VSS.n3702 VSS.n3701 9.01392
R7754 VSS.n3701 VSS.n3700 9.01392
R7755 VSS.n3696 VSS.n3695 9.01392
R7756 VSS.n3695 VSS.n3694 9.01392
R7757 VSS.n3692 VSS.n3691 9.01392
R7758 VSS.n3691 VSS.n3690 9.01392
R7759 VSS.n3688 VSS.n3687 9.01392
R7760 VSS.n3687 VSS.n3686 9.01392
R7761 VSS.n3684 VSS.n3683 9.01392
R7762 VSS.n3683 VSS.n3682 9.01392
R7763 VSS.n3677 VSS.n3676 9.01392
R7764 VSS.n3674 VSS.n3673 9.01392
R7765 VSS.n3673 VSS.n3672 9.01392
R7766 VSS.n3670 VSS.n3669 9.01392
R7767 VSS.n3669 VSS.n3668 9.01392
R7768 VSS.n3663 VSS.n3662 9.01392
R7769 VSS.n3660 VSS.n3659 9.01392
R7770 VSS.n3659 VSS.n3658 9.01392
R7771 VSS.n3650 VSS.n3436 9.01392
R7772 VSS.n3657 VSS.n3436 9.01392
R7773 VSS.n3656 VSS.n3655 9.01392
R7774 VSS.n3648 VSS.n3647 9.01392
R7775 VSS.n3647 VSS.n3646 9.01392
R7776 VSS.n3642 VSS.n3641 9.01392
R7777 VSS.n3639 VSS.n3638 9.01392
R7778 VSS.n3638 VSS.n3637 9.01392
R7779 VSS.n3635 VSS.n3634 9.01392
R7780 VSS.n3634 VSS.n3633 9.01392
R7781 VSS.n3631 VSS.n3630 9.01392
R7782 VSS.n3630 VSS.n3629 9.01392
R7783 VSS.n3627 VSS.n3626 9.01392
R7784 VSS.n3626 VSS.n3625 9.01392
R7785 VSS.n3621 VSS.n3620 9.01392
R7786 VSS.n3620 VSS.n3619 9.01392
R7787 VSS.n3617 VSS.n3616 9.01392
R7788 VSS.n3616 VSS.n3615 9.01392
R7789 VSS.n3613 VSS.n3612 9.01392
R7790 VSS.n3612 VSS.n3611 9.01392
R7791 VSS.n3609 VSS.n3608 9.01392
R7792 VSS.n3608 VSS.n3607 9.01392
R7793 VSS.n3604 VSS.n3603 9.01392
R7794 VSS.n3603 VSS.n3602 9.01392
R7795 VSS.n3600 VSS.n3599 9.01392
R7796 VSS.n3599 VSS.n3598 9.01392
R7797 VSS.n3596 VSS.n3595 9.01392
R7798 VSS.n3595 VSS.n3594 9.01392
R7799 VSS.n3592 VSS.n3591 9.01392
R7800 VSS.n3591 VSS.n3590 9.01392
R7801 VSS.n3588 VSS.n3587 9.01392
R7802 VSS.n3587 VSS.n3586 9.01392
R7803 VSS.n3582 VSS.n3581 9.01392
R7804 VSS.n3581 VSS.n3580 9.01392
R7805 VSS.n3578 VSS.n3577 9.01392
R7806 VSS.n3577 VSS.n3576 9.01392
R7807 VSS.n3574 VSS.n3573 9.01392
R7808 VSS.n3573 VSS.n3572 9.01392
R7809 VSS.n3570 VSS.n3569 9.01392
R7810 VSS.n3569 VSS.n3568 9.01392
R7811 VSS.n3563 VSS.n3562 9.01392
R7812 VSS.n3560 VSS.n3559 9.01392
R7813 VSS.n3559 VSS.n3558 9.01392
R7814 VSS.n3556 VSS.n3555 9.01392
R7815 VSS.n3555 VSS.n3554 9.01392
R7816 VSS.n3549 VSS.n3548 9.01392
R7817 VSS.n3546 VSS.n3545 9.01392
R7818 VSS.n3545 VSS.n3544 9.01392
R7819 VSS.n3536 VSS.n3438 9.01392
R7820 VSS.n3543 VSS.n3438 9.01392
R7821 VSS.n3542 VSS.n3541 9.01392
R7822 VSS.n3534 VSS.n3533 9.01392
R7823 VSS.n3533 VSS.n3532 9.01392
R7824 VSS.n3528 VSS.n3527 9.01392
R7825 VSS.n3525 VSS.n3524 9.01392
R7826 VSS.n3524 VSS.n3523 9.01392
R7827 VSS.n3521 VSS.n3520 9.01392
R7828 VSS.n3520 VSS.n3519 9.01392
R7829 VSS.n3517 VSS.n3516 9.01392
R7830 VSS.n3516 VSS.n3515 9.01392
R7831 VSS.n3513 VSS.n3512 9.01392
R7832 VSS.n3512 VSS.n3511 9.01392
R7833 VSS.n3507 VSS.n3506 9.01392
R7834 VSS.n3506 VSS.n3505 9.01392
R7835 VSS.n3503 VSS.n3502 9.01392
R7836 VSS.n3502 VSS.n3501 9.01392
R7837 VSS.n3499 VSS.n3498 9.01392
R7838 VSS.n3498 VSS.n3497 9.01392
R7839 VSS.n3495 VSS.n3494 9.01392
R7840 VSS.n3494 VSS.n3493 9.01392
R7841 VSS.n3490 VSS.n3489 9.01392
R7842 VSS.n3489 VSS.n3488 9.01392
R7843 VSS.n3486 VSS.n3485 9.01392
R7844 VSS.n3485 VSS.n3484 9.01392
R7845 VSS.n3482 VSS.n3481 9.01392
R7846 VSS.n3481 VSS.n3480 9.01392
R7847 VSS.n3478 VSS.n3477 9.01392
R7848 VSS.n3477 VSS.n3476 9.01392
R7849 VSS.n3474 VSS.n3473 9.01392
R7850 VSS.n3473 VSS.n3472 9.01392
R7851 VSS.n3468 VSS.n3467 9.01392
R7852 VSS.n3467 VSS.n3466 9.01392
R7853 VSS.n3464 VSS.n3463 9.01392
R7854 VSS.n3463 VSS.n3462 9.01392
R7855 VSS.n3460 VSS.n3459 9.01392
R7856 VSS.n3459 VSS.n3458 9.01392
R7857 VSS.n3456 VSS.n3455 9.01392
R7858 VSS.n3455 VSS.n3454 9.01392
R7859 VSS.n3449 VSS.n3448 9.01392
R7860 VSS.n3446 VSS.n3445 9.01392
R7861 VSS.n3445 VSS.n3444 9.01392
R7862 VSS.n3442 VSS.n3441 9.01392
R7863 VSS.n3441 VSS.n3440 9.01392
R7864 VSS.n2 VSS.n1 9.01392
R7865 VSS.n4286 VSS.n4285 9.01392
R7866 VSS.n4285 VSS.n4284 9.01392
R7867 VSS.n4282 VSS.n4281 9.01392
R7868 VSS.n4283 VSS.n4282 9.01392
R7869 VSS.n4280 VSS.n4279 9.01392
R7870 VSS.n4274 VSS.n4273 9.01392
R7871 VSS.n4273 VSS.n4272 9.01392
R7872 VSS.n4268 VSS.n4267 9.01392
R7873 VSS.n4265 VSS.n4264 9.01392
R7874 VSS.n4264 VSS.n4263 9.01392
R7875 VSS.n4261 VSS.n4260 9.01392
R7876 VSS.n4260 VSS.n4259 9.01392
R7877 VSS.n4257 VSS.n4256 9.01392
R7878 VSS.n4256 VSS.n4255 9.01392
R7879 VSS.n4253 VSS.n4252 9.01392
R7880 VSS.n4252 VSS.n4251 9.01392
R7881 VSS.n4247 VSS.n4246 9.01392
R7882 VSS.n4246 VSS.n4245 9.01392
R7883 VSS.n4243 VSS.n4242 9.01392
R7884 VSS.n4242 VSS.n4241 9.01392
R7885 VSS.n4239 VSS.n4238 9.01392
R7886 VSS.n4238 VSS.n4237 9.01392
R7887 VSS.n4235 VSS.n4234 9.01392
R7888 VSS.n4234 VSS.n4233 9.01392
R7889 VSS.n4230 VSS.n4229 9.01392
R7890 VSS.n4229 VSS.n4228 9.01392
R7891 VSS.n4226 VSS.n4225 9.01392
R7892 VSS.n4225 VSS.n4224 9.01392
R7893 VSS.n4222 VSS.n4221 9.01392
R7894 VSS.n4221 VSS.n4220 9.01392
R7895 VSS.n4218 VSS.n4217 9.01392
R7896 VSS.n4217 VSS.n4216 9.01392
R7897 VSS.n4214 VSS.n4213 9.01392
R7898 VSS.n4213 VSS.n4212 9.01392
R7899 VSS.n4208 VSS.n4207 9.01392
R7900 VSS.n4207 VSS.n4206 9.01392
R7901 VSS.n4204 VSS.n4203 9.01392
R7902 VSS.n4203 VSS.n4202 9.01392
R7903 VSS.n4200 VSS.n4199 9.01392
R7904 VSS.n4199 VSS.n4198 9.01392
R7905 VSS.n4196 VSS.n4195 9.01392
R7906 VSS.n4195 VSS.n4194 9.01392
R7907 VSS.n4189 VSS.n4188 9.01392
R7908 VSS.n4186 VSS.n4185 9.01392
R7909 VSS.n4185 VSS.n4184 9.01392
R7910 VSS.n4182 VSS.n4181 9.01392
R7911 VSS.n4181 VSS.n4180 9.01392
R7912 VSS.n4171 VSS.n4170 9.01392
R7913 VSS VSS.n1994 8.8005
R7914 VSS.n2032 VSS.t497 8.8005
R7915 VSS VSS.n2109 8.8005
R7916 VSS.n2147 VSS.t40 8.8005
R7917 VSS.n2453 VSS.t157 8.8005
R7918 VSS.n2481 VSS.t119 8.8005
R7919 VSS.n2805 VSS.t147 8.8005
R7920 VSS.n2833 VSS.t219 8.8005
R7921 VSS.n3333 VSS.n82 8.8005
R7922 VSS.n265 VSS.n262 8.76429
R7923 VSS.n272 VSS.n271 8.76429
R7924 VSS.n1997 VSS 8.6074
R7925 VSS.n2065 VSS.n2062 8.6074
R7926 VSS.n2112 VSS 8.6074
R7927 VSS.n2359 VSS 8.6074
R7928 VSS.n2711 VSS 8.6074
R7929 VSS.n3322 VSS.n3321 8.6074
R7930 VSS.n1375 VSS.n1372 8.6074
R7931 VSS.n1920 VSS.n1917 8.6074
R7932 VSS.n1819 VSS.n1816 8.6074
R7933 VSS.n1718 VSS.n1715 8.6074
R7934 VSS.n1617 VSS.n1614 8.6074
R7935 VSS.n1516 VSS.n1513 8.6074
R7936 VSS.n4214 VSS.n4211 8.6074
R7937 VSS.n3474 VSS.n3471 8.6074
R7938 VSS.n3588 VSS.n3585 8.6074
R7939 VSS.n3702 VSS.n3699 8.6074
R7940 VSS.n3816 VSS.n3813 8.6074
R7941 VSS.t283 VSS.n21 8.5775
R7942 VSS.n1313 VSS.t76 8.5775
R7943 VSS.n1220 VSS 8.5775
R7944 VSS.t32 VSS.n1112 8.5775
R7945 VSS.t129 VSS.n794 8.5775
R7946 VSS.t53 VSS.n476 8.5775
R7947 VSS.n3157 VSS.n3156 7.72464
R7948 VSS.n2329 VSS.n2328 7.57647
R7949 VSS.n2681 VSS.n2680 7.57647
R7950 VSS.n3033 VSS.n3032 7.57647
R7951 VSS.n168 VSS.n167 7.57501
R7952 VSS.n194 VSS.n193 7.57501
R7953 VSS.n213 VSS.n212 7.57501
R7954 VSS.n239 VSS.n238 7.57501
R7955 VSS.n258 VSS.n257 7.57501
R7956 VSS.n158 VSS.n157 7.57431
R7957 VSS.n203 VSS.n202 7.57431
R7958 VSS.n248 VSS.n247 7.57431
R7959 VSS.n2442 VSS.n2441 7.50395
R7960 VSS.n2794 VSS.n2793 7.50395
R7961 VSS.n1251 VSS.n1246 7.45502
R7962 VSS.n1230 VSS.n1225 7.43981
R7963 VSS.n1186 VSS.n1181 7.43981
R7964 VSS.n496 VSS.n495 6.84188
R7965 VSS.n814 VSS.n813 6.84188
R7966 VSS.n1132 VSS.n1131 6.84188
R7967 VSS.n266 VSS 6.66075
R7968 VSS.n4164 VSS.n4163 6.62119
R7969 VSS.n3287 VSS.t353 6.37269
R7970 VSS.n3138 VSS.t533 6.37269
R7971 VSS.n3375 VSS.n76 6.30775
R7972 VSS.n10 VSS.n9 5.71609
R7973 VSS.n267 VSS 5.58923
R7974 VSS.n60 VSS.n59 5.51774
R7975 VSS.n54 VSS.n53 5.51774
R7976 VSS.n1984 VSS 5.26996
R7977 VSS.n1947 VSS.t175 5.26996
R7978 VSS.n1883 VSS 5.26996
R7979 VSS.n1846 VSS.t688 5.26996
R7980 VSS.n1782 VSS 5.26996
R7981 VSS.n1745 VSS.t287 5.26996
R7982 VSS.n1681 VSS 5.26996
R7983 VSS.n1644 VSS.t459 5.26996
R7984 VSS.n1580 VSS 5.26996
R7985 VSS.n1543 VSS.t305 5.26996
R7986 VSS.n271 VSS.n270 5.25868
R7987 VSS.n3292 VSS.n3291 5.07636
R7988 VSS.n3021 VSS.n3020 4.6505
R7989 VSS.n2176 VSS.n2175 4.6505
R7990 VSS.n2190 VSS.n2189 4.6505
R7991 VSS.n2204 VSS.n2203 4.6505
R7992 VSS.n2220 VSS.n2219 4.6505
R7993 VSS.n2234 VSS.n2233 4.6505
R7994 VSS.n2248 VSS.n2247 4.6505
R7995 VSS.n2262 VSS.n2261 4.6505
R7996 VSS.n2276 VSS.n2275 4.6505
R7997 VSS.n2303 VSS.n2302 4.6505
R7998 VSS.n2317 VSS.n2316 4.6505
R7999 VSS.n2346 VSS.n2345 4.6505
R8000 VSS.n2351 VSS.n2350 4.6505
R8001 VSS.n2375 VSS.n2374 4.6505
R8002 VSS.n2401 VSS.n2400 4.6505
R8003 VSS.n2415 VSS.n2414 4.6505
R8004 VSS.n2429 VSS.n2428 4.6505
R8005 VSS.n2444 VSS.n2443 4.6505
R8006 VSS.n2458 VSS.n2457 4.6505
R8007 VSS.n2472 VSS.n2471 4.6505
R8008 VSS.n2486 VSS.n2485 4.6505
R8009 VSS.n2501 VSS.n2500 4.6505
R8010 VSS.n2514 VSS.n2513 4.6505
R8011 VSS.n2528 VSS.n2527 4.6505
R8012 VSS.n2542 VSS.n2541 4.6505
R8013 VSS.n2556 VSS.n2555 4.6505
R8014 VSS.n2572 VSS.n2571 4.6505
R8015 VSS.n2586 VSS.n2585 4.6505
R8016 VSS.n2600 VSS.n2599 4.6505
R8017 VSS.n2614 VSS.n2613 4.6505
R8018 VSS.n2628 VSS.n2627 4.6505
R8019 VSS.n2655 VSS.n2654 4.6505
R8020 VSS.n2669 VSS.n2668 4.6505
R8021 VSS.n2698 VSS.n2697 4.6505
R8022 VSS.n2703 VSS.n2702 4.6505
R8023 VSS.n2727 VSS.n2726 4.6505
R8024 VSS.n2753 VSS.n2752 4.6505
R8025 VSS.n2767 VSS.n2766 4.6505
R8026 VSS.n2781 VSS.n2780 4.6505
R8027 VSS.n2796 VSS.n2795 4.6505
R8028 VSS.n2810 VSS.n2809 4.6505
R8029 VSS.n2824 VSS.n2823 4.6505
R8030 VSS.n2838 VSS.n2837 4.6505
R8031 VSS.n2853 VSS.n2852 4.6505
R8032 VSS.n2866 VSS.n2865 4.6505
R8033 VSS.n2880 VSS.n2879 4.6505
R8034 VSS.n2894 VSS.n2893 4.6505
R8035 VSS.n2908 VSS.n2907 4.6505
R8036 VSS.n2924 VSS.n2923 4.6505
R8037 VSS.n2938 VSS.n2937 4.6505
R8038 VSS.n2952 VSS.n2951 4.6505
R8039 VSS.n2966 VSS.n2965 4.6505
R8040 VSS.n2980 VSS.n2979 4.6505
R8041 VSS.n3007 VSS.n3006 4.6505
R8042 VSS.n3040 VSS.n3039 4.6505
R8043 VSS.n3054 VSS.n3053 4.6505
R8044 VSS.n3068 VSS.n3067 4.6505
R8045 VSS.n3082 VSS.n3081 4.6505
R8046 VSS.n3328 VSS.n3327 4.6505
R8047 VSS.n3324 VSS.n3323 4.6505
R8048 VSS.n3308 VSS.n3307 4.6505
R8049 VSS.n3294 VSS.n3293 4.6505
R8050 VSS.n3278 VSS.n3277 4.6505
R8051 VSS.n3265 VSS.n3264 4.6505
R8052 VSS.n3249 VSS.n3248 4.6505
R8053 VSS.n3235 VSS.n3234 4.6505
R8054 VSS.n3219 VSS.n3218 4.6505
R8055 VSS.n3205 VSS.n3204 4.6505
R8056 VSS.n3189 VSS.n3188 4.6505
R8057 VSS.n3175 VSS.n3174 4.6505
R8058 VSS.n3159 VSS.n3158 4.6505
R8059 VSS.n3143 VSS.n3142 4.6505
R8060 VSS.n3129 VSS.n3128 4.6505
R8061 VSS.n3113 VSS.n3112 4.6505
R8062 VSS.n3099 VSS.n3098 4.6505
R8063 VSS.n3384 VSS.n3383 4.6505
R8064 VSS.n3389 VSS.n3388 4.6505
R8065 VSS.n4150 VSS.n4149 4.6505
R8066 VSS.n4145 VSS.n4144 4.6505
R8067 VSS.n4131 VSS.n4130 4.6505
R8068 VSS.n4115 VSS.n4114 4.6505
R8069 VSS.n4103 VSS.n4102 4.6505
R8070 VSS.n4089 VSS.n4088 4.6505
R8071 VSS.n4075 VSS.n4074 4.6505
R8072 VSS.n4058 VSS.n4057 4.6505
R8073 VSS.n4046 VSS.n4045 4.6505
R8074 VSS.n4032 VSS.n4031 4.6505
R8075 VSS.n4018 VSS.n4017 4.6505
R8076 VSS.n4004 VSS.n4003 4.6505
R8077 VSS.n3989 VSS.n3988 4.6505
R8078 VSS.n3975 VSS.n3974 4.6505
R8079 VSS.n3960 VSS.n3959 4.6505
R8080 VSS.n3946 VSS.n3945 4.6505
R8081 VSS.n1148 VSS.n1147 4.6505
R8082 VSS.n1134 VSS.n1133 4.6505
R8083 VSS.n1118 VSS.n1117 4.6505
R8084 VSS.n1104 VSS.n1103 4.6505
R8085 VSS.n1090 VSS.n1089 4.6505
R8086 VSS.n1076 VSS.n1075 4.6505
R8087 VSS.n1062 VSS.n1061 4.6505
R8088 VSS.n1048 VSS.n1047 4.6505
R8089 VSS.n1034 VSS.n1033 4.6505
R8090 VSS.n1020 VSS.n1019 4.6505
R8091 VSS.n1006 VSS.n1005 4.6505
R8092 VSS.n990 VSS.n989 4.6505
R8093 VSS.n976 VSS.n975 4.6505
R8094 VSS.n962 VSS.n961 4.6505
R8095 VSS.n945 VSS.n944 4.6505
R8096 VSS.n928 VSS.n927 4.6505
R8097 VSS.n910 VSS.n909 4.6505
R8098 VSS.n903 VSS.n902 4.6505
R8099 VSS.n889 VSS.n888 4.6505
R8100 VSS.n872 VSS.n871 4.6505
R8101 VSS.n858 VSS.n857 4.6505
R8102 VSS.n844 VSS.n843 4.6505
R8103 VSS.n830 VSS.n829 4.6505
R8104 VSS.n816 VSS.n815 4.6505
R8105 VSS.n800 VSS.n799 4.6505
R8106 VSS.n786 VSS.n785 4.6505
R8107 VSS.n772 VSS.n771 4.6505
R8108 VSS.n758 VSS.n757 4.6505
R8109 VSS.n744 VSS.n743 4.6505
R8110 VSS.n730 VSS.n729 4.6505
R8111 VSS.n716 VSS.n715 4.6505
R8112 VSS.n702 VSS.n701 4.6505
R8113 VSS.n688 VSS.n687 4.6505
R8114 VSS.n672 VSS.n671 4.6505
R8115 VSS.n658 VSS.n657 4.6505
R8116 VSS.n644 VSS.n643 4.6505
R8117 VSS.n627 VSS.n626 4.6505
R8118 VSS.n610 VSS.n609 4.6505
R8119 VSS.n592 VSS.n591 4.6505
R8120 VSS.n585 VSS.n584 4.6505
R8121 VSS.n571 VSS.n570 4.6505
R8122 VSS.n554 VSS.n553 4.6505
R8123 VSS.n540 VSS.n539 4.6505
R8124 VSS.n526 VSS.n525 4.6505
R8125 VSS.n512 VSS.n511 4.6505
R8126 VSS.n498 VSS.n497 4.6505
R8127 VSS.n482 VSS.n481 4.6505
R8128 VSS.n468 VSS.n467 4.6505
R8129 VSS.n454 VSS.n453 4.6505
R8130 VSS.n440 VSS.n439 4.6505
R8131 VSS.n426 VSS.n425 4.6505
R8132 VSS.n412 VSS.n411 4.6505
R8133 VSS.n398 VSS.n397 4.6505
R8134 VSS.n384 VSS.n383 4.6505
R8135 VSS.n370 VSS.n369 4.6505
R8136 VSS.n354 VSS.n353 4.6505
R8137 VSS.n340 VSS.n339 4.6505
R8138 VSS.n326 VSS.n325 4.6505
R8139 VSS.n309 VSS.n308 4.6505
R8140 VSS.n290 VSS.n289 4.6505
R8141 VSS.n3343 VSS.n3342 4.6505
R8142 VSS.n3373 VSS.n3372 4.6505
R8143 VSS.n3371 VSS.n3370 4.6505
R8144 VSS.n3365 VSS.n3364 4.6505
R8145 VSS.n3361 VSS.n3360 4.6505
R8146 VSS.n3355 VSS.n3354 4.6505
R8147 VSS.n3348 VSS.n3347 4.6505
R8148 VSS.n3346 VSS.n3345 4.6505
R8149 VSS.n3375 VSS.n3374 4.6505
R8150 VSS.n262 VSS.n261 4.46346
R8151 VSS.n2739 VSS.n2738 4.43314
R8152 VSS.n2387 VSS.n2386 4.43314
R8153 VSS.n948 VSS.n159 4.43314
R8154 VSS.n630 VSS.n204 4.43314
R8155 VSS.n312 VSS.n249 4.43314
R8156 VSS.n2993 VSS.n2992 4.42059
R8157 VSS.n2713 VSS.n2712 4.42059
R8158 VSS.n2641 VSS.n2640 4.42059
R8159 VSS.n2361 VSS.n2360 4.42059
R8160 VSS.n2289 VSS.n2288 4.42059
R8161 VSS.n4118 VSS.n27 4.42059
R8162 VSS.n4061 VSS.n40 4.42059
R8163 VSS.n4154 VSS.n4153 4.42059
R8164 VSS.n931 VSS.n169 4.42059
R8165 VSS.n875 VSS.n195 4.42059
R8166 VSS.n613 VSS.n214 4.42059
R8167 VSS.n557 VSS.n240 4.42059
R8168 VSS.n295 VSS.n259 4.42059
R8169 VSS.n2683 VSS.n2682 4.39476
R8170 VSS.n2331 VSS.n2330 4.39476
R8171 VSS.n3035 VSS.n3034 4.39476
R8172 VSS.n906 VSS.n185 4.39476
R8173 VSS.n588 VSS.n230 4.39476
R8174 VSS.n3127 VSS.n3126 4.1936
R8175 VSS.n1992 VSS 3.97291
R8176 VSS.n2107 VSS 3.97291
R8177 VSS.n1175 VSS.n1170 3.75222
R8178 VSS.n1165 VSS.n1160 3.75222
R8179 VSS.n1155 VSS.n1150 3.75222
R8180 VSS.n1206 VSS.n1201 3.75222
R8181 VSS.n1196 VSS.n1191 3.75222
R8182 VSS.n134 VSS.n133 3.75222
R8183 VSS.n1216 VSS.n140 3.75222
R8184 VSS.n1240 VSS.n1235 3.75222
R8185 VSS.n1322 VSS.n1317 3.75222
R8186 VSS.n1312 VSS.n1307 3.75222
R8187 VSS.n1302 VSS.n1297 3.75222
R8188 VSS.n1292 VSS.n1287 3.75222
R8189 VSS.n1280 VSS.n1275 3.75222
R8190 VSS.n1270 VSS.n1265 3.75222
R8191 VSS.n1260 VSS.n1255 3.75222
R8192 VSS.n1362 VSS.n1357 3.75222
R8193 VSS.n1352 VSS.n1347 3.75222
R8194 VSS.n1342 VSS.n1337 3.75222
R8195 VSS.n3416 VSS 3.53153
R8196 VSS.n3905 VSS 3.53153
R8197 VSS.n1222 VSS 3.53153
R8198 VSS.n4281 VSS 3.53153
R8199 VSS.n3536 VSS 3.53153
R8200 VSS.n3650 VSS 3.53153
R8201 VSS.n3764 VSS 3.53153
R8202 VSS.n3885 VSS 3.53153
R8203 VSS.n148 VSS.n145 3.42435
R8204 VSS.n3370 VSS.n3367 3.33963
R8205 VSS.n3430 VSS 3.31084
R8206 VSS.n3891 VSS 3.31084
R8207 VSS.n359 VSS.n358 3.31084
R8208 VSS.n677 VSS.n676 3.31084
R8209 VSS.n995 VSS.n994 3.31084
R8210 VSS.n1287 VSS.n1286 3.31084
R8211 VSS.n294 VSS.n266 3.19691
R8212 VSS.n3256 VSS.t349 3.1866
R8213 VSS.n2330 VSS.n2329 3.11687
R8214 VSS.n2682 VSS.n2681 3.11687
R8215 VSS.n3034 VSS.n3033 3.11687
R8216 VSS.n230 VSS.n228 3.11687
R8217 VSS.n185 VSS.n183 3.11687
R8218 VSS.n3430 VSS.n3429 3.1005
R8219 VSS.n3900 VSS.n3899 3.1005
R8220 VSS.n3892 VSS.n3891 3.1005
R8221 VSS.n3906 VSS.n3905 3.1005
R8222 VSS.n3912 VSS.n3911 3.1005
R8223 VSS.n3916 VSS.n3915 3.1005
R8224 VSS.n3927 VSS.n3924 3.1005
R8225 VSS.n1407 VSS.n1406 3.1005
R8226 VSS.n1485 VSS.n1484 3.1005
R8227 VSS.n1987 VSS.n1986 3.1005
R8228 VSS.n1977 VSS.n1976 3.1005
R8229 VSS.n1972 VSS.n1971 3.1005
R8230 VSS.n1968 VSS.n1967 3.1005
R8231 VSS.n1964 VSS.n1963 3.1005
R8232 VSS.n1960 VSS.n1959 3.1005
R8233 VSS.n1954 VSS.n1953 3.1005
R8234 VSS.n1950 VSS.n1949 3.1005
R8235 VSS.n1946 VSS.n1945 3.1005
R8236 VSS.n1942 VSS.n1941 3.1005
R8237 VSS.n1937 VSS.n1936 3.1005
R8238 VSS.n1933 VSS.n1932 3.1005
R8239 VSS.n1929 VSS.n1928 3.1005
R8240 VSS.n1925 VSS.n1924 3.1005
R8241 VSS.n1921 VSS.n1920 3.1005
R8242 VSS.n1915 VSS.n1914 3.1005
R8243 VSS.n1911 VSS.n1910 3.1005
R8244 VSS.n1907 VSS.n1906 3.1005
R8245 VSS.n1903 VSS.n1902 3.1005
R8246 VSS.n1898 VSS.n1897 3.1005
R8247 VSS.n1894 VSS.n1893 3.1005
R8248 VSS.n1889 VSS.n1888 3.1005
R8249 VSS.n1885 VSS.n1422 3.1005
R8250 VSS.n1876 VSS.n1875 3.1005
R8251 VSS.n1871 VSS.n1870 3.1005
R8252 VSS.n1867 VSS.n1866 3.1005
R8253 VSS.n1863 VSS.n1862 3.1005
R8254 VSS.n1859 VSS.n1858 3.1005
R8255 VSS.n1853 VSS.n1852 3.1005
R8256 VSS.n1849 VSS.n1848 3.1005
R8257 VSS.n1845 VSS.n1844 3.1005
R8258 VSS.n1841 VSS.n1840 3.1005
R8259 VSS.n1836 VSS.n1835 3.1005
R8260 VSS.n1832 VSS.n1831 3.1005
R8261 VSS.n1828 VSS.n1827 3.1005
R8262 VSS.n1824 VSS.n1823 3.1005
R8263 VSS.n1820 VSS.n1819 3.1005
R8264 VSS.n1814 VSS.n1813 3.1005
R8265 VSS.n1810 VSS.n1809 3.1005
R8266 VSS.n1806 VSS.n1805 3.1005
R8267 VSS.n1802 VSS.n1801 3.1005
R8268 VSS.n1797 VSS.n1796 3.1005
R8269 VSS.n1793 VSS.n1792 3.1005
R8270 VSS.n1788 VSS.n1787 3.1005
R8271 VSS.n1784 VSS.n1437 3.1005
R8272 VSS.n1775 VSS.n1774 3.1005
R8273 VSS.n1770 VSS.n1769 3.1005
R8274 VSS.n1766 VSS.n1765 3.1005
R8275 VSS.n1762 VSS.n1761 3.1005
R8276 VSS.n1758 VSS.n1757 3.1005
R8277 VSS.n1752 VSS.n1751 3.1005
R8278 VSS.n1748 VSS.n1747 3.1005
R8279 VSS.n1744 VSS.n1743 3.1005
R8280 VSS.n1740 VSS.n1739 3.1005
R8281 VSS.n1735 VSS.n1734 3.1005
R8282 VSS.n1731 VSS.n1730 3.1005
R8283 VSS.n1727 VSS.n1726 3.1005
R8284 VSS.n1723 VSS.n1722 3.1005
R8285 VSS.n1719 VSS.n1718 3.1005
R8286 VSS.n1713 VSS.n1712 3.1005
R8287 VSS.n1709 VSS.n1708 3.1005
R8288 VSS.n1705 VSS.n1704 3.1005
R8289 VSS.n1701 VSS.n1700 3.1005
R8290 VSS.n1696 VSS.n1695 3.1005
R8291 VSS.n1692 VSS.n1691 3.1005
R8292 VSS.n1687 VSS.n1686 3.1005
R8293 VSS.n1683 VSS.n1452 3.1005
R8294 VSS.n1674 VSS.n1673 3.1005
R8295 VSS.n1669 VSS.n1668 3.1005
R8296 VSS.n1665 VSS.n1664 3.1005
R8297 VSS.n1661 VSS.n1660 3.1005
R8298 VSS.n1657 VSS.n1656 3.1005
R8299 VSS.n1651 VSS.n1650 3.1005
R8300 VSS.n1647 VSS.n1646 3.1005
R8301 VSS.n1643 VSS.n1642 3.1005
R8302 VSS.n1639 VSS.n1638 3.1005
R8303 VSS.n1634 VSS.n1633 3.1005
R8304 VSS.n1630 VSS.n1629 3.1005
R8305 VSS.n1626 VSS.n1625 3.1005
R8306 VSS.n1622 VSS.n1621 3.1005
R8307 VSS.n1618 VSS.n1617 3.1005
R8308 VSS.n1612 VSS.n1611 3.1005
R8309 VSS.n1608 VSS.n1607 3.1005
R8310 VSS.n1604 VSS.n1603 3.1005
R8311 VSS.n1600 VSS.n1599 3.1005
R8312 VSS.n1595 VSS.n1594 3.1005
R8313 VSS.n1591 VSS.n1590 3.1005
R8314 VSS.n1586 VSS.n1585 3.1005
R8315 VSS.n1582 VSS.n1467 3.1005
R8316 VSS.n1573 VSS.n1572 3.1005
R8317 VSS.n1568 VSS.n1567 3.1005
R8318 VSS.n1564 VSS.n1563 3.1005
R8319 VSS.n1560 VSS.n1559 3.1005
R8320 VSS.n1556 VSS.n1555 3.1005
R8321 VSS.n1550 VSS.n1549 3.1005
R8322 VSS.n1546 VSS.n1545 3.1005
R8323 VSS.n1542 VSS.n1541 3.1005
R8324 VSS.n1538 VSS.n1537 3.1005
R8325 VSS.n1533 VSS.n1532 3.1005
R8326 VSS.n1529 VSS.n1528 3.1005
R8327 VSS.n1525 VSS.n1524 3.1005
R8328 VSS.n1521 VSS.n1520 3.1005
R8329 VSS.n1517 VSS.n1516 3.1005
R8330 VSS.n1511 VSS.n1510 3.1005
R8331 VSS.n1507 VSS.n1506 3.1005
R8332 VSS.n1503 VSS.n1502 3.1005
R8333 VSS.n1499 VSS.n1498 3.1005
R8334 VSS.n1494 VSS.n1493 3.1005
R8335 VSS.n1490 VSS.n1489 3.1005
R8336 VSS.n3397 VSS.n3396 3.1005
R8337 VSS.n3408 VSS.n3407 3.1005
R8338 VSS.n3414 VSS.n3413 3.1005
R8339 VSS.n3416 VSS.n3415 3.1005
R8340 VSS.n3422 VSS.n3421 3.1005
R8341 VSS.n1401 VSS.n1400 3.1005
R8342 VSS.n1392 VSS.n1391 3.1005
R8343 VSS.n1384 VSS.n1383 3.1005
R8344 VSS.n1380 VSS.n1379 3.1005
R8345 VSS.n1370 VSS.n1369 3.1005
R8346 VSS.n1366 VSS.n1365 3.1005
R8347 VSS.n1356 VSS.n1355 3.1005
R8348 VSS.n1336 VSS.n1335 3.1005
R8349 VSS.n1326 VSS.n1325 3.1005
R8350 VSS.n1316 VSS.n1315 3.1005
R8351 VSS.n1296 VSS.n1295 3.1005
R8352 VSS.n1284 VSS.n1283 3.1005
R8353 VSS.n1274 VSS.n1273 3.1005
R8354 VSS.n1244 VSS.n1243 3.1005
R8355 VSS.n1215 VSS.n1212 3.1005
R8356 VSS.n1210 VSS.n1209 3.1005
R8357 VSS.n1179 VSS.n1178 3.1005
R8358 VSS.n1169 VSS.n1168 3.1005
R8359 VSS.n287 VSS.n278 3.1005
R8360 VSS.n80 VSS.n79 3.1005
R8361 VSS.n3337 VSS.n3336 3.1005
R8362 VSS.n1159 VSS.n1158 3.1005
R8363 VSS.n1200 VSS.n1199 3.1005
R8364 VSS.n1223 VSS.n1222 3.1005
R8365 VSS.n1264 VSS.n1263 3.1005
R8366 VSS.n1306 VSS.n1305 3.1005
R8367 VSS.n1346 VSS.n1345 3.1005
R8368 VSS.n1376 VSS.n1375 3.1005
R8369 VSS.n1388 VSS.n1387 3.1005
R8370 VSS.n1397 VSS.n1396 3.1005
R8371 VSS.n2004 VSS.n2003 3.1005
R8372 VSS.n2013 VSS.n2012 3.1005
R8373 VSS.n2017 VSS.n2016 3.1005
R8374 VSS.n2021 VSS.n2020 3.1005
R8375 VSS.n2027 VSS.n2026 3.1005
R8376 VSS.n2031 VSS.n2030 3.1005
R8377 VSS.n2035 VSS.n2034 3.1005
R8378 VSS.n2039 VSS.n2038 3.1005
R8379 VSS.n2044 VSS.n2043 3.1005
R8380 VSS.n2048 VSS.n2047 3.1005
R8381 VSS.n2052 VSS.n2051 3.1005
R8382 VSS.n2056 VSS.n2055 3.1005
R8383 VSS.n2060 VSS.n2059 3.1005
R8384 VSS.n2066 VSS.n2065 3.1005
R8385 VSS.n2070 VSS.n2069 3.1005
R8386 VSS.n2074 VSS.n2073 3.1005
R8387 VSS.n2078 VSS.n2077 3.1005
R8388 VSS.n2082 VSS.n2081 3.1005
R8389 VSS.n2092 VSS.n2091 3.1005
R8390 VSS.n2096 VSS.n2095 3.1005
R8391 VSS.n2106 VSS.n2103 3.1005
R8392 VSS.n2107 VSS.n122 3.1005
R8393 VSS.n2119 VSS.n2118 3.1005
R8394 VSS.n2128 VSS.n2127 3.1005
R8395 VSS.n2132 VSS.n2131 3.1005
R8396 VSS.n2136 VSS.n2135 3.1005
R8397 VSS.n2142 VSS.n2141 3.1005
R8398 VSS.n2146 VSS.n2145 3.1005
R8399 VSS.n2150 VSS.n2149 3.1005
R8400 VSS.n2154 VSS.n2153 3.1005
R8401 VSS.n2159 VSS.n2158 3.1005
R8402 VSS.n2163 VSS.n2162 3.1005
R8403 VSS.n1992 VSS.n1990 3.1005
R8404 VSS.n4173 VSS.n4172 3.1005
R8405 VSS.n3885 VSS.n3884 3.1005
R8406 VSS.n3877 VSS.n3876 3.1005
R8407 VSS.n3868 VSS.n3867 3.1005
R8408 VSS.n3864 VSS.n3863 3.1005
R8409 VSS.n3860 VSS.n3859 3.1005
R8410 VSS.n3856 VSS.n3855 3.1005
R8411 VSS.n3850 VSS.n3849 3.1005
R8412 VSS.n3846 VSS.n3845 3.1005
R8413 VSS.n3842 VSS.n3841 3.1005
R8414 VSS.n3838 VSS.n3837 3.1005
R8415 VSS.n3833 VSS.n3832 3.1005
R8416 VSS.n3829 VSS.n3828 3.1005
R8417 VSS.n3825 VSS.n3824 3.1005
R8418 VSS.n3821 VSS.n3820 3.1005
R8419 VSS.n3817 VSS.n3816 3.1005
R8420 VSS.n3811 VSS.n3810 3.1005
R8421 VSS.n3807 VSS.n3806 3.1005
R8422 VSS.n3803 VSS.n3802 3.1005
R8423 VSS.n3799 VSS.n3798 3.1005
R8424 VSS.n3789 VSS.n3788 3.1005
R8425 VSS.n3785 VSS.n3784 3.1005
R8426 VSS.n3775 VSS.n3774 3.1005
R8427 VSS.n3765 VSS.n3764 3.1005
R8428 VSS.n3763 VSS.n3762 3.1005
R8429 VSS.n3754 VSS.n3753 3.1005
R8430 VSS.n3750 VSS.n3749 3.1005
R8431 VSS.n3746 VSS.n3745 3.1005
R8432 VSS.n3742 VSS.n3741 3.1005
R8433 VSS.n3736 VSS.n3735 3.1005
R8434 VSS.n3732 VSS.n3731 3.1005
R8435 VSS.n3728 VSS.n3727 3.1005
R8436 VSS.n3724 VSS.n3723 3.1005
R8437 VSS.n3719 VSS.n3718 3.1005
R8438 VSS.n3715 VSS.n3714 3.1005
R8439 VSS.n3711 VSS.n3710 3.1005
R8440 VSS.n3707 VSS.n3706 3.1005
R8441 VSS.n3703 VSS.n3702 3.1005
R8442 VSS.n3697 VSS.n3696 3.1005
R8443 VSS.n3693 VSS.n3692 3.1005
R8444 VSS.n3689 VSS.n3688 3.1005
R8445 VSS.n3685 VSS.n3684 3.1005
R8446 VSS.n3675 VSS.n3674 3.1005
R8447 VSS.n3671 VSS.n3670 3.1005
R8448 VSS.n3661 VSS.n3660 3.1005
R8449 VSS.n3651 VSS.n3650 3.1005
R8450 VSS.n3649 VSS.n3648 3.1005
R8451 VSS.n3640 VSS.n3639 3.1005
R8452 VSS.n3636 VSS.n3635 3.1005
R8453 VSS.n3632 VSS.n3631 3.1005
R8454 VSS.n3628 VSS.n3627 3.1005
R8455 VSS.n3622 VSS.n3621 3.1005
R8456 VSS.n3618 VSS.n3617 3.1005
R8457 VSS.n3614 VSS.n3613 3.1005
R8458 VSS.n3610 VSS.n3609 3.1005
R8459 VSS.n3605 VSS.n3604 3.1005
R8460 VSS.n3601 VSS.n3600 3.1005
R8461 VSS.n3597 VSS.n3596 3.1005
R8462 VSS.n3593 VSS.n3592 3.1005
R8463 VSS.n3589 VSS.n3588 3.1005
R8464 VSS.n3583 VSS.n3582 3.1005
R8465 VSS.n3579 VSS.n3578 3.1005
R8466 VSS.n3575 VSS.n3574 3.1005
R8467 VSS.n3571 VSS.n3570 3.1005
R8468 VSS.n3561 VSS.n3560 3.1005
R8469 VSS.n3557 VSS.n3556 3.1005
R8470 VSS.n3547 VSS.n3546 3.1005
R8471 VSS.n3537 VSS.n3536 3.1005
R8472 VSS.n3535 VSS.n3534 3.1005
R8473 VSS.n3526 VSS.n3525 3.1005
R8474 VSS.n3522 VSS.n3521 3.1005
R8475 VSS.n3518 VSS.n3517 3.1005
R8476 VSS.n3514 VSS.n3513 3.1005
R8477 VSS.n3508 VSS.n3507 3.1005
R8478 VSS.n3504 VSS.n3503 3.1005
R8479 VSS.n3500 VSS.n3499 3.1005
R8480 VSS.n3496 VSS.n3495 3.1005
R8481 VSS.n3491 VSS.n3490 3.1005
R8482 VSS.n3487 VSS.n3486 3.1005
R8483 VSS.n3483 VSS.n3482 3.1005
R8484 VSS.n3479 VSS.n3478 3.1005
R8485 VSS.n3475 VSS.n3474 3.1005
R8486 VSS.n3469 VSS.n3468 3.1005
R8487 VSS.n3465 VSS.n3464 3.1005
R8488 VSS.n3461 VSS.n3460 3.1005
R8489 VSS.n3457 VSS.n3456 3.1005
R8490 VSS.n3447 VSS.n3446 3.1005
R8491 VSS.n3443 VSS.n3442 3.1005
R8492 VSS.n4287 VSS.n4286 3.1005
R8493 VSS.n4281 VSS.n0 3.1005
R8494 VSS.n4275 VSS.n4274 3.1005
R8495 VSS.n4266 VSS.n4265 3.1005
R8496 VSS.n4262 VSS.n4261 3.1005
R8497 VSS.n4258 VSS.n4257 3.1005
R8498 VSS.n4254 VSS.n4253 3.1005
R8499 VSS.n4248 VSS.n4247 3.1005
R8500 VSS.n4244 VSS.n4243 3.1005
R8501 VSS.n4240 VSS.n4239 3.1005
R8502 VSS.n4236 VSS.n4235 3.1005
R8503 VSS.n4231 VSS.n4230 3.1005
R8504 VSS.n4227 VSS.n4226 3.1005
R8505 VSS.n4223 VSS.n4222 3.1005
R8506 VSS.n4219 VSS.n4218 3.1005
R8507 VSS.n4215 VSS.n4214 3.1005
R8508 VSS.n4209 VSS.n4208 3.1005
R8509 VSS.n4205 VSS.n4204 3.1005
R8510 VSS.n4201 VSS.n4200 3.1005
R8511 VSS.n4197 VSS.n4196 3.1005
R8512 VSS.n4187 VSS.n4186 3.1005
R8513 VSS.n4183 VSS.n4182 3.1005
R8514 VSS.n4162 VSS.n4161 3.09016
R8515 VSS.n4142 VSS.n4135 3.09016
R8516 VSS.n4144 VSS.n4142 3.09016
R8517 VSS.n4128 VSS.n4122 3.09016
R8518 VSS.n4130 VSS.n4128 3.09016
R8519 VSS.n4114 VSS.n4112 3.09016
R8520 VSS.n4100 VSS.n4093 3.09016
R8521 VSS.n4102 VSS.n4100 3.09016
R8522 VSS.n4086 VSS.n4079 3.09016
R8523 VSS.n4088 VSS.n4086 3.09016
R8524 VSS.n4072 VSS.n4065 3.09016
R8525 VSS.n4074 VSS.n4072 3.09016
R8526 VSS.n36 VSS.n29 3.09016
R8527 VSS.n4057 VSS.n4055 3.09016
R8528 VSS.n4043 VSS.n4036 3.09016
R8529 VSS.n4045 VSS.n4043 3.09016
R8530 VSS.n4029 VSS.n4022 3.09016
R8531 VSS.n4031 VSS.n4029 3.09016
R8532 VSS.n4015 VSS.n4008 3.09016
R8533 VSS.n4017 VSS.n4015 3.09016
R8534 VSS.n4000 VSS.n3993 3.09016
R8535 VSS.n4003 VSS.n4000 3.09016
R8536 VSS.n3986 VSS.n3979 3.09016
R8537 VSS.n3988 VSS.n3986 3.09016
R8538 VSS.n3971 VSS.n3964 3.09016
R8539 VSS.n3974 VSS.n3971 3.09016
R8540 VSS.n3957 VSS.n3950 3.09016
R8541 VSS.n3959 VSS.n3957 3.09016
R8542 VSS.n50 VSS.n43 3.09016
R8543 VSS.n3945 VSS.n50 3.09016
R8544 VSS.n1186 VSS.n1185 2.99827
R8545 VSS.n1230 VSS.n1229 2.99827
R8546 VSS.n3354 VSS 2.96862
R8547 VSS.n1251 VSS.n1250 2.8978
R8548 VSS.n26 VSS.n17 2.86947
R8549 VSS.n2288 VSS.n2287 2.7891
R8550 VSS.n2360 VSS.n2359 2.7891
R8551 VSS.n2640 VSS.n2639 2.7891
R8552 VSS.n2712 VSS.n2711 2.7891
R8553 VSS.n2992 VSS.n2991 2.7891
R8554 VSS.n4164 VSS.n4154 2.7891
R8555 VSS.n27 VSS.n26 2.7891
R8556 VSS.n40 VSS.n39 2.7891
R8557 VSS.n259 VSS.n258 2.7891
R8558 VSS.n240 VSS.n239 2.7891
R8559 VSS.n214 VSS.n213 2.7891
R8560 VSS.n195 VSS.n194 2.7891
R8561 VSS.n169 VSS.n168 2.7891
R8562 VSS.n2043 VSS.n2040 2.64878
R8563 VSS.n2158 VSS.n2155 2.64878
R8564 VSS.n2209 VSS.n2208 2.64878
R8565 VSS.n2561 VSS.n2560 2.64878
R8566 VSS.n2913 VSS.n2912 2.64878
R8567 VSS.n1941 VSS.n1938 2.64878
R8568 VSS.n1840 VSS.n1837 2.64878
R8569 VSS.n1739 VSS.n1736 2.64878
R8570 VSS.n1638 VSS.n1635 2.64878
R8571 VSS.n1537 VSS.n1534 2.64878
R8572 VSS.n4235 VSS.n4232 2.64878
R8573 VSS.n3495 VSS.n3492 2.64878
R8574 VSS.n3609 VSS.n3606 2.64878
R8575 VSS.n3723 VSS.n3720 2.64878
R8576 VSS.n3837 VSS.n3834 2.64878
R8577 VSS.n2386 VSS.n2385 2.63101
R8578 VSS.n2738 VSS.n2737 2.63101
R8579 VSS.n249 VSS.n248 2.63101
R8580 VSS.n204 VSS.n203 2.63101
R8581 VSS.n159 VSS.n158 2.63101
R8582 VSS.n3341 VSS 2.5976
R8583 VSS.n2124 VSS.n2123 2.5203
R8584 VSS.n2009 VSS.n2008 2.5203
R8585 VSS.n1254 VSS.n1253 2.5203
R8586 VSS.n1569 VSS.n1471 2.5203
R8587 VSS.n1670 VSS.n1456 2.5203
R8588 VSS.n1771 VSS.n1441 2.5203
R8589 VSS.n1872 VSS.n1426 2.5203
R8590 VSS.n1973 VSS.n1411 2.5203
R8591 VSS.n3873 VSS.n3872 2.5203
R8592 VSS.n3759 VSS.n3758 2.5203
R8593 VSS.n3645 VSS.n3644 2.5203
R8594 VSS.n3531 VSS.n3530 2.5203
R8595 VSS.n4271 VSS.n4270 2.5203
R8596 VSS.n3428 VSS.n3427 2.49102
R8597 VSS.n3404 VSS.n3403 2.49102
R8598 VSS.n2115 VSS.n2114 2.49102
R8599 VSS.n2088 VSS.n2087 2.49102
R8600 VSS.n2000 VSS.n1999 2.49102
R8601 VSS.n3922 VSS.n3921 2.49102
R8602 VSS.n3898 VSS.n3897 2.49102
R8603 VSS.n1234 VSS.n1233 2.49102
R8604 VSS.n1190 VSS.n1189 2.49102
R8605 VSS.n1393 VSS.n132 2.49102
R8606 VSS.n1495 VSS.n1476 2.49102
R8607 VSS.n1576 VSS.n1574 2.49102
R8608 VSS.n1596 VSS.n1461 2.49102
R8609 VSS.n1677 VSS.n1675 2.49102
R8610 VSS.n1697 VSS.n1446 2.49102
R8611 VSS.n1778 VSS.n1776 2.49102
R8612 VSS.n1798 VSS.n1431 2.49102
R8613 VSS.n1879 VSS.n1877 2.49102
R8614 VSS.n1899 VSS.n1416 2.49102
R8615 VSS.n1980 VSS.n1978 2.49102
R8616 VSS.n3883 VSS.n3882 2.49102
R8617 VSS.n3795 VSS.n3794 2.49102
R8618 VSS.n3767 VSS.n3766 2.49102
R8619 VSS.n3681 VSS.n3680 2.49102
R8620 VSS.n3653 VSS.n3652 2.49102
R8621 VSS.n3567 VSS.n3566 2.49102
R8622 VSS.n3539 VSS.n3538 2.49102
R8623 VSS.n3453 VSS.n3452 2.49102
R8624 VSS.n4277 VSS.n4276 2.49102
R8625 VSS.n4193 VSS.n4192 2.49102
R8626 VSS.n2102 VSS.n2101 2.43201
R8627 VSS.n1211 VSS.n150 2.43201
R8628 VSS.n1402 VSS.n127 2.43201
R8629 VSS.n1486 VSS.n1481 2.43201
R8630 VSS.n1587 VSS.n1466 2.43201
R8631 VSS.n1688 VSS.n1451 2.43201
R8632 VSS.n1789 VSS.n1436 2.43201
R8633 VSS.n1890 VSS.n1421 2.43201
R8634 VSS.n3781 VSS.n3780 2.43201
R8635 VSS.n3667 VSS.n3666 2.43201
R8636 VSS.n3553 VSS.n3552 2.43201
R8637 VSS.n6 VSS.n5 2.43201
R8638 VSS.n4179 VSS.n4178 2.43201
R8639 VSS.n121 VSS 2.42809
R8640 VSS.n110 VSS 2.42809
R8641 VSS.n291 VSS.n273 2.38818
R8642 VSS.n3374 VSS 2.29155
R8643 VSS.n273 VSS 2.2358
R8644 VSS.n2173 VSS.n2166 2.2074
R8645 VSS.n2175 VSS.n2173 2.2074
R8646 VSS.n2187 VSS.n2180 2.2074
R8647 VSS.n2189 VSS.n2187 2.2074
R8648 VSS.n2201 VSS.n2194 2.2074
R8649 VSS.n2203 VSS.n2201 2.2074
R8650 VSS.n2217 VSS.n2210 2.2074
R8651 VSS.n2219 VSS.n2217 2.2074
R8652 VSS.n2231 VSS.n2224 2.2074
R8653 VSS.n2233 VSS.n2231 2.2074
R8654 VSS.n2245 VSS.n2238 2.2074
R8655 VSS.n2247 VSS.n2245 2.2074
R8656 VSS.n2259 VSS.n2252 2.2074
R8657 VSS.n2261 VSS.n2259 2.2074
R8658 VSS.n2273 VSS.n2266 2.2074
R8659 VSS.n2275 VSS.n2273 2.2074
R8660 VSS.n2300 VSS.n2293 2.2074
R8661 VSS.n2302 VSS.n2300 2.2074
R8662 VSS.n2314 VSS.n2307 2.2074
R8663 VSS.n2316 VSS.n2314 2.2074
R8664 VSS.n2342 VSS.n2335 2.2074
R8665 VSS.n2345 VSS.n2342 2.2074
R8666 VSS.n2352 VSS.n120 2.2074
R8667 VSS.n2352 VSS.n2351 2.2074
R8668 VSS.n2372 VSS.n2365 2.2074
R8669 VSS.n2374 VSS.n2372 2.2074
R8670 VSS.n2398 VSS.n2391 2.2074
R8671 VSS.n2400 VSS.n2398 2.2074
R8672 VSS.n2412 VSS.n2405 2.2074
R8673 VSS.n2414 VSS.n2412 2.2074
R8674 VSS.n2426 VSS.n2419 2.2074
R8675 VSS.n2428 VSS.n2426 2.2074
R8676 VSS.n2439 VSS.n2433 2.2074
R8677 VSS.n2443 VSS.n2439 2.2074
R8678 VSS.n2455 VSS.n2448 2.2074
R8679 VSS.n2457 VSS.n2455 2.2074
R8680 VSS.n2469 VSS.n2462 2.2074
R8681 VSS.n2471 VSS.n2469 2.2074
R8682 VSS.n2483 VSS.n2476 2.2074
R8683 VSS.n2485 VSS.n2483 2.2074
R8684 VSS.n2497 VSS.n2490 2.2074
R8685 VSS.n2500 VSS.n2497 2.2074
R8686 VSS.n2513 VSS.n2511 2.2074
R8687 VSS.n2525 VSS.n2518 2.2074
R8688 VSS.n2527 VSS.n2525 2.2074
R8689 VSS.n2539 VSS.n2532 2.2074
R8690 VSS.n2541 VSS.n2539 2.2074
R8691 VSS.n2553 VSS.n2546 2.2074
R8692 VSS.n2555 VSS.n2553 2.2074
R8693 VSS.n2569 VSS.n2562 2.2074
R8694 VSS.n2571 VSS.n2569 2.2074
R8695 VSS.n2583 VSS.n2576 2.2074
R8696 VSS.n2585 VSS.n2583 2.2074
R8697 VSS.n2597 VSS.n2590 2.2074
R8698 VSS.n2599 VSS.n2597 2.2074
R8699 VSS.n2611 VSS.n2604 2.2074
R8700 VSS.n2613 VSS.n2611 2.2074
R8701 VSS.n2625 VSS.n2618 2.2074
R8702 VSS.n2627 VSS.n2625 2.2074
R8703 VSS.n2652 VSS.n2645 2.2074
R8704 VSS.n2654 VSS.n2652 2.2074
R8705 VSS.n2666 VSS.n2659 2.2074
R8706 VSS.n2668 VSS.n2666 2.2074
R8707 VSS.n2694 VSS.n2687 2.2074
R8708 VSS.n2697 VSS.n2694 2.2074
R8709 VSS.n2704 VSS.n109 2.2074
R8710 VSS.n2704 VSS.n2703 2.2074
R8711 VSS.n2724 VSS.n2717 2.2074
R8712 VSS.n2726 VSS.n2724 2.2074
R8713 VSS.n2750 VSS.n2743 2.2074
R8714 VSS.n2752 VSS.n2750 2.2074
R8715 VSS.n2764 VSS.n2757 2.2074
R8716 VSS.n2766 VSS.n2764 2.2074
R8717 VSS.n2778 VSS.n2771 2.2074
R8718 VSS.n2780 VSS.n2778 2.2074
R8719 VSS.n2791 VSS.n2785 2.2074
R8720 VSS.n2795 VSS.n2791 2.2074
R8721 VSS.n2807 VSS.n2800 2.2074
R8722 VSS.n2809 VSS.n2807 2.2074
R8723 VSS.n2821 VSS.n2814 2.2074
R8724 VSS.n2823 VSS.n2821 2.2074
R8725 VSS.n2835 VSS.n2828 2.2074
R8726 VSS.n2837 VSS.n2835 2.2074
R8727 VSS.n2849 VSS.n2842 2.2074
R8728 VSS.n2852 VSS.n2849 2.2074
R8729 VSS.n2865 VSS.n2863 2.2074
R8730 VSS.n2877 VSS.n2870 2.2074
R8731 VSS.n2879 VSS.n2877 2.2074
R8732 VSS.n2891 VSS.n2884 2.2074
R8733 VSS.n2893 VSS.n2891 2.2074
R8734 VSS.n2905 VSS.n2898 2.2074
R8735 VSS.n2907 VSS.n2905 2.2074
R8736 VSS.n2921 VSS.n2914 2.2074
R8737 VSS.n2923 VSS.n2921 2.2074
R8738 VSS.n2935 VSS.n2928 2.2074
R8739 VSS.n2937 VSS.n2935 2.2074
R8740 VSS.n2949 VSS.n2942 2.2074
R8741 VSS.n2951 VSS.n2949 2.2074
R8742 VSS.n2963 VSS.n2956 2.2074
R8743 VSS.n2965 VSS.n2963 2.2074
R8744 VSS.n2977 VSS.n2970 2.2074
R8745 VSS.n2979 VSS.n2977 2.2074
R8746 VSS.n3004 VSS.n2997 2.2074
R8747 VSS.n3006 VSS.n3004 2.2074
R8748 VSS.n3018 VSS.n3011 2.2074
R8749 VSS.n3020 VSS.n3018 2.2074
R8750 VSS.n99 VSS.n92 2.2074
R8751 VSS.n3040 VSS.n99 2.2074
R8752 VSS.n3050 VSS.n3043 2.2074
R8753 VSS.n3053 VSS.n3050 2.2074
R8754 VSS.n3067 VSS.n3065 2.2074
R8755 VSS.n3079 VSS.n3072 2.2074
R8756 VSS.n3081 VSS.n3079 2.2074
R8757 VSS.n3329 VSS.n88 2.2074
R8758 VSS.n3329 VSS.n3328 2.2074
R8759 VSS.n3319 VSS.n3312 2.2074
R8760 VSS.n3323 VSS.n3319 2.2074
R8761 VSS.n3305 VSS.n3298 2.2074
R8762 VSS.n3307 VSS.n3305 2.2074
R8763 VSS.n3289 VSS.n3282 2.2074
R8764 VSS.n3293 VSS.n3289 2.2074
R8765 VSS.n3275 VSS.n3269 2.2074
R8766 VSS.n3277 VSS.n3275 2.2074
R8767 VSS.n3260 VSS.n3253 2.2074
R8768 VSS.n3264 VSS.n3260 2.2074
R8769 VSS.n3246 VSS.n3239 2.2074
R8770 VSS.n3248 VSS.n3246 2.2074
R8771 VSS.n3231 VSS.n3224 2.2074
R8772 VSS.n3216 VSS.n3209 2.2074
R8773 VSS.n3218 VSS.n3216 2.2074
R8774 VSS.n3204 VSS.n3202 2.2074
R8775 VSS.n3186 VSS.n3179 2.2074
R8776 VSS.n3188 VSS.n3186 2.2074
R8777 VSS.n3172 VSS.n3165 2.2074
R8778 VSS.n3174 VSS.n3172 2.2074
R8779 VSS.n3154 VSS.n3147 2.2074
R8780 VSS.n3158 VSS.n3154 2.2074
R8781 VSS.n3140 VSS.n3133 2.2074
R8782 VSS.n3142 VSS.n3140 2.2074
R8783 VSS.n3124 VSS.n3117 2.2074
R8784 VSS.n3128 VSS.n3124 2.2074
R8785 VSS.n3110 VSS.n3103 2.2074
R8786 VSS.n3112 VSS.n3110 2.2074
R8787 VSS.n3094 VSS.n3087 2.2074
R8788 VSS.n3098 VSS.n3094 2.2074
R8789 VSS.n3381 VSS.n69 2.2074
R8790 VSS.n3383 VSS.n3381 2.2074
R8791 VSS.n3391 VSS.n66 2.2074
R8792 VSS.n26 VSS.n25 2.2074
R8793 VSS.n277 VSS.n276 2.2074
R8794 VSS.n306 VSS.n299 2.2074
R8795 VSS.n409 VSS.n402 2.2074
R8796 VSS.n395 VSS.n388 2.2074
R8797 VSS.n381 VSS.n374 2.2074
R8798 VSS.n367 VSS.n360 2.2074
R8799 VSS.n351 VSS.n344 2.2074
R8800 VSS.n337 VSS.n330 2.2074
R8801 VSS.n323 VSS.n316 2.2074
R8802 VSS.n551 VSS.n544 2.2074
R8803 VSS.n537 VSS.n530 2.2074
R8804 VSS.n523 VSS.n516 2.2074
R8805 VSS.n509 VSS.n502 2.2074
R8806 VSS.n493 VSS.n486 2.2074
R8807 VSS.n479 VSS.n472 2.2074
R8808 VSS.n465 VSS.n458 2.2074
R8809 VSS.n451 VSS.n444 2.2074
R8810 VSS.n437 VSS.n430 2.2074
R8811 VSS.n582 VSS.n575 2.2074
R8812 VSS.n568 VSS.n561 2.2074
R8813 VSS.n218 VSS.n217 2.2074
R8814 VSS.n606 VSS.n605 2.2074
R8815 VSS.n624 VSS.n617 2.2074
R8816 VSS.n727 VSS.n720 2.2074
R8817 VSS.n713 VSS.n706 2.2074
R8818 VSS.n699 VSS.n692 2.2074
R8819 VSS.n685 VSS.n678 2.2074
R8820 VSS.n669 VSS.n662 2.2074
R8821 VSS.n655 VSS.n648 2.2074
R8822 VSS.n641 VSS.n634 2.2074
R8823 VSS.n869 VSS.n862 2.2074
R8824 VSS.n855 VSS.n848 2.2074
R8825 VSS.n841 VSS.n834 2.2074
R8826 VSS.n827 VSS.n820 2.2074
R8827 VSS.n811 VSS.n804 2.2074
R8828 VSS.n797 VSS.n790 2.2074
R8829 VSS.n783 VSS.n776 2.2074
R8830 VSS.n769 VSS.n762 2.2074
R8831 VSS.n755 VSS.n748 2.2074
R8832 VSS.n900 VSS.n893 2.2074
R8833 VSS.n886 VSS.n879 2.2074
R8834 VSS.n173 VSS.n172 2.2074
R8835 VSS.n924 VSS.n923 2.2074
R8836 VSS.n942 VSS.n935 2.2074
R8837 VSS.n1045 VSS.n1038 2.2074
R8838 VSS.n1031 VSS.n1024 2.2074
R8839 VSS.n1017 VSS.n1010 2.2074
R8840 VSS.n1003 VSS.n996 2.2074
R8841 VSS.n987 VSS.n980 2.2074
R8842 VSS.n973 VSS.n966 2.2074
R8843 VSS.n959 VSS.n952 2.2074
R8844 VSS.n1145 VSS.n1138 2.2074
R8845 VSS.n1129 VSS.n1122 2.2074
R8846 VSS.n1115 VSS.n1108 2.2074
R8847 VSS.n1101 VSS.n1094 2.2074
R8848 VSS.n1087 VSS.n1080 2.2074
R8849 VSS.n1073 VSS.n1066 2.2074
R8850 VSS.n3413 VSS.n3410 1.98671
R8851 VSS.n3911 VSS.n3908 1.98671
R8852 VSS.n289 VSS.n277 1.98671
R8853 VSS.n308 VSS.n306 1.98671
R8854 VSS.n425 VSS.n423 1.98671
R8855 VSS.n411 VSS.n409 1.98671
R8856 VSS.n397 VSS.n395 1.98671
R8857 VSS.n383 VSS.n381 1.98671
R8858 VSS.n369 VSS.n367 1.98671
R8859 VSS.n353 VSS.n351 1.98671
R8860 VSS.n339 VSS.n337 1.98671
R8861 VSS.n325 VSS.n323 1.98671
R8862 VSS.n553 VSS.n551 1.98671
R8863 VSS.n539 VSS.n537 1.98671
R8864 VSS.n525 VSS.n523 1.98671
R8865 VSS.n511 VSS.n509 1.98671
R8866 VSS.n497 VSS.n493 1.98671
R8867 VSS.n481 VSS.n479 1.98671
R8868 VSS.n467 VSS.n465 1.98671
R8869 VSS.n453 VSS.n451 1.98671
R8870 VSS.n439 VSS.n437 1.98671
R8871 VSS.n584 VSS.n582 1.98671
R8872 VSS.n570 VSS.n568 1.98671
R8873 VSS.n609 VSS.n218 1.98671
R8874 VSS.n605 VSS.n592 1.98671
R8875 VSS.n626 VSS.n624 1.98671
R8876 VSS.n743 VSS.n741 1.98671
R8877 VSS.n729 VSS.n727 1.98671
R8878 VSS.n715 VSS.n713 1.98671
R8879 VSS.n701 VSS.n699 1.98671
R8880 VSS.n687 VSS.n685 1.98671
R8881 VSS.n671 VSS.n669 1.98671
R8882 VSS.n657 VSS.n655 1.98671
R8883 VSS.n643 VSS.n641 1.98671
R8884 VSS.n871 VSS.n869 1.98671
R8885 VSS.n857 VSS.n855 1.98671
R8886 VSS.n843 VSS.n841 1.98671
R8887 VSS.n829 VSS.n827 1.98671
R8888 VSS.n815 VSS.n811 1.98671
R8889 VSS.n799 VSS.n797 1.98671
R8890 VSS.n785 VSS.n783 1.98671
R8891 VSS.n771 VSS.n769 1.98671
R8892 VSS.n757 VSS.n755 1.98671
R8893 VSS.n902 VSS.n900 1.98671
R8894 VSS.n888 VSS.n886 1.98671
R8895 VSS.n927 VSS.n173 1.98671
R8896 VSS.n923 VSS.n910 1.98671
R8897 VSS.n944 VSS.n942 1.98671
R8898 VSS.n1061 VSS.n1059 1.98671
R8899 VSS.n1047 VSS.n1045 1.98671
R8900 VSS.n1033 VSS.n1031 1.98671
R8901 VSS.n1019 VSS.n1017 1.98671
R8902 VSS.n1005 VSS.n1003 1.98671
R8903 VSS.n989 VSS.n987 1.98671
R8904 VSS.n975 VSS.n973 1.98671
R8905 VSS.n961 VSS.n959 1.98671
R8906 VSS.n1178 VSS.n1175 1.98671
R8907 VSS.n1168 VSS.n1165 1.98671
R8908 VSS.n1158 VSS.n1155 1.98671
R8909 VSS.n1147 VSS.n1145 1.98671
R8910 VSS.n1133 VSS.n1129 1.98671
R8911 VSS.n1117 VSS.n1115 1.98671
R8912 VSS.n1103 VSS.n1101 1.98671
R8913 VSS.n1089 VSS.n1087 1.98671
R8914 VSS.n1075 VSS.n1073 1.98671
R8915 VSS.n1209 VSS.n1206 1.98671
R8916 VSS.n1199 VSS.n1196 1.98671
R8917 VSS.n1222 VSS.n134 1.98671
R8918 VSS.n1216 VSS.n1215 1.98671
R8919 VSS.n1243 VSS.n1240 1.98671
R8920 VSS.n1335 VSS.n1332 1.98671
R8921 VSS.n1325 VSS.n1322 1.98671
R8922 VSS.n1315 VSS.n1312 1.98671
R8923 VSS.n1305 VSS.n1302 1.98671
R8924 VSS.n1295 VSS.n1292 1.98671
R8925 VSS.n1283 VSS.n1280 1.98671
R8926 VSS.n1273 VSS.n1270 1.98671
R8927 VSS.n1263 VSS.n1260 1.98671
R8928 VSS.n1365 VSS.n1362 1.98671
R8929 VSS.n1355 VSS.n1352 1.98671
R8930 VSS.n1345 VSS.n1342 1.98671
R8931 VSS.n268 VSS.n267 1.9836
R8932 VSS.n264 VSS.n263 1.87367
R8933 VSS.n3232 VSS.n3231 1.76602
R8934 VSS.n3202 VSS.n3195 1.76602
R8935 VSS.n39 VSS.n36 1.76602
R8936 VSS.n289 VSS.n288 1.76602
R8937 VSS.n288 VSS 1.76602
R8938 VSS.n308 VSS.n307 1.76602
R8939 VSS.n425 VSS.n424 1.76602
R8940 VSS.n411 VSS.n410 1.76602
R8941 VSS.n397 VSS.n396 1.76602
R8942 VSS.n383 VSS.n382 1.76602
R8943 VSS.n369 VSS.n368 1.76602
R8944 VSS.n353 VSS.n352 1.76602
R8945 VSS.n339 VSS.n338 1.76602
R8946 VSS.n325 VSS.n324 1.76602
R8947 VSS.n553 VSS.n552 1.76602
R8948 VSS.n539 VSS.n538 1.76602
R8949 VSS.n525 VSS.n524 1.76602
R8950 VSS.n511 VSS.n510 1.76602
R8951 VSS.n497 VSS.n496 1.76602
R8952 VSS.n481 VSS.n480 1.76602
R8953 VSS.n467 VSS.n466 1.76602
R8954 VSS.n453 VSS.n452 1.76602
R8955 VSS.n439 VSS.n438 1.76602
R8956 VSS.n584 VSS.n583 1.76602
R8957 VSS.n570 VSS.n569 1.76602
R8958 VSS.n609 VSS.n608 1.76602
R8959 VSS.n608 VSS 1.76602
R8960 VSS.n592 VSS.n219 1.76602
R8961 VSS.n626 VSS.n625 1.76602
R8962 VSS.n743 VSS.n742 1.76602
R8963 VSS.n729 VSS.n728 1.76602
R8964 VSS.n715 VSS.n714 1.76602
R8965 VSS.n701 VSS.n700 1.76602
R8966 VSS.n687 VSS.n686 1.76602
R8967 VSS.n671 VSS.n670 1.76602
R8968 VSS.n657 VSS.n656 1.76602
R8969 VSS.n643 VSS.n642 1.76602
R8970 VSS.n871 VSS.n870 1.76602
R8971 VSS.n857 VSS.n856 1.76602
R8972 VSS.n843 VSS.n842 1.76602
R8973 VSS.n829 VSS.n828 1.76602
R8974 VSS.n815 VSS.n814 1.76602
R8975 VSS.n799 VSS.n798 1.76602
R8976 VSS.n785 VSS.n784 1.76602
R8977 VSS.n771 VSS.n770 1.76602
R8978 VSS.n757 VSS.n756 1.76602
R8979 VSS.n902 VSS.n901 1.76602
R8980 VSS.n888 VSS.n887 1.76602
R8981 VSS.n927 VSS.n926 1.76602
R8982 VSS.n926 VSS 1.76602
R8983 VSS.n910 VSS.n174 1.76602
R8984 VSS.n944 VSS.n943 1.76602
R8985 VSS.n1061 VSS.n1060 1.76602
R8986 VSS.n1047 VSS.n1046 1.76602
R8987 VSS.n1033 VSS.n1032 1.76602
R8988 VSS.n1019 VSS.n1018 1.76602
R8989 VSS.n1005 VSS.n1004 1.76602
R8990 VSS.n989 VSS.n988 1.76602
R8991 VSS.n975 VSS.n974 1.76602
R8992 VSS.n961 VSS.n960 1.76602
R8993 VSS.n1147 VSS.n1146 1.76602
R8994 VSS.n1133 VSS.n1132 1.76602
R8995 VSS.n1117 VSS.n1116 1.76602
R8996 VSS.n1103 VSS.n1102 1.76602
R8997 VSS.n1089 VSS.n1088 1.76602
R8998 VSS.n1075 VSS.n1074 1.76602
R8999 VSS.n1421 VSS.n1419 1.72554
R9000 VSS.n1436 VSS.n1434 1.72554
R9001 VSS.n1451 VSS.n1449 1.72554
R9002 VSS.n1466 VSS.n1464 1.72554
R9003 VSS.n1481 VSS.n1479 1.72554
R9004 VSS.n127 VSS.n125 1.72554
R9005 VSS.n150 VSS.n148 1.72554
R9006 VSS.n2101 VSS.n2099 1.72554
R9007 VSS.n3780 VSS.n3778 1.72554
R9008 VSS.n3666 VSS.n3664 1.72554
R9009 VSS.n3552 VSS.n3550 1.72554
R9010 VSS.n5 VSS.n3 1.72554
R9011 VSS.n4178 VSS.n4176 1.72554
R9012 VSS.n3360 VSS.n3357 1.67007
R9013 VSS.n3897 VSS.n3895 1.57241
R9014 VSS.n3921 VSS.n3919 1.57241
R9015 VSS.n1981 VSS.n1980 1.57241
R9016 VSS.n1416 VSS.n1414 1.57241
R9017 VSS.n1880 VSS.n1879 1.57241
R9018 VSS.n1431 VSS.n1429 1.57241
R9019 VSS.n1779 VSS.n1778 1.57241
R9020 VSS.n1446 VSS.n1444 1.57241
R9021 VSS.n1678 VSS.n1677 1.57241
R9022 VSS.n1461 VSS.n1459 1.57241
R9023 VSS.n1577 VSS.n1576 1.57241
R9024 VSS.n1476 VSS.n1474 1.57241
R9025 VSS.n3403 VSS.n3401 1.57241
R9026 VSS.n3427 VSS.n3425 1.57241
R9027 VSS.n132 VSS.n130 1.57241
R9028 VSS.n1233 VSS.n1231 1.57241
R9029 VSS.n1189 VSS.n1187 1.57241
R9030 VSS.n1999 VSS.n1997 1.57241
R9031 VSS.n2087 VSS.n2085 1.57241
R9032 VSS.n2114 VSS.n2112 1.57241
R9033 VSS.n4192 VSS.n4190 1.57241
R9034 VSS.n4278 VSS.n4277 1.57241
R9035 VSS.n3452 VSS.n3450 1.57241
R9036 VSS.n3540 VSS.n3539 1.57241
R9037 VSS.n3566 VSS.n3564 1.57241
R9038 VSS.n3654 VSS.n3653 1.57241
R9039 VSS.n3680 VSS.n3678 1.57241
R9040 VSS.n3768 VSS.n3767 1.57241
R9041 VSS.n3794 VSS.n3792 1.57241
R9042 VSS.n3882 VSS.n3880 1.57241
R9043 VSS.n2166 VSS.n2165 1.54533
R9044 VSS.n2175 VSS.n2174 1.54533
R9045 VSS.n2180 VSS.n2179 1.54533
R9046 VSS.n2189 VSS.n2188 1.54533
R9047 VSS.n2194 VSS.n2193 1.54533
R9048 VSS.n2203 VSS.n2202 1.54533
R9049 VSS.n2210 VSS.n2209 1.54533
R9050 VSS.n2219 VSS.n2218 1.54533
R9051 VSS.n2224 VSS.n2223 1.54533
R9052 VSS.n2233 VSS.n2232 1.54533
R9053 VSS.n2238 VSS.n2237 1.54533
R9054 VSS.n2247 VSS.n2246 1.54533
R9055 VSS.n2252 VSS.n2251 1.54533
R9056 VSS.n2261 VSS.n2260 1.54533
R9057 VSS.n2266 VSS.n2265 1.54533
R9058 VSS.n2275 VSS.n2274 1.54533
R9059 VSS.n2293 VSS.n2292 1.54533
R9060 VSS.n2302 VSS.n2301 1.54533
R9061 VSS.n2307 VSS.n2306 1.54533
R9062 VSS.n2316 VSS.n2315 1.54533
R9063 VSS.n2335 VSS.n2334 1.54533
R9064 VSS.n2345 VSS.n2344 1.54533
R9065 VSS.n2343 VSS.n120 1.54533
R9066 VSS.n2351 VSS.n121 1.54533
R9067 VSS.n2365 VSS.n2364 1.54533
R9068 VSS.n2374 VSS.n2373 1.54533
R9069 VSS.n2391 VSS.n2390 1.54533
R9070 VSS.n2400 VSS.n2399 1.54533
R9071 VSS.n2405 VSS.n2404 1.54533
R9072 VSS.n2414 VSS.n2413 1.54533
R9073 VSS.n2419 VSS.n2418 1.54533
R9074 VSS.n2428 VSS.n2427 1.54533
R9075 VSS.n2433 VSS.n2432 1.54533
R9076 VSS.n2443 VSS.n2442 1.54533
R9077 VSS.n2448 VSS.n2447 1.54533
R9078 VSS.n2457 VSS.n2456 1.54533
R9079 VSS.n2462 VSS.n2461 1.54533
R9080 VSS.n2471 VSS.n2470 1.54533
R9081 VSS.n2476 VSS.n2475 1.54533
R9082 VSS.n2485 VSS.n2484 1.54533
R9083 VSS.n2490 VSS.n2489 1.54533
R9084 VSS.n2500 VSS.n2499 1.54533
R9085 VSS.n2513 VSS.n2512 1.54533
R9086 VSS.n2518 VSS.n2517 1.54533
R9087 VSS.n2527 VSS.n2526 1.54533
R9088 VSS.n2532 VSS.n2531 1.54533
R9089 VSS.n2541 VSS.n2540 1.54533
R9090 VSS.n2546 VSS.n2545 1.54533
R9091 VSS.n2555 VSS.n2554 1.54533
R9092 VSS.n2562 VSS.n2561 1.54533
R9093 VSS.n2571 VSS.n2570 1.54533
R9094 VSS.n2576 VSS.n2575 1.54533
R9095 VSS.n2585 VSS.n2584 1.54533
R9096 VSS.n2590 VSS.n2589 1.54533
R9097 VSS.n2599 VSS.n2598 1.54533
R9098 VSS.n2604 VSS.n2603 1.54533
R9099 VSS.n2613 VSS.n2612 1.54533
R9100 VSS.n2618 VSS.n2617 1.54533
R9101 VSS.n2627 VSS.n2626 1.54533
R9102 VSS.n2645 VSS.n2644 1.54533
R9103 VSS.n2654 VSS.n2653 1.54533
R9104 VSS.n2659 VSS.n2658 1.54533
R9105 VSS.n2668 VSS.n2667 1.54533
R9106 VSS.n2687 VSS.n2686 1.54533
R9107 VSS.n2697 VSS.n2696 1.54533
R9108 VSS.n2695 VSS.n109 1.54533
R9109 VSS.n2703 VSS.n110 1.54533
R9110 VSS.n2717 VSS.n2716 1.54533
R9111 VSS.n2726 VSS.n2725 1.54533
R9112 VSS.n2743 VSS.n2742 1.54533
R9113 VSS.n2752 VSS.n2751 1.54533
R9114 VSS.n2757 VSS.n2756 1.54533
R9115 VSS.n2766 VSS.n2765 1.54533
R9116 VSS.n2771 VSS.n2770 1.54533
R9117 VSS.n2780 VSS.n2779 1.54533
R9118 VSS.n2785 VSS.n2784 1.54533
R9119 VSS.n2795 VSS.n2794 1.54533
R9120 VSS.n2800 VSS.n2799 1.54533
R9121 VSS.n2809 VSS.n2808 1.54533
R9122 VSS.n2814 VSS.n2813 1.54533
R9123 VSS.n2823 VSS.n2822 1.54533
R9124 VSS.n2828 VSS.n2827 1.54533
R9125 VSS.n2837 VSS.n2836 1.54533
R9126 VSS.n2842 VSS.n2841 1.54533
R9127 VSS.n2852 VSS.n2851 1.54533
R9128 VSS.n2865 VSS.n2864 1.54533
R9129 VSS.n2870 VSS.n2869 1.54533
R9130 VSS.n2879 VSS.n2878 1.54533
R9131 VSS.n2884 VSS.n2883 1.54533
R9132 VSS.n2893 VSS.n2892 1.54533
R9133 VSS.n2898 VSS.n2897 1.54533
R9134 VSS.n2907 VSS.n2906 1.54533
R9135 VSS.n2914 VSS.n2913 1.54533
R9136 VSS.n2923 VSS.n2922 1.54533
R9137 VSS.n2928 VSS.n2927 1.54533
R9138 VSS.n2937 VSS.n2936 1.54533
R9139 VSS.n2942 VSS.n2941 1.54533
R9140 VSS.n2951 VSS.n2950 1.54533
R9141 VSS.n2956 VSS.n2955 1.54533
R9142 VSS.n2965 VSS.n2964 1.54533
R9143 VSS.n2970 VSS.n2969 1.54533
R9144 VSS.n2979 VSS.n2978 1.54533
R9145 VSS.n2997 VSS.n2996 1.54533
R9146 VSS.n3006 VSS.n3005 1.54533
R9147 VSS.n3011 VSS.n3010 1.54533
R9148 VSS.n3020 VSS.n3019 1.54533
R9149 VSS.n92 VSS.n91 1.54533
R9150 VSS.n3041 VSS.n3040 1.54533
R9151 VSS.n3043 VSS.n3042 1.54533
R9152 VSS.n3053 VSS.n3052 1.54533
R9153 VSS.n3067 VSS.n3066 1.54533
R9154 VSS.n3072 VSS.n3071 1.54533
R9155 VSS.n3081 VSS.n3080 1.54533
R9156 VSS.n88 VSS.n87 1.54533
R9157 VSS.n3328 VSS.n89 1.54533
R9158 VSS.n3312 VSS.n3311 1.54533
R9159 VSS.n3323 VSS.n3322 1.54533
R9160 VSS.n3298 VSS.n3297 1.54533
R9161 VSS.n3307 VSS.n3306 1.54533
R9162 VSS.n3282 VSS.n3281 1.54533
R9163 VSS.n3293 VSS.n3292 1.54533
R9164 VSS.n3269 VSS.n3268 1.54533
R9165 VSS.n3277 VSS.n3276 1.54533
R9166 VSS.n3253 VSS.n3252 1.54533
R9167 VSS.n3264 VSS.n3263 1.54533
R9168 VSS.n3263 VSS.n3262 1.54533
R9169 VSS.n3239 VSS.n3238 1.54533
R9170 VSS.n3248 VSS.n3247 1.54533
R9171 VSS.n3224 VSS.n3223 1.54533
R9172 VSS.n3234 VSS.n3233 1.54533
R9173 VSS.n3209 VSS.n3208 1.54533
R9174 VSS.n3218 VSS.n3217 1.54533
R9175 VSS.n3194 VSS.n3193 1.54533
R9176 VSS.n3204 VSS.n3203 1.54533
R9177 VSS.n3179 VSS.n3178 1.54533
R9178 VSS.n3188 VSS.n3187 1.54533
R9179 VSS.n3164 VSS.n3163 1.54533
R9180 VSS.n3165 VSS.n3164 1.54533
R9181 VSS.n3174 VSS.n3173 1.54533
R9182 VSS.n3147 VSS.n3146 1.54533
R9183 VSS.n3158 VSS.n3157 1.54533
R9184 VSS.n3133 VSS.n3132 1.54533
R9185 VSS.n3142 VSS.n3141 1.54533
R9186 VSS.n3117 VSS.n3116 1.54533
R9187 VSS.n3128 VSS.n3127 1.54533
R9188 VSS.n3103 VSS.n3102 1.54533
R9189 VSS.n3112 VSS.n3111 1.54533
R9190 VSS.n3087 VSS.n3086 1.54533
R9191 VSS.n3098 VSS.n3097 1.54533
R9192 VSS.n69 VSS.n68 1.54533
R9193 VSS.n3383 VSS.n3382 1.54533
R9194 VSS.n66 VSS.n65 1.54533
R9195 VSS.n3389 VSS.n56 1.54533
R9196 VSS.n276 VSS.n275 1.54533
R9197 VSS.n299 VSS.n298 1.54533
R9198 VSS.n402 VSS.n401 1.54533
R9199 VSS.n388 VSS.n387 1.54533
R9200 VSS.n374 VSS.n373 1.54533
R9201 VSS.n360 VSS.n359 1.54533
R9202 VSS.n344 VSS.n343 1.54533
R9203 VSS.n330 VSS.n329 1.54533
R9204 VSS.n316 VSS.n315 1.54533
R9205 VSS.n544 VSS.n543 1.54533
R9206 VSS.n530 VSS.n529 1.54533
R9207 VSS.n516 VSS.n515 1.54533
R9208 VSS.n502 VSS.n501 1.54533
R9209 VSS.n486 VSS.n485 1.54533
R9210 VSS.n472 VSS.n471 1.54533
R9211 VSS.n458 VSS.n457 1.54533
R9212 VSS.n444 VSS.n443 1.54533
R9213 VSS.n430 VSS.n429 1.54533
R9214 VSS.n575 VSS.n574 1.54533
R9215 VSS.n561 VSS.n560 1.54533
R9216 VSS.n217 VSS.n216 1.54533
R9217 VSS.n607 VSS.n606 1.54533
R9218 VSS.n617 VSS.n616 1.54533
R9219 VSS.n720 VSS.n719 1.54533
R9220 VSS.n706 VSS.n705 1.54533
R9221 VSS.n692 VSS.n691 1.54533
R9222 VSS.n678 VSS.n677 1.54533
R9223 VSS.n662 VSS.n661 1.54533
R9224 VSS.n648 VSS.n647 1.54533
R9225 VSS.n634 VSS.n633 1.54533
R9226 VSS.n862 VSS.n861 1.54533
R9227 VSS.n848 VSS.n847 1.54533
R9228 VSS.n834 VSS.n833 1.54533
R9229 VSS.n820 VSS.n819 1.54533
R9230 VSS.n804 VSS.n803 1.54533
R9231 VSS.n790 VSS.n789 1.54533
R9232 VSS.n776 VSS.n775 1.54533
R9233 VSS.n762 VSS.n761 1.54533
R9234 VSS.n748 VSS.n747 1.54533
R9235 VSS.n893 VSS.n892 1.54533
R9236 VSS.n879 VSS.n878 1.54533
R9237 VSS.n172 VSS.n171 1.54533
R9238 VSS.n925 VSS.n924 1.54533
R9239 VSS.n935 VSS.n934 1.54533
R9240 VSS.n1038 VSS.n1037 1.54533
R9241 VSS.n1024 VSS.n1023 1.54533
R9242 VSS.n1010 VSS.n1009 1.54533
R9243 VSS.n996 VSS.n995 1.54533
R9244 VSS.n980 VSS.n979 1.54533
R9245 VSS.n966 VSS.n965 1.54533
R9246 VSS.n952 VSS.n951 1.54533
R9247 VSS.n1138 VSS.n1137 1.54533
R9248 VSS.n1122 VSS.n1121 1.54533
R9249 VSS.n1108 VSS.n1107 1.54533
R9250 VSS.n1094 VSS.n1093 1.54533
R9251 VSS.n1080 VSS.n1079 1.54533
R9252 VSS.n1066 VSS.n1065 1.54533
R9253 VSS.n1411 VSS.n1410 1.49652
R9254 VSS.n1426 VSS.n1425 1.49652
R9255 VSS.n1441 VSS.n1440 1.49652
R9256 VSS.n1456 VSS.n1455 1.49652
R9257 VSS.n1471 VSS.n1470 1.49652
R9258 VSS.n1253 VSS.n1252 1.49652
R9259 VSS.n2008 VSS.n2007 1.49652
R9260 VSS.n2123 VSS.n2122 1.49652
R9261 VSS.n4270 VSS.n4269 1.49652
R9262 VSS.n3530 VSS.n3529 1.49652
R9263 VSS.n3644 VSS.n3643 1.49652
R9264 VSS.n3758 VSS.n3757 1.49652
R9265 VSS.n3872 VSS.n3871 1.49652
R9266 VSS.n157 VSS.n154 1.48887
R9267 VSS.n202 VSS.n199 1.48887
R9268 VSS.n247 VSS.n244 1.48887
R9269 VSS.n167 VSS.n164 1.48827
R9270 VSS.n193 VSS.n190 1.48827
R9271 VSS.n212 VSS.n209 1.48827
R9272 VSS.n238 VSS.n235 1.48827
R9273 VSS.n257 VSS.n254 1.48827
R9274 VSS.n2328 VSS.n2325 1.48702
R9275 VSS.n2680 VSS.n2677 1.48702
R9276 VSS.n3032 VSS.n3029 1.48702
R9277 VSS.n1155 VSS.n1154 1.4204
R9278 VSS.n1154 VSS.n1153 1.4204
R9279 VSS.n1165 VSS.n1164 1.4204
R9280 VSS.n1164 VSS.n1163 1.4204
R9281 VSS.n1175 VSS.n1174 1.4204
R9282 VSS.n1174 VSS.n1173 1.4204
R9283 VSS.n1185 VSS.n1184 1.4204
R9284 VSS.n1196 VSS.n1195 1.4204
R9285 VSS.n1195 VSS.n1194 1.4204
R9286 VSS.n1206 VSS.n1205 1.4204
R9287 VSS.n1205 VSS.n1204 1.4204
R9288 VSS.n144 VSS.n143 1.4204
R9289 VSS.n1217 VSS.n1216 1.4204
R9290 VSS.n1218 VSS.n1217 1.4204
R9291 VSS.n138 VSS.n134 1.4204
R9292 VSS.n139 VSS.n138 1.4204
R9293 VSS.n1229 VSS.n1228 1.4204
R9294 VSS.n1240 VSS.n1239 1.4204
R9295 VSS.n1239 VSS.n1238 1.4204
R9296 VSS.n1250 VSS.n1249 1.4204
R9297 VSS.n1260 VSS.n1259 1.4204
R9298 VSS.n1259 VSS.n1258 1.4204
R9299 VSS.n1270 VSS.n1269 1.4204
R9300 VSS.n1269 VSS.n1268 1.4204
R9301 VSS.n1280 VSS.n1279 1.4204
R9302 VSS.n1279 VSS.n1278 1.4204
R9303 VSS.n1292 VSS.n1291 1.4204
R9304 VSS.n1291 VSS.n1290 1.4204
R9305 VSS.n1302 VSS.n1301 1.4204
R9306 VSS.n1301 VSS.n1300 1.4204
R9307 VSS.n1312 VSS.n1311 1.4204
R9308 VSS.n1311 VSS.n1310 1.4204
R9309 VSS.n1322 VSS.n1321 1.4204
R9310 VSS.n1321 VSS.n1320 1.4204
R9311 VSS.n1332 VSS.n1331 1.4204
R9312 VSS.n1331 VSS.n1330 1.4204
R9313 VSS.n1342 VSS.n1341 1.4204
R9314 VSS.n1341 VSS.n1340 1.4204
R9315 VSS.n1352 VSS.n1351 1.4204
R9316 VSS.n1351 VSS.n1350 1.4204
R9317 VSS.n1362 VSS.n1361 1.4204
R9318 VSS.n1361 VSS.n1360 1.4204
R9319 VSS.n3058 VSS.n3057 1.32464
R9320 VSS.n3390 VSS.n3389 1.32464
R9321 VSS.n2499 VSS.n2498 1.10395
R9322 VSS.n2851 VSS.n2850 1.10395
R9323 VSS.n272 VSS.n268 1.08219
R9324 VSS.n3065 VSS.n3058 0.883259
R9325 VSS.n3391 VSS.n3390 0.883259
R9326 VSS.n273 VSS.n272 0.821308
R9327 VSS.n265 VSS.n264 0.780988
R9328 VSS.n266 VSS.n265 0.723468
R9329 VSS.n2329 VSS.n2321 0.662569
R9330 VSS.n2681 VSS.n2673 0.662569
R9331 VSS.n3033 VSS.n3025 0.662569
R9332 VSS.n87 VSS.n86 0.662569
R9333 VSS.n3097 VSS.n3096 0.662569
R9334 VSS.n4163 VSS.n4162 0.662569
R9335 VSS.n4149 VSS.n4148 0.662569
R9336 VSS.n4135 VSS.n4134 0.662569
R9337 VSS.n4144 VSS.n4143 0.662569
R9338 VSS.n4122 VSS.n4121 0.662569
R9339 VSS.n4130 VSS.n4129 0.662569
R9340 VSS.n17 VSS.n16 0.662569
R9341 VSS.n25 VSS.n24 0.662569
R9342 VSS.n4114 VSS.n4113 0.662569
R9343 VSS.n4093 VSS.n4092 0.662569
R9344 VSS.n4102 VSS.n4101 0.662569
R9345 VSS.n4079 VSS.n4078 0.662569
R9346 VSS.n4088 VSS.n4087 0.662569
R9347 VSS.n4065 VSS.n4064 0.662569
R9348 VSS.n4074 VSS.n4073 0.662569
R9349 VSS.n29 VSS.n28 0.662569
R9350 VSS.n38 VSS.n37 0.662569
R9351 VSS.n4057 VSS.n4056 0.662569
R9352 VSS.n4036 VSS.n4035 0.662569
R9353 VSS.n4045 VSS.n4044 0.662569
R9354 VSS.n4022 VSS.n4021 0.662569
R9355 VSS.n4031 VSS.n4030 0.662569
R9356 VSS.n4008 VSS.n4007 0.662569
R9357 VSS.n4017 VSS.n4016 0.662569
R9358 VSS.n3993 VSS.n3992 0.662569
R9359 VSS.n4003 VSS.n4002 0.662569
R9360 VSS.n3979 VSS.n3978 0.662569
R9361 VSS.n3988 VSS.n3987 0.662569
R9362 VSS.n3964 VSS.n3963 0.662569
R9363 VSS.n3974 VSS.n3973 0.662569
R9364 VSS.n3950 VSS.n3949 0.662569
R9365 VSS.n3959 VSS.n3958 0.662569
R9366 VSS.n43 VSS.n42 0.662569
R9367 VSS.n423 VSS.n415 0.662569
R9368 VSS.n741 VSS.n733 0.662569
R9369 VSS.n1059 VSS.n1051 0.662569
R9370 VSS.n1332 VSS.n1327 0.662569
R9371 VSS.n3924 VSS 0.622896
R9372 VSS.n145 VSS.n144 0.577409
R9373 VSS.n1231 VSS.n1230 0.535538
R9374 VSS.n1187 VSS.n1186 0.535538
R9375 VSS.n1252 VSS.n1251 0.517621
R9376 VSS.n3234 VSS.n3232 0.441879
R9377 VSS.n3195 VSS.n3194 0.441879
R9378 VSS.n3945 VSS.n3944 0.441879
R9379 VSS.n1988 VSS.n1987 0.268864
R9380 VSS.n3396 VSS.n60 0.22119
R9381 VSS.n39 VSS.n38 0.22119
R9382 VSS.n3944 VSS.n3943 0.22119
R9383 VSS.n3927 VSS.n54 0.22119
R9384 VSS.n4173 VSS.n8 0.208232
R9385 VSS.n1988 VSS.n1407 0.188667
R9386 VSS.n3342 VSS.n3341 0.186007
R9387 VSS.n1990 VSS.n1989 0.182006
R9388 VSS.n263 VSS 0.156598
R9389 VSS.n2000 VSS.n1990 0.120292
R9390 VSS.n2004 VSS.n2000 0.120292
R9391 VSS.n2009 VSS.n2004 0.120292
R9392 VSS.n2013 VSS.n2009 0.120292
R9393 VSS.n2017 VSS.n2013 0.120292
R9394 VSS.n2021 VSS.n2017 0.120292
R9395 VSS.n2027 VSS.n2021 0.120292
R9396 VSS.n2031 VSS.n2027 0.120292
R9397 VSS.n2035 VSS.n2031 0.120292
R9398 VSS.n2039 VSS.n2035 0.120292
R9399 VSS.n2044 VSS.n2039 0.120292
R9400 VSS.n2048 VSS.n2044 0.120292
R9401 VSS.n2052 VSS.n2048 0.120292
R9402 VSS.n2056 VSS.n2052 0.120292
R9403 VSS.n2060 VSS.n2056 0.120292
R9404 VSS.n2066 VSS.n2060 0.120292
R9405 VSS.n2070 VSS.n2066 0.120292
R9406 VSS.n2074 VSS.n2070 0.120292
R9407 VSS.n2078 VSS.n2074 0.120292
R9408 VSS.n2082 VSS.n2078 0.120292
R9409 VSS.n2088 VSS.n2082 0.120292
R9410 VSS.n2092 VSS.n2088 0.120292
R9411 VSS.n2096 VSS.n2092 0.120292
R9412 VSS.n2102 VSS.n2096 0.120292
R9413 VSS.n2103 VSS.n2102 0.120292
R9414 VSS.n2115 VSS.n122 0.120292
R9415 VSS.n2119 VSS.n2115 0.120292
R9416 VSS.n2124 VSS.n2119 0.120292
R9417 VSS.n2128 VSS.n2124 0.120292
R9418 VSS.n2132 VSS.n2128 0.120292
R9419 VSS.n2136 VSS.n2132 0.120292
R9420 VSS.n2142 VSS.n2136 0.120292
R9421 VSS.n2146 VSS.n2142 0.120292
R9422 VSS.n2150 VSS.n2146 0.120292
R9423 VSS.n2154 VSS.n2150 0.120292
R9424 VSS.n2159 VSS.n2154 0.120292
R9425 VSS.n2163 VSS.n2159 0.120292
R9426 VSS.n3398 VSS.n3397 0.120292
R9427 VSS.n3404 VSS.n3398 0.120292
R9428 VSS.n3408 VSS.n3404 0.120292
R9429 VSS.n3414 VSS.n3408 0.120292
R9430 VSS.n3415 VSS.n3414 0.120292
R9431 VSS.n3428 VSS.n3422 0.120292
R9432 VSS.n3429 VSS.n3428 0.120292
R9433 VSS.n3924 VSS.n3923 0.120292
R9434 VSS.n3923 VSS.n3922 0.120292
R9435 VSS.n3922 VSS.n3916 0.120292
R9436 VSS.n3916 VSS.n3912 0.120292
R9437 VSS.n3912 VSS.n3906 0.120292
R9438 VSS.n3899 VSS.n3898 0.120292
R9439 VSS.n3898 VSS.n3892 0.120292
R9440 VSS.n1407 VSS.n1402 0.120292
R9441 VSS.n1402 VSS.n1401 0.120292
R9442 VSS.n1401 VSS.n1397 0.120292
R9443 VSS.n1397 VSS.n1393 0.120292
R9444 VSS.n1393 VSS.n1392 0.120292
R9445 VSS.n1392 VSS.n1388 0.120292
R9446 VSS.n1388 VSS.n1384 0.120292
R9447 VSS.n1384 VSS.n1380 0.120292
R9448 VSS.n1380 VSS.n1376 0.120292
R9449 VSS.n1376 VSS.n1370 0.120292
R9450 VSS.n1370 VSS.n1366 0.120292
R9451 VSS.n1366 VSS.n1356 0.120292
R9452 VSS.n1356 VSS.n1346 0.120292
R9453 VSS.n1346 VSS.n1336 0.120292
R9454 VSS.n1336 VSS.n1326 0.120292
R9455 VSS.n1326 VSS.n1316 0.120292
R9456 VSS.n1316 VSS.n1306 0.120292
R9457 VSS.n1306 VSS.n1296 0.120292
R9458 VSS.n1296 VSS.n1284 0.120292
R9459 VSS.n1284 VSS.n1274 0.120292
R9460 VSS.n1274 VSS.n1264 0.120292
R9461 VSS.n1264 VSS.n1254 0.120292
R9462 VSS.n1254 VSS.n1244 0.120292
R9463 VSS.n1244 VSS.n1234 0.120292
R9464 VSS.n1234 VSS.n1223 0.120292
R9465 VSS.n1212 VSS.n1211 0.120292
R9466 VSS.n1211 VSS.n1210 0.120292
R9467 VSS.n1210 VSS.n1200 0.120292
R9468 VSS.n1200 VSS.n1190 0.120292
R9469 VSS.n1190 VSS.n1179 0.120292
R9470 VSS.n1179 VSS.n1169 0.120292
R9471 VSS.n1169 VSS.n1159 0.120292
R9472 VSS.n278 VSS.n80 0.120292
R9473 VSS.n3337 VSS.n80 0.120292
R9474 VSS.n1978 VSS.n1977 0.120292
R9475 VSS.n1977 VSS.n1973 0.120292
R9476 VSS.n1973 VSS.n1972 0.120292
R9477 VSS.n1972 VSS.n1968 0.120292
R9478 VSS.n1968 VSS.n1964 0.120292
R9479 VSS.n1964 VSS.n1960 0.120292
R9480 VSS.n1960 VSS.n1954 0.120292
R9481 VSS.n1954 VSS.n1950 0.120292
R9482 VSS.n1950 VSS.n1946 0.120292
R9483 VSS.n1946 VSS.n1942 0.120292
R9484 VSS.n1942 VSS.n1937 0.120292
R9485 VSS.n1937 VSS.n1933 0.120292
R9486 VSS.n1933 VSS.n1929 0.120292
R9487 VSS.n1929 VSS.n1925 0.120292
R9488 VSS.n1925 VSS.n1921 0.120292
R9489 VSS.n1921 VSS.n1915 0.120292
R9490 VSS.n1915 VSS.n1911 0.120292
R9491 VSS.n1911 VSS.n1907 0.120292
R9492 VSS.n1907 VSS.n1903 0.120292
R9493 VSS.n1903 VSS.n1899 0.120292
R9494 VSS.n1899 VSS.n1898 0.120292
R9495 VSS.n1898 VSS.n1894 0.120292
R9496 VSS.n1894 VSS.n1890 0.120292
R9497 VSS.n1890 VSS.n1889 0.120292
R9498 VSS.n1877 VSS.n1876 0.120292
R9499 VSS.n1876 VSS.n1872 0.120292
R9500 VSS.n1872 VSS.n1871 0.120292
R9501 VSS.n1871 VSS.n1867 0.120292
R9502 VSS.n1867 VSS.n1863 0.120292
R9503 VSS.n1863 VSS.n1859 0.120292
R9504 VSS.n1859 VSS.n1853 0.120292
R9505 VSS.n1853 VSS.n1849 0.120292
R9506 VSS.n1849 VSS.n1845 0.120292
R9507 VSS.n1845 VSS.n1841 0.120292
R9508 VSS.n1841 VSS.n1836 0.120292
R9509 VSS.n1836 VSS.n1832 0.120292
R9510 VSS.n1832 VSS.n1828 0.120292
R9511 VSS.n1828 VSS.n1824 0.120292
R9512 VSS.n1824 VSS.n1820 0.120292
R9513 VSS.n1820 VSS.n1814 0.120292
R9514 VSS.n1814 VSS.n1810 0.120292
R9515 VSS.n1810 VSS.n1806 0.120292
R9516 VSS.n1806 VSS.n1802 0.120292
R9517 VSS.n1802 VSS.n1798 0.120292
R9518 VSS.n1798 VSS.n1797 0.120292
R9519 VSS.n1797 VSS.n1793 0.120292
R9520 VSS.n1793 VSS.n1789 0.120292
R9521 VSS.n1789 VSS.n1788 0.120292
R9522 VSS.n1776 VSS.n1775 0.120292
R9523 VSS.n1775 VSS.n1771 0.120292
R9524 VSS.n1771 VSS.n1770 0.120292
R9525 VSS.n1770 VSS.n1766 0.120292
R9526 VSS.n1766 VSS.n1762 0.120292
R9527 VSS.n1762 VSS.n1758 0.120292
R9528 VSS.n1758 VSS.n1752 0.120292
R9529 VSS.n1752 VSS.n1748 0.120292
R9530 VSS.n1748 VSS.n1744 0.120292
R9531 VSS.n1744 VSS.n1740 0.120292
R9532 VSS.n1740 VSS.n1735 0.120292
R9533 VSS.n1735 VSS.n1731 0.120292
R9534 VSS.n1731 VSS.n1727 0.120292
R9535 VSS.n1727 VSS.n1723 0.120292
R9536 VSS.n1723 VSS.n1719 0.120292
R9537 VSS.n1719 VSS.n1713 0.120292
R9538 VSS.n1713 VSS.n1709 0.120292
R9539 VSS.n1709 VSS.n1705 0.120292
R9540 VSS.n1705 VSS.n1701 0.120292
R9541 VSS.n1701 VSS.n1697 0.120292
R9542 VSS.n1697 VSS.n1696 0.120292
R9543 VSS.n1696 VSS.n1692 0.120292
R9544 VSS.n1692 VSS.n1688 0.120292
R9545 VSS.n1688 VSS.n1687 0.120292
R9546 VSS.n1675 VSS.n1674 0.120292
R9547 VSS.n1674 VSS.n1670 0.120292
R9548 VSS.n1670 VSS.n1669 0.120292
R9549 VSS.n1669 VSS.n1665 0.120292
R9550 VSS.n1665 VSS.n1661 0.120292
R9551 VSS.n1661 VSS.n1657 0.120292
R9552 VSS.n1657 VSS.n1651 0.120292
R9553 VSS.n1651 VSS.n1647 0.120292
R9554 VSS.n1647 VSS.n1643 0.120292
R9555 VSS.n1643 VSS.n1639 0.120292
R9556 VSS.n1639 VSS.n1634 0.120292
R9557 VSS.n1634 VSS.n1630 0.120292
R9558 VSS.n1630 VSS.n1626 0.120292
R9559 VSS.n1626 VSS.n1622 0.120292
R9560 VSS.n1622 VSS.n1618 0.120292
R9561 VSS.n1618 VSS.n1612 0.120292
R9562 VSS.n1612 VSS.n1608 0.120292
R9563 VSS.n1608 VSS.n1604 0.120292
R9564 VSS.n1604 VSS.n1600 0.120292
R9565 VSS.n1600 VSS.n1596 0.120292
R9566 VSS.n1596 VSS.n1595 0.120292
R9567 VSS.n1595 VSS.n1591 0.120292
R9568 VSS.n1591 VSS.n1587 0.120292
R9569 VSS.n1587 VSS.n1586 0.120292
R9570 VSS.n1574 VSS.n1573 0.120292
R9571 VSS.n1573 VSS.n1569 0.120292
R9572 VSS.n1569 VSS.n1568 0.120292
R9573 VSS.n1568 VSS.n1564 0.120292
R9574 VSS.n1564 VSS.n1560 0.120292
R9575 VSS.n1560 VSS.n1556 0.120292
R9576 VSS.n1556 VSS.n1550 0.120292
R9577 VSS.n1550 VSS.n1546 0.120292
R9578 VSS.n1546 VSS.n1542 0.120292
R9579 VSS.n1542 VSS.n1538 0.120292
R9580 VSS.n1538 VSS.n1533 0.120292
R9581 VSS.n1533 VSS.n1529 0.120292
R9582 VSS.n1529 VSS.n1525 0.120292
R9583 VSS.n1525 VSS.n1521 0.120292
R9584 VSS.n1521 VSS.n1517 0.120292
R9585 VSS.n1517 VSS.n1511 0.120292
R9586 VSS.n1511 VSS.n1507 0.120292
R9587 VSS.n1507 VSS.n1503 0.120292
R9588 VSS.n1503 VSS.n1499 0.120292
R9589 VSS.n1499 VSS.n1495 0.120292
R9590 VSS.n1495 VSS.n1494 0.120292
R9591 VSS.n1494 VSS.n1490 0.120292
R9592 VSS.n1490 VSS.n1486 0.120292
R9593 VSS.n1486 VSS.n1485 0.120292
R9594 VSS.n4179 VSS.n4173 0.120292
R9595 VSS.n4183 VSS.n4179 0.120292
R9596 VSS.n4187 VSS.n4183 0.120292
R9597 VSS.n4193 VSS.n4187 0.120292
R9598 VSS.n4197 VSS.n4193 0.120292
R9599 VSS.n4201 VSS.n4197 0.120292
R9600 VSS.n4205 VSS.n4201 0.120292
R9601 VSS.n4209 VSS.n4205 0.120292
R9602 VSS.n4215 VSS.n4209 0.120292
R9603 VSS.n4219 VSS.n4215 0.120292
R9604 VSS.n4223 VSS.n4219 0.120292
R9605 VSS.n4227 VSS.n4223 0.120292
R9606 VSS.n4231 VSS.n4227 0.120292
R9607 VSS.n4236 VSS.n4231 0.120292
R9608 VSS.n4240 VSS.n4236 0.120292
R9609 VSS.n4244 VSS.n4240 0.120292
R9610 VSS.n4248 VSS.n4244 0.120292
R9611 VSS.n4254 VSS.n4248 0.120292
R9612 VSS.n4258 VSS.n4254 0.120292
R9613 VSS.n4262 VSS.n4258 0.120292
R9614 VSS.n4266 VSS.n4262 0.120292
R9615 VSS.n4271 VSS.n4266 0.120292
R9616 VSS.n4275 VSS.n4271 0.120292
R9617 VSS.n4276 VSS.n4275 0.120292
R9618 VSS.n4276 VSS.n0 0.120292
R9619 VSS.n4287 VSS.n6 0.120292
R9620 VSS.n3443 VSS.n6 0.120292
R9621 VSS.n3447 VSS.n3443 0.120292
R9622 VSS.n3453 VSS.n3447 0.120292
R9623 VSS.n3457 VSS.n3453 0.120292
R9624 VSS.n3461 VSS.n3457 0.120292
R9625 VSS.n3465 VSS.n3461 0.120292
R9626 VSS.n3469 VSS.n3465 0.120292
R9627 VSS.n3475 VSS.n3469 0.120292
R9628 VSS.n3479 VSS.n3475 0.120292
R9629 VSS.n3483 VSS.n3479 0.120292
R9630 VSS.n3487 VSS.n3483 0.120292
R9631 VSS.n3491 VSS.n3487 0.120292
R9632 VSS.n3496 VSS.n3491 0.120292
R9633 VSS.n3500 VSS.n3496 0.120292
R9634 VSS.n3504 VSS.n3500 0.120292
R9635 VSS.n3508 VSS.n3504 0.120292
R9636 VSS.n3514 VSS.n3508 0.120292
R9637 VSS.n3518 VSS.n3514 0.120292
R9638 VSS.n3522 VSS.n3518 0.120292
R9639 VSS.n3526 VSS.n3522 0.120292
R9640 VSS.n3531 VSS.n3526 0.120292
R9641 VSS.n3535 VSS.n3531 0.120292
R9642 VSS.n3538 VSS.n3535 0.120292
R9643 VSS.n3538 VSS.n3537 0.120292
R9644 VSS.n3553 VSS.n3547 0.120292
R9645 VSS.n3557 VSS.n3553 0.120292
R9646 VSS.n3561 VSS.n3557 0.120292
R9647 VSS.n3567 VSS.n3561 0.120292
R9648 VSS.n3571 VSS.n3567 0.120292
R9649 VSS.n3575 VSS.n3571 0.120292
R9650 VSS.n3579 VSS.n3575 0.120292
R9651 VSS.n3583 VSS.n3579 0.120292
R9652 VSS.n3589 VSS.n3583 0.120292
R9653 VSS.n3593 VSS.n3589 0.120292
R9654 VSS.n3597 VSS.n3593 0.120292
R9655 VSS.n3601 VSS.n3597 0.120292
R9656 VSS.n3605 VSS.n3601 0.120292
R9657 VSS.n3610 VSS.n3605 0.120292
R9658 VSS.n3614 VSS.n3610 0.120292
R9659 VSS.n3618 VSS.n3614 0.120292
R9660 VSS.n3622 VSS.n3618 0.120292
R9661 VSS.n3628 VSS.n3622 0.120292
R9662 VSS.n3632 VSS.n3628 0.120292
R9663 VSS.n3636 VSS.n3632 0.120292
R9664 VSS.n3640 VSS.n3636 0.120292
R9665 VSS.n3645 VSS.n3640 0.120292
R9666 VSS.n3649 VSS.n3645 0.120292
R9667 VSS.n3652 VSS.n3649 0.120292
R9668 VSS.n3652 VSS.n3651 0.120292
R9669 VSS.n3667 VSS.n3661 0.120292
R9670 VSS.n3671 VSS.n3667 0.120292
R9671 VSS.n3675 VSS.n3671 0.120292
R9672 VSS.n3681 VSS.n3675 0.120292
R9673 VSS.n3685 VSS.n3681 0.120292
R9674 VSS.n3689 VSS.n3685 0.120292
R9675 VSS.n3693 VSS.n3689 0.120292
R9676 VSS.n3697 VSS.n3693 0.120292
R9677 VSS.n3703 VSS.n3697 0.120292
R9678 VSS.n3707 VSS.n3703 0.120292
R9679 VSS.n3711 VSS.n3707 0.120292
R9680 VSS.n3715 VSS.n3711 0.120292
R9681 VSS.n3719 VSS.n3715 0.120292
R9682 VSS.n3724 VSS.n3719 0.120292
R9683 VSS.n3728 VSS.n3724 0.120292
R9684 VSS.n3732 VSS.n3728 0.120292
R9685 VSS.n3736 VSS.n3732 0.120292
R9686 VSS.n3742 VSS.n3736 0.120292
R9687 VSS.n3746 VSS.n3742 0.120292
R9688 VSS.n3750 VSS.n3746 0.120292
R9689 VSS.n3754 VSS.n3750 0.120292
R9690 VSS.n3759 VSS.n3754 0.120292
R9691 VSS.n3763 VSS.n3759 0.120292
R9692 VSS.n3766 VSS.n3763 0.120292
R9693 VSS.n3766 VSS.n3765 0.120292
R9694 VSS.n3781 VSS.n3775 0.120292
R9695 VSS.n3785 VSS.n3781 0.120292
R9696 VSS.n3789 VSS.n3785 0.120292
R9697 VSS.n3795 VSS.n3789 0.120292
R9698 VSS.n3799 VSS.n3795 0.120292
R9699 VSS.n3803 VSS.n3799 0.120292
R9700 VSS.n3807 VSS.n3803 0.120292
R9701 VSS.n3811 VSS.n3807 0.120292
R9702 VSS.n3817 VSS.n3811 0.120292
R9703 VSS.n3821 VSS.n3817 0.120292
R9704 VSS.n3825 VSS.n3821 0.120292
R9705 VSS.n3829 VSS.n3825 0.120292
R9706 VSS.n3833 VSS.n3829 0.120292
R9707 VSS.n3838 VSS.n3833 0.120292
R9708 VSS.n3842 VSS.n3838 0.120292
R9709 VSS.n3846 VSS.n3842 0.120292
R9710 VSS.n3850 VSS.n3846 0.120292
R9711 VSS.n3856 VSS.n3850 0.120292
R9712 VSS.n3860 VSS.n3856 0.120292
R9713 VSS.n3864 VSS.n3860 0.120292
R9714 VSS.n3868 VSS.n3864 0.120292
R9715 VSS.n3873 VSS.n3868 0.120292
R9716 VSS.n3877 VSS.n3873 0.120292
R9717 VSS.n3883 VSS.n3877 0.120292
R9718 VSS.n3884 VSS.n3883 0.120292
R9719 VSS.n3374 VSS.n3373 0.119057
R9720 VSS.n3373 VSS.n3371 0.119057
R9721 VSS.n3371 VSS.n3365 0.119057
R9722 VSS.n3365 VSS.n3361 0.119057
R9723 VSS.n3361 VSS.n3355 0.119057
R9724 VSS.n3347 VSS.n3346 0.119057
R9725 VSS.n3346 VSS.n3343 0.119057
R9726 VSS.n1159 VSS.n1149 0.108573
R9727 VSS.n2164 VSS.n2163 0.107271
R9728 VSS.n2178 VSS.n2177 0.0981562
R9729 VSS.n2192 VSS.n2191 0.0981562
R9730 VSS.n2206 VSS.n2205 0.0981562
R9731 VSS.n2222 VSS.n2221 0.0981562
R9732 VSS.n2236 VSS.n2235 0.0981562
R9733 VSS.n2250 VSS.n2249 0.0981562
R9734 VSS.n2264 VSS.n2263 0.0981562
R9735 VSS.n2278 VSS.n2277 0.0981562
R9736 VSS.n2291 VSS.n2290 0.0981562
R9737 VSS.n2305 VSS.n2304 0.0981562
R9738 VSS.n2319 VSS.n2318 0.0981562
R9739 VSS.n2333 VSS.n2332 0.0981562
R9740 VSS.n2349 VSS.n111 0.0981562
R9741 VSS.n2363 VSS.n2362 0.0981562
R9742 VSS.n2377 VSS.n2376 0.0981562
R9743 VSS.n2389 VSS.n2388 0.0981562
R9744 VSS.n2403 VSS.n2402 0.0981562
R9745 VSS.n2417 VSS.n2416 0.0981562
R9746 VSS.n2431 VSS.n2430 0.0981562
R9747 VSS.n2446 VSS.n2445 0.0981562
R9748 VSS.n2460 VSS.n2459 0.0981562
R9749 VSS.n2474 VSS.n2473 0.0981562
R9750 VSS.n2488 VSS.n2487 0.0981562
R9751 VSS.n2503 VSS.n2502 0.0981562
R9752 VSS.n2516 VSS.n2515 0.0981562
R9753 VSS.n2530 VSS.n2529 0.0981562
R9754 VSS.n2544 VSS.n2543 0.0981562
R9755 VSS.n2558 VSS.n2557 0.0981562
R9756 VSS.n2574 VSS.n2573 0.0981562
R9757 VSS.n2588 VSS.n2587 0.0981562
R9758 VSS.n2602 VSS.n2601 0.0981562
R9759 VSS.n2616 VSS.n2615 0.0981562
R9760 VSS.n2630 VSS.n2629 0.0981562
R9761 VSS.n2643 VSS.n2642 0.0981562
R9762 VSS.n2657 VSS.n2656 0.0981562
R9763 VSS.n2671 VSS.n2670 0.0981562
R9764 VSS.n2685 VSS.n2684 0.0981562
R9765 VSS.n2701 VSS.n100 0.0981562
R9766 VSS.n2715 VSS.n2714 0.0981562
R9767 VSS.n2729 VSS.n2728 0.0981562
R9768 VSS.n2741 VSS.n2740 0.0981562
R9769 VSS.n2755 VSS.n2754 0.0981562
R9770 VSS.n2769 VSS.n2768 0.0981562
R9771 VSS.n2783 VSS.n2782 0.0981562
R9772 VSS.n2798 VSS.n2797 0.0981562
R9773 VSS.n2812 VSS.n2811 0.0981562
R9774 VSS.n2826 VSS.n2825 0.0981562
R9775 VSS.n2840 VSS.n2839 0.0981562
R9776 VSS.n2855 VSS.n2854 0.0981562
R9777 VSS.n2868 VSS.n2867 0.0981562
R9778 VSS.n2882 VSS.n2881 0.0981562
R9779 VSS.n2896 VSS.n2895 0.0981562
R9780 VSS.n2910 VSS.n2909 0.0981562
R9781 VSS.n2926 VSS.n2925 0.0981562
R9782 VSS.n2940 VSS.n2939 0.0981562
R9783 VSS.n2954 VSS.n2953 0.0981562
R9784 VSS.n2968 VSS.n2967 0.0981562
R9785 VSS.n2982 VSS.n2981 0.0981562
R9786 VSS.n2995 VSS.n2994 0.0981562
R9787 VSS.n3009 VSS.n3008 0.0981562
R9788 VSS.n3023 VSS.n3022 0.0981562
R9789 VSS.n3037 VSS.n3036 0.0981562
R9790 VSS.n3056 VSS.n3055 0.0981562
R9791 VSS.n3070 VSS.n3069 0.0981562
R9792 VSS.n3084 VSS.n3083 0.0981562
R9793 VSS.n3326 VSS.n3325 0.0981562
R9794 VSS.n3310 VSS.n3309 0.0981562
R9795 VSS.n3296 VSS.n3295 0.0981562
R9796 VSS.n3280 VSS.n3279 0.0981562
R9797 VSS.n3267 VSS.n3266 0.0981562
R9798 VSS.n3251 VSS.n3250 0.0981562
R9799 VSS.n3237 VSS.n3236 0.0981562
R9800 VSS.n3221 VSS.n3220 0.0981562
R9801 VSS.n3207 VSS.n3206 0.0981562
R9802 VSS.n3191 VSS.n3190 0.0981562
R9803 VSS.n3177 VSS.n3176 0.0981562
R9804 VSS.n3161 VSS.n3160 0.0981562
R9805 VSS.n3145 VSS.n3144 0.0981562
R9806 VSS.n3131 VSS.n3130 0.0981562
R9807 VSS.n3115 VSS.n3114 0.0981562
R9808 VSS.n3101 VSS.n3100 0.0981562
R9809 VSS.n3085 VSS.n67 0.0981562
R9810 VSS.n3386 VSS.n3385 0.0981562
R9811 VSS.n4152 VSS.n4151 0.0981562
R9812 VSS.n4147 VSS.n4146 0.0981562
R9813 VSS.n4133 VSS.n4132 0.0981562
R9814 VSS.n4120 VSS.n4119 0.0981562
R9815 VSS.n4117 VSS.n4116 0.0981562
R9816 VSS.n4105 VSS.n4104 0.0981562
R9817 VSS.n4091 VSS.n4090 0.0981562
R9818 VSS.n4077 VSS.n4076 0.0981562
R9819 VSS.n4063 VSS.n4062 0.0981562
R9820 VSS.n4060 VSS.n4059 0.0981562
R9821 VSS.n4048 VSS.n4047 0.0981562
R9822 VSS.n4034 VSS.n4033 0.0981562
R9823 VSS.n4020 VSS.n4019 0.0981562
R9824 VSS.n4006 VSS.n4005 0.0981562
R9825 VSS.n3991 VSS.n3990 0.0981562
R9826 VSS.n3977 VSS.n3976 0.0981562
R9827 VSS.n3962 VSS.n3961 0.0981562
R9828 VSS.n3948 VSS.n3947 0.0981562
R9829 VSS.n1136 VSS.n1135 0.0981562
R9830 VSS.n1120 VSS.n1119 0.0981562
R9831 VSS.n1106 VSS.n1105 0.0981562
R9832 VSS.n1092 VSS.n1091 0.0981562
R9833 VSS.n1078 VSS.n1077 0.0981562
R9834 VSS.n1064 VSS.n1063 0.0981562
R9835 VSS.n1050 VSS.n1049 0.0981562
R9836 VSS.n1036 VSS.n1035 0.0981562
R9837 VSS.n1022 VSS.n1021 0.0981562
R9838 VSS.n1008 VSS.n1007 0.0981562
R9839 VSS.n992 VSS.n991 0.0981562
R9840 VSS.n978 VSS.n977 0.0981562
R9841 VSS.n964 VSS.n963 0.0981562
R9842 VSS.n950 VSS.n949 0.0981562
R9843 VSS.n947 VSS.n946 0.0981562
R9844 VSS.n933 VSS.n932 0.0981562
R9845 VSS.n930 VSS.n929 0.0981562
R9846 VSS.n908 VSS.n907 0.0981562
R9847 VSS.n905 VSS.n904 0.0981562
R9848 VSS.n891 VSS.n890 0.0981562
R9849 VSS.n877 VSS.n876 0.0981562
R9850 VSS.n874 VSS.n873 0.0981562
R9851 VSS.n860 VSS.n859 0.0981562
R9852 VSS.n846 VSS.n845 0.0981562
R9853 VSS.n832 VSS.n831 0.0981562
R9854 VSS.n818 VSS.n817 0.0981562
R9855 VSS.n802 VSS.n801 0.0981562
R9856 VSS.n788 VSS.n787 0.0981562
R9857 VSS.n774 VSS.n773 0.0981562
R9858 VSS.n760 VSS.n759 0.0981562
R9859 VSS.n746 VSS.n745 0.0981562
R9860 VSS.n732 VSS.n731 0.0981562
R9861 VSS.n718 VSS.n717 0.0981562
R9862 VSS.n704 VSS.n703 0.0981562
R9863 VSS.n690 VSS.n689 0.0981562
R9864 VSS.n674 VSS.n673 0.0981562
R9865 VSS.n660 VSS.n659 0.0981562
R9866 VSS.n646 VSS.n645 0.0981562
R9867 VSS.n632 VSS.n631 0.0981562
R9868 VSS.n629 VSS.n628 0.0981562
R9869 VSS.n615 VSS.n614 0.0981562
R9870 VSS.n612 VSS.n611 0.0981562
R9871 VSS.n590 VSS.n589 0.0981562
R9872 VSS.n587 VSS.n586 0.0981562
R9873 VSS.n573 VSS.n572 0.0981562
R9874 VSS.n559 VSS.n558 0.0981562
R9875 VSS.n556 VSS.n555 0.0981562
R9876 VSS.n542 VSS.n541 0.0981562
R9877 VSS.n528 VSS.n527 0.0981562
R9878 VSS.n514 VSS.n513 0.0981562
R9879 VSS.n500 VSS.n499 0.0981562
R9880 VSS.n484 VSS.n483 0.0981562
R9881 VSS.n470 VSS.n469 0.0981562
R9882 VSS.n456 VSS.n455 0.0981562
R9883 VSS.n442 VSS.n441 0.0981562
R9884 VSS.n428 VSS.n427 0.0981562
R9885 VSS.n414 VSS.n413 0.0981562
R9886 VSS.n400 VSS.n399 0.0981562
R9887 VSS.n386 VSS.n385 0.0981562
R9888 VSS.n372 VSS.n371 0.0981562
R9889 VSS.n356 VSS.n355 0.0981562
R9890 VSS.n342 VSS.n341 0.0981562
R9891 VSS.n328 VSS.n327 0.0981562
R9892 VSS.n314 VSS.n313 0.0981562
R9893 VSS.n311 VSS.n310 0.0981562
R9894 VSS.n297 VSS.n296 0.0981562
R9895 VSS.n293 VSS.n292 0.0981562
R9896 VSS.n1978 VSS 0.0968542
R9897 VSS.n1877 VSS 0.0968542
R9898 VSS.n1776 VSS 0.0968542
R9899 VSS.n1675 VSS 0.0968542
R9900 VSS.n1574 VSS 0.0968542
R9901 VSS.n1989 VSS.n1988 0.0852709
R9902 VSS.n14 VSS 0.078625
R9903 VSS.n1989 VSS.n8 0.0637239
R9904 VSS.n2103 VSS 0.0603958
R9905 VSS VSS.n122 0.0603958
R9906 VSS.n3415 VSS 0.0603958
R9907 VSS.n3422 VSS 0.0603958
R9908 VSS.n3429 VSS 0.0603958
R9909 VSS.n3906 VSS 0.0603958
R9910 VSS.n3899 VSS 0.0603958
R9911 VSS.n3892 VSS 0.0603958
R9912 VSS.n1223 VSS 0.0603958
R9913 VSS.n1212 VSS 0.0603958
R9914 VSS.n1889 VSS 0.0603958
R9915 VSS.n1422 VSS 0.0603958
R9916 VSS.n1788 VSS 0.0603958
R9917 VSS.n1437 VSS 0.0603958
R9918 VSS.n1687 VSS 0.0603958
R9919 VSS.n1452 VSS 0.0603958
R9920 VSS.n1586 VSS 0.0603958
R9921 VSS.n1467 VSS 0.0603958
R9922 VSS.n1485 VSS 0.0603958
R9923 VSS VSS.n0 0.0603958
R9924 VSS VSS.n4287 0.0603958
R9925 VSS.n3537 VSS 0.0603958
R9926 VSS.n3547 VSS 0.0603958
R9927 VSS.n3651 VSS 0.0603958
R9928 VSS.n3661 VSS 0.0603958
R9929 VSS.n3765 VSS 0.0603958
R9930 VSS.n3775 VSS 0.0603958
R9931 VSS.n3884 VSS 0.0603958
R9932 VSS.n3355 VSS 0.0597784
R9933 VSS.n3347 VSS 0.0597784
R9934 VSS.n3343 VSS 0.0597784
R9935 VSS VSS.n41 0.0564896
R9936 VSS.n11 VSS.n8 0.0537635
R9937 VSS VSS.n2347 0.0512812
R9938 VSS VSS.n2699 0.0512812
R9939 VSS.n3038 VSS 0.0512812
R9940 VSS VSS.n170 0.0499792
R9941 VSS VSS.n215 0.0499792
R9942 VSS VSS.n274 0.0499792
R9943 VSS.n175 VSS 0.0486771
R9944 VSS.n220 VSS 0.0486771
R9945 VSS.n2348 VSS 0.047375
R9946 VSS.n2700 VSS 0.047375
R9947 VSS VSS.n90 0.047375
R9948 VSS.n278 VSS 0.0356562
R9949 VSS.n3397 VSS 0.0343542
R9950 VSS VSS.n12 0.0239375
R9951 VSS.n1987 VSS 0.0239375
R9952 VSS VSS.n1422 0.0239375
R9953 VSS VSS.n1437 0.0239375
R9954 VSS VSS.n1452 0.0239375
R9955 VSS VSS.n1467 0.0239375
R9956 VSS VSS.n3337 0.0226354
R9957 VSS.n4153 VSS.n14 0.0187292
R9958 VSS.n4151 VSS.n4150 0.0187292
R9959 VSS.n4146 VSS.n4145 0.0187292
R9960 VSS.n4132 VSS.n4131 0.0187292
R9961 VSS.n4119 VSS.n4118 0.0187292
R9962 VSS.n4116 VSS.n4115 0.0187292
R9963 VSS.n4104 VSS.n4103 0.0187292
R9964 VSS.n4090 VSS.n4089 0.0187292
R9965 VSS.n4076 VSS.n4075 0.0187292
R9966 VSS.n4062 VSS.n4061 0.0187292
R9967 VSS.n4059 VSS.n4058 0.0187292
R9968 VSS.n4047 VSS.n4046 0.0187292
R9969 VSS.n4033 VSS.n4032 0.0187292
R9970 VSS.n4019 VSS.n4018 0.0187292
R9971 VSS.n4005 VSS.n4004 0.0187292
R9972 VSS.n3990 VSS.n3989 0.0187292
R9973 VSS.n3976 VSS.n3975 0.0187292
R9974 VSS.n3961 VSS.n3960 0.0187292
R9975 VSS.n3947 VSS.n3946 0.0187292
R9976 VSS.n2176 VSS.n2164 0.0135208
R9977 VSS.n2190 VSS.n2178 0.0135208
R9978 VSS.n2204 VSS.n2192 0.0135208
R9979 VSS.n2220 VSS.n2206 0.0135208
R9980 VSS.n2234 VSS.n2222 0.0135208
R9981 VSS.n2248 VSS.n2236 0.0135208
R9982 VSS.n2262 VSS.n2250 0.0135208
R9983 VSS.n2276 VSS.n2264 0.0135208
R9984 VSS.n2289 VSS.n2278 0.0135208
R9985 VSS.n2303 VSS.n2291 0.0135208
R9986 VSS.n2317 VSS.n2305 0.0135208
R9987 VSS.n2331 VSS.n2319 0.0135208
R9988 VSS.n2346 VSS.n2333 0.0135208
R9989 VSS.n2350 VSS.n2348 0.0135208
R9990 VSS.n2361 VSS.n111 0.0135208
R9991 VSS.n2375 VSS.n2363 0.0135208
R9992 VSS.n2387 VSS.n2377 0.0135208
R9993 VSS.n2401 VSS.n2389 0.0135208
R9994 VSS.n2415 VSS.n2403 0.0135208
R9995 VSS.n2429 VSS.n2417 0.0135208
R9996 VSS.n2444 VSS.n2431 0.0135208
R9997 VSS.n2458 VSS.n2446 0.0135208
R9998 VSS.n2472 VSS.n2460 0.0135208
R9999 VSS.n2486 VSS.n2474 0.0135208
R10000 VSS.n2501 VSS.n2488 0.0135208
R10001 VSS.n2514 VSS.n2503 0.0135208
R10002 VSS.n2528 VSS.n2516 0.0135208
R10003 VSS.n2542 VSS.n2530 0.0135208
R10004 VSS.n2556 VSS.n2544 0.0135208
R10005 VSS.n2572 VSS.n2558 0.0135208
R10006 VSS.n2586 VSS.n2574 0.0135208
R10007 VSS.n2600 VSS.n2588 0.0135208
R10008 VSS.n2614 VSS.n2602 0.0135208
R10009 VSS.n2628 VSS.n2616 0.0135208
R10010 VSS.n2641 VSS.n2630 0.0135208
R10011 VSS.n2655 VSS.n2643 0.0135208
R10012 VSS.n2669 VSS.n2657 0.0135208
R10013 VSS.n2683 VSS.n2671 0.0135208
R10014 VSS.n2698 VSS.n2685 0.0135208
R10015 VSS.n2702 VSS.n2700 0.0135208
R10016 VSS.n2713 VSS.n100 0.0135208
R10017 VSS.n2727 VSS.n2715 0.0135208
R10018 VSS.n2739 VSS.n2729 0.0135208
R10019 VSS.n2753 VSS.n2741 0.0135208
R10020 VSS.n2767 VSS.n2755 0.0135208
R10021 VSS.n2781 VSS.n2769 0.0135208
R10022 VSS.n2796 VSS.n2783 0.0135208
R10023 VSS.n2810 VSS.n2798 0.0135208
R10024 VSS.n2824 VSS.n2812 0.0135208
R10025 VSS.n2838 VSS.n2826 0.0135208
R10026 VSS.n2853 VSS.n2840 0.0135208
R10027 VSS.n2866 VSS.n2855 0.0135208
R10028 VSS.n2880 VSS.n2868 0.0135208
R10029 VSS.n2894 VSS.n2882 0.0135208
R10030 VSS.n2908 VSS.n2896 0.0135208
R10031 VSS.n2924 VSS.n2910 0.0135208
R10032 VSS.n2938 VSS.n2926 0.0135208
R10033 VSS.n2952 VSS.n2940 0.0135208
R10034 VSS.n2966 VSS.n2954 0.0135208
R10035 VSS.n2980 VSS.n2968 0.0135208
R10036 VSS.n2993 VSS.n2982 0.0135208
R10037 VSS.n3007 VSS.n2995 0.0135208
R10038 VSS.n3021 VSS.n3009 0.0135208
R10039 VSS.n3035 VSS.n3023 0.0135208
R10040 VSS.n3039 VSS.n3037 0.0135208
R10041 VSS.n3054 VSS.n90 0.0135208
R10042 VSS.n3068 VSS.n3056 0.0135208
R10043 VSS.n3082 VSS.n3070 0.0135208
R10044 VSS.n3327 VSS.n3084 0.0135208
R10045 VSS.n3325 VSS.n3324 0.0135208
R10046 VSS.n3309 VSS.n3308 0.0135208
R10047 VSS.n3295 VSS.n3294 0.0135208
R10048 VSS.n3279 VSS.n3278 0.0135208
R10049 VSS.n3266 VSS.n3265 0.0135208
R10050 VSS.n3250 VSS.n3249 0.0135208
R10051 VSS.n3236 VSS.n3235 0.0135208
R10052 VSS.n3220 VSS.n3219 0.0135208
R10053 VSS.n3206 VSS.n3205 0.0135208
R10054 VSS.n3190 VSS.n3189 0.0135208
R10055 VSS.n3176 VSS.n3175 0.0135208
R10056 VSS.n3160 VSS.n3159 0.0135208
R10057 VSS.n3144 VSS.n3143 0.0135208
R10058 VSS.n3130 VSS.n3129 0.0135208
R10059 VSS.n3114 VSS.n3113 0.0135208
R10060 VSS.n3100 VSS.n3099 0.0135208
R10061 VSS.n3384 VSS.n67 0.0135208
R10062 VSS.n3388 VSS.n3386 0.0135208
R10063 VSS.n3387 VSS 0.0122188
R10064 VSS.n1149 VSS.n1148 0.0122188
R10065 VSS.n1135 VSS.n1134 0.0122188
R10066 VSS.n1119 VSS.n1118 0.0122188
R10067 VSS.n1105 VSS.n1104 0.0122188
R10068 VSS.n1091 VSS.n1090 0.0122188
R10069 VSS.n1077 VSS.n1076 0.0122188
R10070 VSS.n1063 VSS.n1062 0.0122188
R10071 VSS.n1049 VSS.n1048 0.0122188
R10072 VSS.n1035 VSS.n1034 0.0122188
R10073 VSS.n1021 VSS.n1020 0.0122188
R10074 VSS.n1007 VSS.n1006 0.0122188
R10075 VSS.n991 VSS.n990 0.0122188
R10076 VSS.n977 VSS.n976 0.0122188
R10077 VSS.n963 VSS.n962 0.0122188
R10078 VSS.n949 VSS.n948 0.0122188
R10079 VSS.n946 VSS.n945 0.0122188
R10080 VSS.n932 VSS.n931 0.0122188
R10081 VSS.n929 VSS.n928 0.0122188
R10082 VSS.n909 VSS.n175 0.0122188
R10083 VSS.n907 VSS.n906 0.0122188
R10084 VSS.n904 VSS.n903 0.0122188
R10085 VSS.n890 VSS.n889 0.0122188
R10086 VSS.n876 VSS.n875 0.0122188
R10087 VSS.n873 VSS.n872 0.0122188
R10088 VSS.n859 VSS.n858 0.0122188
R10089 VSS.n845 VSS.n844 0.0122188
R10090 VSS.n831 VSS.n830 0.0122188
R10091 VSS.n817 VSS.n816 0.0122188
R10092 VSS.n801 VSS.n800 0.0122188
R10093 VSS.n787 VSS.n786 0.0122188
R10094 VSS.n773 VSS.n772 0.0122188
R10095 VSS.n759 VSS.n758 0.0122188
R10096 VSS.n745 VSS.n744 0.0122188
R10097 VSS.n731 VSS.n730 0.0122188
R10098 VSS.n717 VSS.n716 0.0122188
R10099 VSS.n703 VSS.n702 0.0122188
R10100 VSS.n689 VSS.n688 0.0122188
R10101 VSS.n673 VSS.n672 0.0122188
R10102 VSS.n659 VSS.n658 0.0122188
R10103 VSS.n645 VSS.n644 0.0122188
R10104 VSS.n631 VSS.n630 0.0122188
R10105 VSS.n628 VSS.n627 0.0122188
R10106 VSS.n614 VSS.n613 0.0122188
R10107 VSS.n611 VSS.n610 0.0122188
R10108 VSS.n591 VSS.n220 0.0122188
R10109 VSS.n589 VSS.n588 0.0122188
R10110 VSS.n586 VSS.n585 0.0122188
R10111 VSS.n572 VSS.n571 0.0122188
R10112 VSS.n558 VSS.n557 0.0122188
R10113 VSS.n555 VSS.n554 0.0122188
R10114 VSS.n541 VSS.n540 0.0122188
R10115 VSS.n527 VSS.n526 0.0122188
R10116 VSS.n513 VSS.n512 0.0122188
R10117 VSS.n499 VSS.n498 0.0122188
R10118 VSS.n483 VSS.n482 0.0122188
R10119 VSS.n469 VSS.n468 0.0122188
R10120 VSS.n455 VSS.n454 0.0122188
R10121 VSS.n441 VSS.n440 0.0122188
R10122 VSS.n427 VSS.n426 0.0122188
R10123 VSS.n413 VSS.n412 0.0122188
R10124 VSS.n399 VSS.n398 0.0122188
R10125 VSS.n385 VSS.n384 0.0122188
R10126 VSS.n371 VSS.n370 0.0122188
R10127 VSS.n355 VSS.n354 0.0122188
R10128 VSS.n341 VSS.n340 0.0122188
R10129 VSS.n327 VSS.n326 0.0122188
R10130 VSS.n313 VSS.n312 0.0122188
R10131 VSS.n310 VSS.n309 0.0122188
R10132 VSS.n296 VSS.n295 0.0122188
R10133 VSS.n1148 VSS.n1136 0.0109167
R10134 VSS.n1134 VSS.n1120 0.0109167
R10135 VSS.n1118 VSS.n1106 0.0109167
R10136 VSS.n1104 VSS.n1092 0.0109167
R10137 VSS.n1090 VSS.n1078 0.0109167
R10138 VSS.n1076 VSS.n1064 0.0109167
R10139 VSS.n1062 VSS.n1050 0.0109167
R10140 VSS.n1048 VSS.n1036 0.0109167
R10141 VSS.n1034 VSS.n1022 0.0109167
R10142 VSS.n1020 VSS.n1008 0.0109167
R10143 VSS.n1006 VSS.n992 0.0109167
R10144 VSS.n990 VSS.n978 0.0109167
R10145 VSS.n976 VSS.n964 0.0109167
R10146 VSS.n962 VSS.n950 0.0109167
R10147 VSS.n948 VSS.n947 0.0109167
R10148 VSS.n945 VSS.n933 0.0109167
R10149 VSS.n931 VSS.n930 0.0109167
R10150 VSS.n928 VSS.n170 0.0109167
R10151 VSS.n909 VSS.n908 0.0109167
R10152 VSS.n906 VSS.n905 0.0109167
R10153 VSS.n903 VSS.n891 0.0109167
R10154 VSS.n889 VSS.n877 0.0109167
R10155 VSS.n875 VSS.n874 0.0109167
R10156 VSS.n872 VSS.n860 0.0109167
R10157 VSS.n858 VSS.n846 0.0109167
R10158 VSS.n844 VSS.n832 0.0109167
R10159 VSS.n830 VSS.n818 0.0109167
R10160 VSS.n816 VSS.n802 0.0109167
R10161 VSS.n800 VSS.n788 0.0109167
R10162 VSS.n786 VSS.n774 0.0109167
R10163 VSS.n772 VSS.n760 0.0109167
R10164 VSS.n758 VSS.n746 0.0109167
R10165 VSS.n744 VSS.n732 0.0109167
R10166 VSS.n730 VSS.n718 0.0109167
R10167 VSS.n716 VSS.n704 0.0109167
R10168 VSS.n702 VSS.n690 0.0109167
R10169 VSS.n688 VSS.n674 0.0109167
R10170 VSS.n672 VSS.n660 0.0109167
R10171 VSS.n658 VSS.n646 0.0109167
R10172 VSS.n644 VSS.n632 0.0109167
R10173 VSS.n630 VSS.n629 0.0109167
R10174 VSS.n627 VSS.n615 0.0109167
R10175 VSS.n613 VSS.n612 0.0109167
R10176 VSS.n610 VSS.n215 0.0109167
R10177 VSS.n591 VSS.n590 0.0109167
R10178 VSS.n588 VSS.n587 0.0109167
R10179 VSS.n585 VSS.n573 0.0109167
R10180 VSS.n571 VSS.n559 0.0109167
R10181 VSS.n557 VSS.n556 0.0109167
R10182 VSS.n554 VSS.n542 0.0109167
R10183 VSS.n540 VSS.n528 0.0109167
R10184 VSS.n526 VSS.n514 0.0109167
R10185 VSS.n512 VSS.n500 0.0109167
R10186 VSS.n498 VSS.n484 0.0109167
R10187 VSS.n482 VSS.n470 0.0109167
R10188 VSS.n468 VSS.n456 0.0109167
R10189 VSS.n454 VSS.n442 0.0109167
R10190 VSS.n440 VSS.n428 0.0109167
R10191 VSS.n426 VSS.n414 0.0109167
R10192 VSS.n412 VSS.n400 0.0109167
R10193 VSS.n398 VSS.n386 0.0109167
R10194 VSS.n384 VSS.n372 0.0109167
R10195 VSS.n370 VSS.n356 0.0109167
R10196 VSS.n354 VSS.n342 0.0109167
R10197 VSS.n340 VSS.n328 0.0109167
R10198 VSS.n326 VSS.n314 0.0109167
R10199 VSS.n312 VSS.n311 0.0109167
R10200 VSS.n309 VSS.n297 0.0109167
R10201 VSS.n292 VSS.n291 0.0109167
R10202 VSS.n290 VSS.n274 0.0109167
R10203 VSS.n2177 VSS.n2176 0.00961458
R10204 VSS.n2191 VSS.n2190 0.00961458
R10205 VSS.n2205 VSS.n2204 0.00961458
R10206 VSS.n2221 VSS.n2220 0.00961458
R10207 VSS.n2235 VSS.n2234 0.00961458
R10208 VSS.n2249 VSS.n2248 0.00961458
R10209 VSS.n2263 VSS.n2262 0.00961458
R10210 VSS.n2277 VSS.n2276 0.00961458
R10211 VSS.n2290 VSS.n2289 0.00961458
R10212 VSS.n2304 VSS.n2303 0.00961458
R10213 VSS.n2318 VSS.n2317 0.00961458
R10214 VSS.n2332 VSS.n2331 0.00961458
R10215 VSS.n2347 VSS.n2346 0.00961458
R10216 VSS.n2350 VSS.n2349 0.00961458
R10217 VSS.n2362 VSS.n2361 0.00961458
R10218 VSS.n2376 VSS.n2375 0.00961458
R10219 VSS.n2388 VSS.n2387 0.00961458
R10220 VSS.n2402 VSS.n2401 0.00961458
R10221 VSS.n2416 VSS.n2415 0.00961458
R10222 VSS.n2430 VSS.n2429 0.00961458
R10223 VSS.n2445 VSS.n2444 0.00961458
R10224 VSS.n2459 VSS.n2458 0.00961458
R10225 VSS.n2473 VSS.n2472 0.00961458
R10226 VSS.n2487 VSS.n2486 0.00961458
R10227 VSS.n2502 VSS.n2501 0.00961458
R10228 VSS.n2515 VSS.n2514 0.00961458
R10229 VSS.n2529 VSS.n2528 0.00961458
R10230 VSS.n2543 VSS.n2542 0.00961458
R10231 VSS.n2557 VSS.n2556 0.00961458
R10232 VSS.n2573 VSS.n2572 0.00961458
R10233 VSS.n2587 VSS.n2586 0.00961458
R10234 VSS.n2601 VSS.n2600 0.00961458
R10235 VSS.n2615 VSS.n2614 0.00961458
R10236 VSS.n2629 VSS.n2628 0.00961458
R10237 VSS.n2642 VSS.n2641 0.00961458
R10238 VSS.n2656 VSS.n2655 0.00961458
R10239 VSS.n2670 VSS.n2669 0.00961458
R10240 VSS.n2684 VSS.n2683 0.00961458
R10241 VSS.n2699 VSS.n2698 0.00961458
R10242 VSS.n2702 VSS.n2701 0.00961458
R10243 VSS.n2714 VSS.n2713 0.00961458
R10244 VSS.n2728 VSS.n2727 0.00961458
R10245 VSS.n2740 VSS.n2739 0.00961458
R10246 VSS.n2754 VSS.n2753 0.00961458
R10247 VSS.n2768 VSS.n2767 0.00961458
R10248 VSS.n2782 VSS.n2781 0.00961458
R10249 VSS.n2797 VSS.n2796 0.00961458
R10250 VSS.n2811 VSS.n2810 0.00961458
R10251 VSS.n2825 VSS.n2824 0.00961458
R10252 VSS.n2839 VSS.n2838 0.00961458
R10253 VSS.n2854 VSS.n2853 0.00961458
R10254 VSS.n2867 VSS.n2866 0.00961458
R10255 VSS.n2881 VSS.n2880 0.00961458
R10256 VSS.n2895 VSS.n2894 0.00961458
R10257 VSS.n2909 VSS.n2908 0.00961458
R10258 VSS.n2925 VSS.n2924 0.00961458
R10259 VSS.n2939 VSS.n2938 0.00961458
R10260 VSS.n2953 VSS.n2952 0.00961458
R10261 VSS.n2967 VSS.n2966 0.00961458
R10262 VSS.n2981 VSS.n2980 0.00961458
R10263 VSS.n2994 VSS.n2993 0.00961458
R10264 VSS.n3008 VSS.n3007 0.00961458
R10265 VSS.n3022 VSS.n3021 0.00961458
R10266 VSS.n3036 VSS.n3035 0.00961458
R10267 VSS.n3039 VSS.n3038 0.00961458
R10268 VSS.n3055 VSS.n3054 0.00961458
R10269 VSS.n3069 VSS.n3068 0.00961458
R10270 VSS.n3083 VSS.n3082 0.00961458
R10271 VSS.n3327 VSS.n3326 0.00961458
R10272 VSS.n3324 VSS.n3310 0.00961458
R10273 VSS.n3308 VSS.n3296 0.00961458
R10274 VSS.n3294 VSS.n3280 0.00961458
R10275 VSS.n3278 VSS.n3267 0.00961458
R10276 VSS.n3265 VSS.n3251 0.00961458
R10277 VSS.n3249 VSS.n3237 0.00961458
R10278 VSS.n3235 VSS.n3221 0.00961458
R10279 VSS.n3219 VSS.n3207 0.00961458
R10280 VSS.n3205 VSS.n3191 0.00961458
R10281 VSS.n3189 VSS.n3177 0.00961458
R10282 VSS.n3175 VSS.n3161 0.00961458
R10283 VSS.n3159 VSS.n3145 0.00961458
R10284 VSS.n3143 VSS.n3131 0.00961458
R10285 VSS.n3129 VSS.n3115 0.00961458
R10286 VSS.n3113 VSS.n3101 0.00961458
R10287 VSS.n3099 VSS.n3085 0.00961458
R10288 VSS.n3385 VSS.n3384 0.00961458
R10289 VSS.n3388 VSS.n3387 0.00961458
R10290 VSS.n294 VSS.n293 0.00701042
R10291 VSS.n11 VSS 0.00673818
R10292 VSS.n4153 VSS.n4152 0.00440625
R10293 VSS.n4150 VSS.n4147 0.00440625
R10294 VSS.n4145 VSS.n4133 0.00440625
R10295 VSS.n4131 VSS.n4120 0.00440625
R10296 VSS.n4118 VSS.n4117 0.00440625
R10297 VSS.n4115 VSS.n4105 0.00440625
R10298 VSS.n4103 VSS.n4091 0.00440625
R10299 VSS.n4089 VSS.n4077 0.00440625
R10300 VSS.n4075 VSS.n4063 0.00440625
R10301 VSS.n4061 VSS.n4060 0.00440625
R10302 VSS.n4058 VSS.n4048 0.00440625
R10303 VSS.n4046 VSS.n4034 0.00440625
R10304 VSS.n4032 VSS.n4020 0.00440625
R10305 VSS.n4018 VSS.n4006 0.00440625
R10306 VSS.n4004 VSS.n3991 0.00440625
R10307 VSS.n3989 VSS.n3977 0.00440625
R10308 VSS.n3975 VSS.n3962 0.00440625
R10309 VSS.n3960 VSS.n3948 0.00440625
R10310 VSS.n3946 VSS.n41 0.00440625
R10311 VSS.n295 VSS.n294 0.00440625
R10312 VSS.n291 VSS.n290 0.00180208
R10313 x5.X.n3 x5.X.t24 269.921
R10314 x5.X.n48 x5.X.t14 267.291
R10315 x5.X.n32 x5.X.t17 267.291
R10316 x5.X.n14 x5.X.t13 267.291
R10317 x5.X.n65 x5.X.t12 265.538
R10318 x5.X.n57 x5.X.t23 265.538
R10319 x5.X.n41 x5.X.t22 265.538
R10320 x5.X.n25 x5.X.t21 265.538
R10321 x5.X.n7 x5.X.t15 264.663
R10322 x5.X.n3 x5.X.t11 234.573
R10323 x5.X.n9 x5.X.t20 224.934
R10324 x5.X.n67 x5.X.t16 224.058
R10325 x5.X.n59 x5.X.t10 224.058
R10326 x5.X.n43 x5.X.t9 224.058
R10327 x5.X.n27 x5.X.t8 224.058
R10328 x5.X.n50 x5.X.t19 222.304
R10329 x5.X.n34 x5.X.t25 222.304
R10330 x5.X.n16 x5.X.t18 222.304
R10331 x5.X.n74 x5.X.n72 197.595
R10332 x5.X.n74 x5.X.n73 167.416
R10333 x5.X.n78 x5.X.n76 138.054
R10334 x5.X x5.X.n77 106.453
R10335 x5.X.n4 x5.X.n3 76.0005
R10336 x5.X.n72 x5.X.t2 26.5955
R10337 x5.X.n72 x5.X.t0 26.5955
R10338 x5.X.n73 x5.X.t3 26.5955
R10339 x5.X.n73 x5.X.t1 26.5955
R10340 x5.X.n76 x5.X.t4 24.9236
R10341 x5.X.n76 x5.X.t6 24.9236
R10342 x5.X.n77 x5.X.t5 24.9236
R10343 x5.X.n77 x5.X.t7 24.9236
R10344 x5.X.n22 x5.X 21.2667
R10345 x5.X.n75 x5.X.n71 12.466
R10346 x5.X.n50 x5.X.n49 12.2696
R10347 x5.X.n34 x5.X.n33 12.2696
R10348 x5.X.n16 x5.X.n15 12.2696
R10349 x5.X.n38 x5.X.n22 10.5535
R10350 x5.X.n54 x5.X.n38 10.5535
R10351 x5.X.n67 x5.X.n66 10.5169
R10352 x5.X.n59 x5.X.n58 10.5169
R10353 x5.X.n43 x5.X.n42 10.5169
R10354 x5.X.n27 x5.X.n26 10.5169
R10355 x5.X.n62 x5.X.n54 10.4999
R10356 x5.X.n9 x5.X.n8 9.6405
R10357 x5.X.n44 x5.X.n43 9.3005
R10358 x5.X.n28 x5.X.n27 9.3005
R10359 x5.X.n68 x5.X.n67 8.76429
R10360 x5.X.n60 x5.X.n59 8.76429
R10361 x5.X.n51 x5.X.n50 8.76429
R10362 x5.X.n35 x5.X.n34 8.76429
R10363 x5.X.n10 x5.X.n9 8.76429
R10364 x5.X.n17 x5.X.n16 8.76429
R10365 x5.X.n71 x5.X.n62 7.58473
R10366 x5.X x5.X.n4 7.57233
R10367 x5.X.n53 x5.X.n52 7.52485
R10368 x5.X.n19 x5.X.n18 7.5187
R10369 x5.X.n37 x5.X.n36 7.45404
R10370 x5.X x5.X.n78 7.3702
R10371 x5.X.n71 x5.X.n0 7.19295
R10372 x5.X.n46 x5.X 7.03149
R10373 x5.X.n30 x5.X 7.03149
R10374 x5.X.n12 x5.X 7.03149
R10375 x5.X.n63 x5.X 6.67092
R10376 x5.X.n55 x5.X 6.67092
R10377 x5.X.n39 x5.X 6.67092
R10378 x5.X.n23 x5.X 6.67092
R10379 x5.X.n62 x5.X.n61 6.55969
R10380 x5.X.n5 x5.X 6.49064
R10381 x5.X.n75 x5.X 6.46515
R10382 x5.X.n0 x5.X.n69 5.26654
R10383 x5.X.n8 x5.X.n7 5.25868
R10384 x5.X.n4 x5.X 4.68782
R10385 x5.X.n38 x5.X.n2 4.38498
R10386 x5.X.n66 x5.X.n65 4.38232
R10387 x5.X.n58 x5.X.n57 4.38232
R10388 x5.X.n42 x5.X.n41 4.38232
R10389 x5.X.n26 x5.X.n25 4.38232
R10390 x5.X.n54 x5.X.n1 4.38051
R10391 x5.X.n22 x5.X.n21 4.35575
R10392 x5.X.n2 x5.X.n29 3.43448
R10393 x5.X.n1 x5.X.n45 3.43273
R10394 x5.X.n20 x5.X.n11 5.18552
R10395 x5.X.n49 x5.X.n48 2.62959
R10396 x5.X.n33 x5.X.n32 2.62959
R10397 x5.X.n15 x5.X.n14 2.62959
R10398 x5.X.n51 x5.X.n47 2.52444
R10399 x5.X.n35 x5.X.n31 2.52444
R10400 x5.X.n17 x5.X.n13 2.52444
R10401 x5.X x5.X.n75 2.32777
R10402 x5.X.n69 x5.X.n68 2.27475
R10403 x5.X.n0 x5.X.n70 2.26611
R10404 x5.X.n11 x5.X.n10 2.20216
R10405 x5.X x5.X.n74 2.19848
R10406 x5.X.n68 x5.X.n64 2.16388
R10407 x5.X.n60 x5.X.n56 2.16388
R10408 x5.X.n44 x5.X.n40 2.16388
R10409 x5.X.n28 x5.X.n24 2.16388
R10410 x5.X.n10 x5.X.n6 1.9836
R10411 x5.X.n29 x5.X.n28 1.45136
R10412 x5.X.n78 x5.X 1.42272
R10413 x5.X.n45 x5.X.n44 1.38585
R10414 x5.X.n6 x5.X.n5 1.08219
R10415 x5.X.n61 x5.X.n60 1.0658
R10416 x5.X.n61 x5.X 0.932428
R10417 x5.X.n52 x5.X 0.930853
R10418 x5.X.n18 x5.X 0.919788
R10419 x5.X.n36 x5.X 0.919522
R10420 x5.X.n64 x5.X.n63 0.901908
R10421 x5.X.n56 x5.X.n55 0.901908
R10422 x5.X.n40 x5.X.n39 0.901908
R10423 x5.X.n24 x5.X.n23 0.901908
R10424 x5.X.n36 x5.X.n35 0.850177
R10425 x5.X.n18 x5.X.n17 0.849917
R10426 x5.X.n52 x5.X.n51 0.843446
R10427 x5.X.n45 x5.X 0.801859
R10428 x5.X.n29 x5.X 0.71223
R10429 x5.X.n47 x5.X.n46 0.541345
R10430 x5.X.n31 x5.X.n30 0.541345
R10431 x5.X.n13 x5.X.n12 0.541345
R10432 x5.X.n11 x5.X 0.469125
R10433 x5.X.n69 x5.X 0.242354
R10434 x5.X.n2 x5.X.n37 0.0624655
R10435 x5.X.n1 x5.X.n53 0.0624655
R10436 x5.X.n20 x5.X.n19 0.0421667
R10437 x5.X.n21 x5.X.n20 0.0402727
R10438 x4.X.n38 x4.X.n22 585
R10439 x4.X.n24 x4.X.t66 397.144
R10440 x4.X.n31 x4.X.t50 394.462
R10441 x4.X.n39 x4.X.n37 302.474
R10442 x4.X.n124 x4.X.t41 209.331
R10443 x4.X.n89 x4.X.t36 208.625
R10444 x4.X.n178 x4.X.t59 208.013
R10445 x4.X.n96 x4.X.t33 207.919
R10446 x4.X.n62 x4.X.t58 207.919
R10447 x4.X.n69 x4.X.t55 207.919
R10448 x4.X.n117 x4.X.t42 207.915
R10449 x4.X.n144 x4.X.t56 207.911
R10450 x4.X.n171 x4.X.t47 207.853
R10451 x4.X.n152 x4.X.t53 206.475
R10452 x4.X.n134 x4.X.t61 202.565
R10453 x4.X.n106 x4.X.t49 202.565
R10454 x4.X.n111 x4.X.t67 202.565
R10455 x4.X.n83 x4.X.t60 202.565
R10456 x4.X.n164 x4.X.t62 202.163
R10457 x4.X.n139 x4.X.t43 202.163
R10458 x4.X.n78 x4.X.t39 202.163
R10459 x4.X.n152 x4.X.t40 179.695
R10460 x4.X.n178 x4.X.t44 179.094
R10461 x4.X.n144 x4.X.t35 178.258
R10462 x4.X.n117 x4.X.t64 178.256
R10463 x4.X.n96 x4.X.t63 178.252
R10464 x4.X.n62 x4.X.t45 178.252
R10465 x4.X.n69 x4.X.t51 178.252
R10466 x4.X.n165 x4.X.t48 177.588
R10467 x4.X.n170 x4.X.t68 177.588
R10468 x4.X.n140 x4.X.t65 177.588
R10469 x4.X.n79 x4.X.t34 177.588
R10470 x4.X.n89 x4.X.t57 177.536
R10471 x4.X.n135 x4.X.t46 176.834
R10472 x4.X.n107 x4.X.t69 176.834
R10473 x4.X.n112 x4.X.t52 176.834
R10474 x4.X.n84 x4.X.t54 176.834
R10475 x4.X.n124 x4.X.t38 176.816
R10476 x4.X.n19 x4.X.n17 146.811
R10477 x4.X.n40 x4.X.n39 143.149
R10478 x4.X.n24 x4.X.t32 134.986
R10479 x4.X.n31 x4.X.t37 134.484
R10480 x4.X.n19 x4.X.n18 108.412
R10481 x4.X.n21 x4.X.n20 108.412
R10482 x4.X.n45 x4.X.n13 108.412
R10483 x4.X.n44 x4.X.n14 108.412
R10484 x4.X.n43 x4.X.n15 108.412
R10485 x4.X.n42 x4.X.n16 108.412
R10486 x4.X.n48 x4.X.n46 90.8321
R10487 x4.X.n48 x4.X.n47 52.4321
R10488 x4.X.n50 x4.X.n49 52.4321
R10489 x4.X.n52 x4.X.n51 52.4321
R10490 x4.X.n54 x4.X.n53 52.4321
R10491 x4.X.n56 x4.X.n55 52.4321
R10492 x4.X.n58 x4.X.n57 52.4321
R10493 x4.X.n60 x4.X.n59 52.4321
R10494 x4.X.n50 x4.X.n48 38.4005
R10495 x4.X.n52 x4.X.n50 38.4005
R10496 x4.X.n54 x4.X.n52 38.4005
R10497 x4.X.n56 x4.X.n54 38.4005
R10498 x4.X.n58 x4.X.n56 38.4005
R10499 x4.X.n60 x4.X.n58 38.4005
R10500 x4.X.n45 x4.X.n44 38.4005
R10501 x4.X.n44 x4.X.n43 38.4005
R10502 x4.X.n43 x4.X.n42 38.4005
R10503 x4.X.n21 x4.X.n19 38.4005
R10504 x4.X.n41 x4.X.n21 38.4005
R10505 x4.X.n42 x4.X.n41 38.4005
R10506 x4.X x4.X.n45 33.7342
R10507 x4.X.n181 x4.X.n60 30.8711
R10508 x4.X.n13 x4.X.t4 26.5955
R10509 x4.X.n13 x4.X.t10 26.5955
R10510 x4.X.n14 x4.X.t3 26.5955
R10511 x4.X.n14 x4.X.t14 26.5955
R10512 x4.X.n15 x4.X.t11 26.5955
R10513 x4.X.n15 x4.X.t2 26.5955
R10514 x4.X.n16 x4.X.t7 26.5955
R10515 x4.X.n16 x4.X.t0 26.5955
R10516 x4.X.n17 x4.X.t6 26.5955
R10517 x4.X.n17 x4.X.t1 26.5955
R10518 x4.X.n18 x4.X.t8 26.5955
R10519 x4.X.n18 x4.X.t12 26.5955
R10520 x4.X.n20 x4.X.t9 26.5955
R10521 x4.X.n20 x4.X.t13 26.5955
R10522 x4.X.n46 x4.X.t18 24.9236
R10523 x4.X.n46 x4.X.t29 24.9236
R10524 x4.X.n47 x4.X.t20 24.9236
R10525 x4.X.n47 x4.X.t24 24.9236
R10526 x4.X.n49 x4.X.t21 24.9236
R10527 x4.X.n49 x4.X.t25 24.9236
R10528 x4.X.n51 x4.X.t17 24.9236
R10529 x4.X.n51 x4.X.t27 24.9236
R10530 x4.X.n53 x4.X.t19 24.9236
R10531 x4.X.n53 x4.X.t28 24.9236
R10532 x4.X.n55 x4.X.t23 24.9236
R10533 x4.X.n55 x4.X.t30 24.9236
R10534 x4.X.n57 x4.X.t31 24.9236
R10535 x4.X.n57 x4.X.t26 24.9236
R10536 x4.X.n59 x4.X.t16 24.9236
R10537 x4.X.n59 x4.X.t22 24.9236
R10538 x4.X.n23 x4.X.t5 22.6555
R10539 x4.X.n180 x4.X.n179 19.9012
R10540 x4.X.n10 x4.X.n11 3.58524
R10541 x4.X.n181 x4.X.n180 19.6126
R10542 x4.X.n38 x4.X.t15 13.7905
R10543 x4.X.n27 x4.X 13.6005
R10544 x4.X.n39 x4.X.n38 12.8055
R10545 x4.X.n142 x4.X.n141 10.4992
R10546 x4.X.n114 x4.X.n113 10.4947
R10547 x4.X.n86 x4.X.n85 10.4903
R10548 x4.X.n41 x4.X.n40 9.82233
R10549 x4.X x4.X.n181 9.6005
R10550 x4.X.n8 x4.X.n7 1.83978
R10551 x4.X.n26 x4.X.n25 9.3005
R10552 x4.X.n33 x4.X.n32 9.3005
R10553 x4.X.n166 x4.X.n165 9.3005
R10554 x4.X.n136 x4.X.n135 9.3005
R10555 x4.X.n141 x4.X.n140 9.3005
R10556 x4.X.n108 x4.X.n107 9.3005
R10557 x4.X.n113 x4.X.n112 9.3005
R10558 x4.X.n80 x4.X.n79 9.3005
R10559 x4.X.n85 x4.X.n84 9.3005
R10560 x4.X.n35 x4.X.n22 9.3005
R10561 x4.X.n23 x4.X.n22 9.3005
R10562 x4.X.n179 x4.X 9.18311
R10563 x4.X.n179 x4.X.n178 8.76429
R10564 x4.X.n87 x4.X.n75 8.41509
R10565 x4.X.n40 x4.X.n22 8.16186
R10566 x4.X.n172 x4.X.n171 7.61316
R10567 x4.X.n135 x4.X.n134 7.35553
R10568 x4.X.n107 x4.X.n106 7.35553
R10569 x4.X.n112 x4.X.n111 7.35553
R10570 x4.X.n84 x4.X.n83 7.35553
R10571 x4.X.n153 x4.X.n152 7.32997
R10572 x4.X.n97 x4.X.n96 7.28785
R10573 x4.X.n63 x4.X.n62 7.28785
R10574 x4.X.n70 x4.X.n69 7.28785
R10575 x4.X.n118 x4.X.n117 7.27968
R10576 x4.X.n145 x4.X.n144 7.27145
R10577 x4.X.n90 x4.X.n89 7.25084
R10578 x4.X.n125 x4.X.n124 7.2225
R10579 x4.X.n32 x4.X.n31 6.9915
R10580 x4.X.n26 x4.X.n24 6.95412
R10581 x4.X.n165 x4.X.n164 6.95331
R10582 x4.X.n140 x4.X.n139 6.95331
R10583 x4.X.n79 x4.X.n78 6.95331
R10584 x4.X.n115 x4.X.n103 6.17402
R10585 x4.X.n143 x4.X.n131 6.14277
R10586 x4.X.n177 x4.X.n161 6.12937
R10587 x4.X.n142 x4.X.n136 6.09927
R10588 x4.X.n86 x4.X.n80 6.09034
R10589 x4.X.n176 x4.X.n175 5.93026
R10590 x4.X.n114 x4.X.n108 5.83458
R10591 x4.X.n146 x4.X 5.56572
R10592 x4.X.n154 x4.X 5.56572
R10593 x4.X.n119 x4.X 5.28746
R10594 x4.X.n126 x4.X 5.28746
R10595 x4.X.n91 x4.X 5.28746
R10596 x4.X.n132 x4.X 5.0092
R10597 x4.X.n98 x4.X 5.0092
R10598 x4.X.n76 x4.X 5.0092
R10599 x4.X.n81 x4.X 5.0092
R10600 x4.X.n64 x4.X 5.0092
R10601 x4.X.n71 x4.X 5.0092
R10602 x4.X.n162 x4.X 4.73093
R10603 x4.X.n172 x4.X.n169 4.73093
R10604 x4.X.n137 x4.X 4.73093
R10605 x4.X.n104 x4.X 4.73093
R10606 x4.X.n109 x4.X 4.73093
R10607 x4.X.n160 x4.X.n151 4.62479
R10608 x4.X.n102 x4.X.n94 4.61713
R10609 x4.X.n130 x4.X.n122 4.6082
R10610 x4.X.n75 x4.X.n67 4.6082
R10611 x4.X.n36 x4.X.n35 4.5327
R10612 x4.X.n12 x4.X.n22 9.31609
R10613 x4.X x4.X.n11 2.9629
R10614 x4.X.n163 x4.X.n162 4.45267
R10615 x4.X.n169 x4.X 4.45267
R10616 x4.X.n138 x4.X.n137 4.45267
R10617 x4.X.n105 x4.X.n104 4.45267
R10618 x4.X.n110 x4.X.n109 4.45267
R10619 x4.X.n176 x4.X.n166 4.42753
R10620 x4.X.n161 x4.X.n143 4.25884
R10621 x4.X.n131 x4.X.n115 4.24991
R10622 x4.X.n103 x4.X.n87 4.21866
R10623 x4.X.n133 x4.X.n132 4.17441
R10624 x4.X.n77 x4.X.n76 4.17441
R10625 x4.X.n82 x4.X.n81 4.17441
R10626 x4.X.n39 x4.X.n23 3.9405
R10627 x4.X.n147 x4.X.n146 3.61789
R10628 x4.X.n155 x4.X.n154 3.33963
R10629 x4.X.n120 x4.X.n119 3.33963
R10630 x4.X.n127 x4.X.n126 3.06137
R10631 x4.X.n92 x4.X.n91 3.06137
R10632 x4.X.n99 x4.X.n98 3.06137
R10633 x4.X.n65 x4.X.n64 3.06137
R10634 x4.X.n72 x4.X.n71 3.06137
R10635 x4.X.n149 x4.X.n147 3.04032
R10636 x4.X.n174 x4.X.n173 3.035
R10637 x4.X.n157 x4.X.n155 3.035
R10638 x4.X.n5 x4.X.n120 3.03311
R10639 x4.X.n0 x4.X.n127 3.03311
R10640 x4.X.n1 x4.X.n92 3.03311
R10641 x4.X.n2 x4.X.n99 3.03311
R10642 x4.X.n3 x4.X.n65 3.03311
R10643 x4.X.n4 x4.X.n72 3.03311
R10644 x4.X.n29 x4.X.n28 3.00943
R10645 x4.X.n8 x4.X 4.1629
R10646 x4.X.n37 x4.X.n9 2.62757
R10647 x4.X.n27 x4.X.n26 2.52171
R10648 x4.X.n32 x4.X.n8 1.54783
R10649 x4.X.n12 x4.X.n36 1.50334
R10650 x4.X.n87 x4.X.n86 2.2505
R10651 x4.X.n103 x4.X.n102 2.2505
R10652 x4.X.n115 x4.X.n114 2.2505
R10653 x4.X.n131 x4.X.n130 2.2505
R10654 x4.X.n143 x4.X.n142 2.2505
R10655 x4.X.n161 x4.X.n160 2.2505
R10656 x4.X.n177 x4.X.n176 2.2505
R10657 x4.X.n175 x4.X.n174 2.23927
R10658 x4.X.n34 x4.X.n9 2.23869
R10659 x4.X.n180 x4.X.n177 2.16478
R10660 x4.X.n160 x4.X.n159 2.07162
R10661 x4.X.n75 x4.X.n74 2.045
R10662 x4.X.n102 x4.X.n101 2.04053
R10663 x4.X.n130 x4.X.n129 2.02268
R10664 x4.X.n37 x4.X.n22 1.76715
R10665 x4.X.n29 x4.X 1.72692
R10666 x4.X.n127 x4.X.n125 1.67007
R10667 x4.X.n92 x4.X.n90 1.67007
R10668 x4.X.n99 x4.X.n97 1.67007
R10669 x4.X.n65 x4.X.n63 1.67007
R10670 x4.X.n72 x4.X.n70 1.67007
R10671 x4.X.n34 x4.X.n6 1.57957
R10672 x4.X.n7 x4.X.n6 0.896263
R10673 x4.X.n121 x4.X.n5 1.50237
R10674 x4.X.n128 x4.X.n0 1.50174
R10675 x4.X.n93 x4.X.n1 1.50174
R10676 x4.X.n100 x4.X.n2 1.50174
R10677 x4.X.n66 x4.X.n3 1.50174
R10678 x4.X.n73 x4.X.n4 1.50174
R10679 x4.X.n159 x4.X.n157 1.49811
R10680 x4.X.n151 x4.X.n149 1.49801
R10681 x4.X.n155 x4.X.n153 1.3918
R10682 x4.X.n120 x4.X.n118 1.3918
R10683 x4.X.n147 x4.X.n145 1.11354
R10684 x4.X.n171 x4.X.n170 0.72374
R10685 x4.X.n136 x4.X.n133 0.557022
R10686 x4.X.n80 x4.X.n77 0.557022
R10687 x4.X.n85 x4.X.n82 0.557022
R10688 x4.X.n27 x4.X.n11 0.300347
R10689 x4.X.n166 x4.X.n163 0.278761
R10690 x4.X.n173 x4.X.n172 0.278761
R10691 x4.X.n141 x4.X.n138 0.278761
R10692 x4.X.n108 x4.X.n105 0.278761
R10693 x4.X.n113 x4.X.n110 0.278761
R10694 x4.X.n28 x4.X 0.259429
R10695 x4.X.n28 x4.X.n10 0.076587
R10696 x4.X.n25 x4.X.n10 0.0466957
R10697 x4.X.n25 x4.X 0.0358261
R10698 x4.X.n7 x4.X.n33 0.0347909
R10699 x4.X.n175 x4.X.n167 0.0291789
R10700 x4.X.n36 x4.X.n34 0.0279871
R10701 x4.X.n122 x4.X.n121 0.0269367
R10702 x4.X.n94 x4.X.n93 0.0269367
R10703 x4.X.n67 x4.X.n66 0.0269367
R10704 x4.X.n129 x4.X.n128 0.0257706
R10705 x4.X.n101 x4.X.n100 0.0257706
R10706 x4.X.n74 x4.X.n73 0.0257706
R10707 x4.X.n6 x4.X.n30 4.51062
R10708 x4.X.n5 x4.X.n116 0.0271977
R10709 x4.X.n4 x4.X.n68 0.0259313
R10710 x4.X.n3 x4.X.n61 0.0259313
R10711 x4.X.n2 x4.X.n95 0.0259313
R10712 x4.X.n1 x4.X.n88 0.0259313
R10713 x4.X.n0 x4.X.n123 0.0259313
R10714 x4.X.n149 x4.X.n148 0.0245385
R10715 x4.X.n9 x4.X.n12 0.00855895
R10716 x4.X.n33 x4.X.n30 0.0217264
R10717 x4.X.n157 x4.X.n156 0.0213333
R10718 x4.X.n30 x4.X 0.0170094
R10719 x4.X.n159 x4.X.n158 0.016693
R10720 x4.X.n174 x4.X.n168 0.0152198
R10721 x4.X.n151 x4.X.n150 0.0144347
R10722 x4.X.n35 x4.X.n9 0.0109693
R10723 x4.X x4.X.n29 0.00993396
R10724 check[5].n1 check[5].t3 331.51
R10725 check[5].n1 check[5].t2 209.403
R10726 check[5].n0 check[5].t0 207.373
R10727 check[5].n2 check[5].n1 76.0005
R10728 check[5].n4 check[5].n3 50.8596
R10729 check[5].n5 check[5].t1 31.153
R10730 check[5].n4 check[5] 18.2949
R10731 check[5].n3 check[5] 13.2142
R10732 check[5].n3 check[5] 12.3082
R10733 check[5] check[5].n0 9.01934
R10734 check[5] check[5].n2 8.58587
R10735 check[5] check[5].n5 7.78567
R10736 check[5].n0 check[5] 7.45876
R10737 check[5].n2 check[5] 2.02977
R10738 check[5].n5 check[5].n4 1.33351
R10739 check[0].n3 check[0].t5 373.283
R10740 check[0].n1 check[0].t3 331.51
R10741 check[0].n1 check[0].t2 209.403
R10742 check[0].n0 check[0].t0 207.373
R10743 check[0].n3 check[0].t4 132.282
R10744 check[0].n4 check[0].n3 84.146
R10745 check[0].n2 check[0].n1 76.0005
R10746 check[0].n8 check[0].n7 48.6767
R10747 check[0].n9 check[0].t1 33.3302
R10748 check[0].n6 check[0].n5 19.508
R10749 check[0].n8 check[0] 15.1737
R10750 check[0].n5 check[0].n4 13.3958
R10751 check[0].n7 check[0] 12.062
R10752 check[0] check[0].n9 9.55531
R10753 check[0] check[0].n0 9.01934
R10754 check[0].n6 check[0] 8.69451
R10755 check[0] check[0].n2 8.58587
R10756 check[0].n0 check[0] 7.45876
R10757 check[0].n5 check[0] 6.84701
R10758 check[0].n4 check[0] 4.07323
R10759 check[0].n7 check[0].n6 3.04048
R10760 check[0].n2 check[0] 2.02977
R10761 check[0].n9 check[0].n8 1.77306
R10762 check[2].n3 check[2].t5 331.51
R10763 check[2].n1 check[2].t3 299.377
R10764 check[2].n3 check[2].t4 209.403
R10765 check[2].n0 check[2].t0 207.373
R10766 check[2].n1 check[2].t2 206.19
R10767 check[2] check[2].n1 105.007
R10768 check[2].n4 check[2].n3 76.0005
R10769 check[2].n7 check[2].n6 49.7951
R10770 check[2].n5 check[2].n2 47.9541
R10771 check[2].n8 check[2].t1 31.8695
R10772 check[2].n7 check[2] 15.2244
R10773 check[2].n6 check[2] 11.8159
R10774 check[2].n2 check[2] 11.1489
R10775 check[2] check[2].n0 9.01934
R10776 check[2] check[2].n8 8.9196
R10777 check[2].n5 check[2] 8.84542
R10778 check[2] check[2].n4 8.58587
R10779 check[2].n0 check[2] 7.45876
R10780 check[2].n6 check[2].n5 3.04357
R10781 check[2].n2 check[2] 2.89082
R10782 check[2].n4 check[2] 2.02977
R10783 check[2].n8 check[2].n7 1.63044
R10784 D[2].n3 D[2].t2 269.921
R10785 D[2].n3 D[2].t3 234.573
R10786 D[2].n10 D[2].t0 207.373
R10787 D[2].n11 D[2] 59.1407
R10788 D[2].n13 D[2].t1 32.581
R10789 D[2] D[2].n13 9.80687
R10790 D[2] D[2].n10 9.01934
R10791 D[2].n4 D[2].n3 8.76429
R10792 D[2].n4 D[2] 7.57233
R10793 D[2].n10 D[2] 7.45876
R10794 D[2].n4 D[2] 4.68782
R10795 D[2].n12 D[2].n11 3.84831
R10796 D[2].n5 D[2].n4 3.77218
R10797 D[2].n6 D[2].n5 3.26839
R10798 D[2].n5 D[2] 3.23635
R10799 D[2].n11 D[2].n9 2.92915
R10800 D[2].n8 D[2].n1 2.26284
R10801 D[2].n7 D[2].n6 2.23869
R10802 D[2].n13 D[2].n12 0.389891
R10803 D[2].n7 D[2].n2 0.0232273
R10804 D[2].n9 D[2].n0 0.00807576
R10805 D[2].n8 D[2].n7 0.00195195
R10806 D[2].n9 D[2].n8 0.00194159
R10807 check[3].n7 check[3].t0 417.519
R10808 check[3].n1 check[3].t3 331.51
R10809 check[3].n1 check[3].t2 209.403
R10810 check[3].t0 check[3].n6 137.702
R10811 check[3].n2 check[3].n1 76.0005
R10812 check[3].n8 check[3] 60.7393
R10813 check[3].n9 check[3].t1 35.4919
R10814 check[3].n8 check[3] 18.329
R10815 check[3].n7 check[3].n0 12.3082
R10816 check[3].n3 check[3] 12.0607
R10817 check[3] check[3].n9 9.48284
R10818 check[3].n4 check[3].n0 9.3005
R10819 check[3].n6 check[3].n3 9.3005
R10820 check[3] check[3].n2 8.58587
R10821 check[3].n5 check[3].n4 4.59955
R10822 check[3] check[3].n0 2.70819
R10823 check[3].n2 check[3] 2.02977
R10824 check[3].n9 check[3].n8 1.84729
R10825 check[3] check[3].n7 1.72358
R10826 check[3].n5 check[3] 1.353
R10827 check[3].n6 check[3].n5 0.122715
R10828 check[3].n4 check[3].n3 0.00847872
R10829 check[6].n3 check[6].t3 331.51
R10830 check[6].n3 check[6].t2 209.403
R10831 check[6].n2 check[6].t0 207.373
R10832 check[6].n4 check[6].n3 76.0005
R10833 check[6].n6 check[6].n5 48.5667
R10834 check[6].n9 check[6].t1 31.8564
R10835 check[6].n0 check[6] 16.649
R10836 check[6].n5 check[6] 13.5264
R10837 check[6].n5 check[6] 11.8159
R10838 check[6] check[6].n2 9.01934
R10839 check[6] check[6].n9 8.94887
R10840 check[6] check[6].n4 8.58587
R10841 check[6].n2 check[6] 7.45876
R10842 check[6].n6 check[6].n1 4.3624
R10843 check[6].n8 check[6].n7 2.95435
R10844 check[6].n4 check[6] 2.02977
R10845 check[6].n7 check[6].n6 0.578192
R10846 check[6].n9 check[6].n8 0.290433
R10847 check[6].n1 check[6].n0 0.0421667
R10848 D[1].n8 D[1].t2 269.921
R10849 D[1].n8 D[1].t3 234.573
R10850 D[1].n7 D[1].t0 207.373
R10851 D[1].n9 D[1].n8 76.0005
R10852 D[1].n13 D[1].t1 33.3405
R10853 D[1].n11 D[1].n10 23.4
R10854 D[1].n10 D[1] 22.0971
R10855 D[1].n10 D[1].n9 14.9338
R10856 D[1] D[1].n13 9.32876
R10857 D[1] D[1].n7 9.01934
R10858 D[1].n9 D[1] 7.57233
R10859 D[1].n7 D[1] 7.45876
R10860 D[1].n3 D[1] 6.54947
R10861 D[1].n9 D[1] 4.68782
R10862 D[1].n12 D[1].n11 3.67573
R10863 D[1].n11 D[1].n6 2.87957
R10864 D[1].n5 D[1].n1 2.26284
R10865 D[1].n4 D[1].n3 2.23869
R10866 D[1].n13 D[1].n12 0.391757
R10867 D[1].n4 D[1].n2 0.0213333
R10868 D[1].n6 D[1].n0 0.0099697
R10869 D[1].n5 D[1].n4 0.00195195
R10870 D[1].n6 D[1].n5 0.00194159
R10871 reset.n0 reset.t0 259.634
R10872 reset.n0 reset.t1 175.183
R10873 reset.n1 reset.n0 8.19557
R10874 reset.n1 reset 2.53088
R10875 reset reset.n1 2.48048
R10876 check[4].n1 check[4].t3 331.51
R10877 check[4].n1 check[4].t2 209.403
R10878 check[4].n0 check[4].t0 207.373
R10879 check[4].n2 check[4].n1 76.0005
R10880 check[4].n4 check[4].n3 48.1851
R10881 check[4].n5 check[4].t1 34.0601
R10882 check[4].n4 check[4] 18.3315
R10883 check[4].n3 check[4] 13.0581
R10884 check[4].n3 check[4] 12.5543
R10885 check[4] check[4].n5 9.53084
R10886 check[4] check[4].n0 9.01934
R10887 check[4] check[4].n2 8.58587
R10888 check[4].n0 check[4] 7.45876
R10889 check[4].n2 check[4] 2.02977
R10890 check[4].n5 check[4].n4 1.79774
R10891 D[5].n8 D[5].t2 269.921
R10892 D[5].n8 D[5].t3 234.573
R10893 D[5].n7 D[5].t0 207.373
R10894 D[5].n9 D[5].n8 76.0005
R10895 D[5].n14 D[5].t1 34.8263
R10896 D[5].n11 D[5] 23.5855
R10897 D[5].n12 D[5].n11 23.0768
R10898 D[5].n11 D[5].n10 14.6672
R10899 D[5] D[5].n7 9.01934
R10900 D[5] D[5].n14 8.60331
R10901 D[5].n9 D[5] 7.57233
R10902 D[5].n7 D[5] 7.45876
R10903 D[5].n10 D[5] 3.78642
R10904 D[5].n13 D[5].n12 3.14374
R10905 D[5].n3 D[5] 3.01822
R10906 D[5].n12 D[5].n6 2.74043
R10907 D[5].n5 D[5].n1 2.26284
R10908 D[5].n4 D[5].n3 2.23869
R10909 D[5].n10 D[5].n9 0.901908
R10910 D[5].n14 D[5].n13 0.398471
R10911 D[5].n6 D[5].n0 0.0232273
R10912 D[5].n4 D[5].n2 0.00807576
R10913 D[5].n5 D[5].n4 0.00195195
R10914 D[5].n6 D[5].n5 0.00194159
R10915 D[4].n8 D[4].t2 269.921
R10916 D[4].n8 D[4].t3 234.573
R10917 D[4].n7 D[4].t0 207.373
R10918 D[4].n9 D[4].n8 76.0005
R10919 D[4].n14 D[4].t1 33.3509
R10920 D[4].n11 D[4] 23.2878
R10921 D[4].n12 D[4].n11 22.7446
R10922 D[4].n11 D[4].n10 14.6672
R10923 D[4] D[4].n14 9.10171
R10924 D[4] D[4].n7 9.01934
R10925 D[4].n9 D[4] 7.57233
R10926 D[4].n7 D[4] 7.45876
R10927 D[4].n10 D[4] 3.9667
R10928 D[4].n13 D[4].n12 3.32332
R10929 D[4].n12 D[4].n6 2.78529
R10930 D[4].n3 D[4] 2.75482
R10931 D[4].n5 D[4].n1 2.26284
R10932 D[4].n4 D[4].n3 2.23869
R10933 D[4].n10 D[4].n9 0.721627
R10934 D[4].n14 D[4].n13 0.379298
R10935 D[4].n6 D[4].n0 0.0251212
R10936 D[4].n4 D[4].n2 0.00618182
R10937 D[4].n5 D[4].n4 0.00195195
R10938 D[4].n6 D[4].n5 0.00194159
R10939 sel_bit[1].t1 sel_bit[1].t3 769.593
R10940 sel_bit[1].n4 sel_bit[1].t2 367.928
R10941 sel_bit[1].n2 sel_bit[1].t1 339.695
R10942 sel_bit[1].n4 sel_bit[1].t0 112.237
R10943 sel_bit[1].n5 sel_bit[1].n4 22.0348
R10944 sel_bit[1].n7 sel_bit[1] 15.3177
R10945 sel_bit[1].n5 sel_bit[1].n3 12.3948
R10946 sel_bit[1].n3 sel_bit[1].n2 11.0176
R10947 sel_bit[1].n6 sel_bit[1].n5 8.76429
R10948 sel_bit[1].n0 sel_bit[1] 5.95912
R10949 sel_bit[1] sel_bit[1].n7 3.41725
R10950 sel_bit[1].n6 sel_bit[1].n1 1.98671
R10951 sel_bit[1].n1 sel_bit[1].n0 1.76602
R10952 sel_bit[1].n7 sel_bit[1].n6 1.07617
R10953 D[7].n0 D[7].t0 207.373
R10954 D[7].n1 D[7] 66.6056
R10955 D[7].n1 D[7].t1 34.2054
R10956 D[7] D[7].n0 9.01934
R10957 D[7].n0 D[7] 7.45876
R10958 D[7].n10 D[7].n9 4.18512
R10959 D[7].n9 D[7].n8 3.02821
R10960 D[7].n4 D[7] 2.91107
R10961 D[7].n6 D[7].n2 2.26284
R10962 D[7].n5 D[7].n4 2.23869
R10963 D[7] D[7].n10 2.21588
R10964 D[7].n9 D[7].n1 0.253183
R10965 D[7].n8 D[7].n7 0.00901436
R10966 D[7].n5 D[7].n3 0.00618182
R10967 D[7].n6 D[7].n5 0.00195195
R10968 D[7].n7 D[7].n6 0.00194159
R10969 D[6].n8 D[6].t2 269.921
R10970 D[6].n8 D[6].t3 234.573
R10971 D[6].n7 D[6].t0 207.373
R10972 D[6].n9 D[6].n8 76.0005
R10973 D[6].n14 D[6].t1 34.0928
R10974 D[6].n11 D[6] 24.4785
R10975 D[6].n12 D[6].n11 21.9377
R10976 D[6].n11 D[6].n10 14.6672
R10977 D[6] D[6].n7 9.01934
R10978 D[6] D[6].n14 8.85188
R10979 D[6].n9 D[6] 7.57233
R10980 D[6].n7 D[6] 7.45876
R10981 D[6].n10 D[6] 3.24557
R10982 D[6].n13 D[6].n12 3.14374
R10983 D[6].n3 D[6] 3.01375
R10984 D[6].n12 D[6].n6 2.74043
R10985 D[6].n5 D[6].n1 2.26284
R10986 D[6].n4 D[6].n3 2.23869
R10987 D[6].n10 D[6].n9 1.44275
R10988 D[6].n14 D[6].n13 0.389863
R10989 D[6].n6 D[6].n0 0.0232273
R10990 D[6].n4 D[6].n2 0.00807576
R10991 D[6].n5 D[6].n4 0.00195195
R10992 D[6].n6 D[6].n5 0.00194159
R10993 sel_bit[0].n4 sel_bit[0].t2 445.048
R10994 sel_bit[0].n12 sel_bit[0].t0 432.193
R10995 sel_bit[0].n7 sel_bit[0].t4 287.995
R10996 sel_bit[0].n12 sel_bit[0].t3 254.389
R10997 sel_bit[0].n2 sel_bit[0].t1 252.248
R10998 sel_bit[0].n7 sel_bit[0].t5 194.809
R10999 sel_bit[0].n4 sel_bit[0].n3 152
R11000 sel_bit[0].n2 sel_bit[0].n1 152
R11001 sel_bit[0].n13 sel_bit[0].n12 76.0005
R11002 sel_bit[0].n8 sel_bit[0].n7 76.0005
R11003 sel_bit[0] sel_bit[0].n8 20.2672
R11004 sel_bit[0].n6 sel_bit[0].n5 15.6271
R11005 sel_bit[0].n5 sel_bit[0].n4 14.4605
R11006 sel_bit[0].n5 sel_bit[0].n2 12.8538
R11007 sel_bit[0].n14 sel_bit[0].n13 9.16815
R11008 sel_bit[0].n3 sel_bit[0] 9.03579
R11009 sel_bit[0].n13 sel_bit[0] 6.21226
R11010 sel_bit[0].n1 sel_bit[0] 5.64756
R11011 sel_bit[0].n10 sel_bit[0].n6 5.18664
R11012 sel_bit[0].n6 sel_bit[0].n0 4.88604
R11013 sel_bit[0].n9 sel_bit[0] 4.77729
R11014 sel_bit[0].n11 sel_bit[0] 4.25943
R11015 sel_bit[0].n8 sel_bit[0] 3.91161
R11016 sel_bit[0].n3 sel_bit[0].n0 3.01226
R11017 sel_bit[0].n1 sel_bit[0].n0 0.753441
R11018 sel_bit[0].n9 sel_bit[0] 0.563
R11019 sel_bit[0].n11 sel_bit[0] 0.259429
R11020 sel_bit[0].n10 sel_bit[0].n9 0.101633
R11021 sel_bit[0].n14 sel_bit[0].n11 0.0793043
R11022 sel_bit[0] sel_bit[0].n14 0.0793043
R11023 sel_bit[0] sel_bit[0].n10 0.0588664
R11024 clk_sar.n0 clk_sar.t0 259.031
R11025 clk_sar.n0 clk_sar.t1 175.778
R11026 clk_sar.n1 clk_sar.n0 8.08213
R11027 clk_sar.n1 clk_sar 4.54939
R11028 clk_sar clk_sar.n1 2.70993
R11029 comparator_out.n5 comparator_out.t1 255.085
R11030 comparator_out.n6 comparator_out.t0 174.536
R11031 comparator_out.n7 comparator_out.n6 9.3005
R11032 comparator_out.n6 comparator_out.n5 5.54501
R11033 comparator_out.n1 comparator_out 4.24368
R11034 comparator_out.n9 comparator_out.n8 2.76807
R11035 comparator_out.n7 comparator_out.n4 2.59138
R11036 comparator_out comparator_out.n9 1.55726
R11037 comparator_out.n3 comparator_out.n1 1.12138
R11038 comparator_out.n8 comparator_out.n7 0.173473
R11039 comparator_out.n1 comparator_out.n0 0.0114596
R11040 comparator_out.n4 comparator_out.n3 0.00870471
R11041 comparator_out.n3 comparator_out.n2 0.00290385
C0 x4.X a_10794_3239# 0.0425f
C1 a_7073_4801# a_6305_4112# 3.76e-19
C2 a_5845_4801# x45.Q_N 3.67e-20
C3 a_6760_4775# a_6845_4386# 7.46e-19
C4 a_2463_4775# a_3619_4801# 3.31e-19
C5 a_2289_4801# a_3453_4801# 6.38e-20
C6 a_6199_4801# a_5992_4086# 3.44e-19
C7 x4.X a_9872_3521# 0.00103f
C8 x30.Q_N x7.X 0.274f
C9 a_1415_4801# a_1616_4801# 3.67e-19
C10 a_1976_4775# x20.Q_N 0.0094f
C11 a_2463_4775# a_2697_5083# 0.00945f
C12 a_2289_4801# a_2194_4801# 0.00276f
C13 x33.Q_N a_8803_4112# 2.89e-22
C14 check[5] a_7049_2340# 7.15e-20
C15 x27.Q_N a_3618_3239# 3.65e-19
C16 check[6] x77.Y 3.89e-20
C17 a_7246_3213# a_8683_3605# 7.98e-21
C18 a_4453_2340# a_4657_2340# 0.117f
C19 a_4452_2640# a_4925_2550# 0.145f
C20 a_4154_2340# x54.Q_N 9.58e-21
C21 a_9639_4775# a_9464_3239# 1.33e-23
C22 a_6759_3213# a_9151_3213# 3.6e-20
C23 a_9465_4801# a_9638_3213# 4.82e-21
C24 a_8998_4801# a_9370_4801# 3.34e-19
C25 a_7072_3239# x72.Q_N 9.58e-21
C26 VDD a_5372_4112# 0.11f
C27 x4.X a_6985_4112# 6.8e-19
C28 x36.Q_N a_11183_3239# 6.74e-20
C29 a_6845_4386# a_9238_4086# 2.9e-21
C30 VDD x27.Q_N 0.452f
C31 a_3900_5167# a_3913_4112# 2.81e-19
C32 a_4074_4775# a_4155_4086# 8.83e-20
C33 a_3619_4801# a_4453_4386# 7.24e-20
C34 a_3453_4801# a_4454_4086# 1.15e-19
C35 x45.Q_N a_8384_4086# 5.27e-21
C36 a_4368_4775# a_3600_4086# 0.0018f
C37 x20.Q_N a_4155_4086# 2.32e-19
C38 check[0] a_6505_4394# 9.42e-20
C39 VDD x36.Q_N 0.419f
C40 a_6400_4801# check[5] 5.31e-21
C41 D[5] a_6845_2340# 1.11e-19
C42 a_8236_3239# a_10345_3239# 1.03e-19
C43 a_1112_2340# a_2060_2640# 7.7e-21
C44 D[7] a_1762_2340# 8.38e-19
C45 D[0] a_8791_3239# 1.27e-19
C46 x33.Q_N D[1] 3.29e-19
C47 check[4] a_11184_4801# 9.44e-20
C48 a_5170_4478# a_5372_4112# 8.94e-19
C49 x77.Y a_4317_3521# 4.28e-20
C50 a_4019_4112# a_4389_4112# 4.11e-20
C51 x4.X a_3900_5167# 0.00135f
C52 a_5992_4086# x7.X 0.00201f
C53 check[2] a_5845_4801# 1.76e-19
C54 VDD a_2533_2550# 0.194f
C55 x4.X a_11076_5167# 0.00135f
C56 comparator_out a_929_3238# 0.00685f
C57 check[2] a_11075_3605# 8.1e-20
C58 a_8289_4086# D[0] 0.00123f
C59 a_5089_5083# x27.Q_N 2.02e-20
C60 x39.Q_N a_11493_3521# 0.00136f
C61 a_10628_3239# a_11075_3605# 0.15f
C62 a_6844_2640# a_8696_2366# 1.79e-19
C63 a_7049_2340# a_7185_2366# 0.07f
C64 a_6845_2340# a_8383_2340# 0.00116f
C65 a_10794_3239# a_11249_3213# 0.153f
C66 x30.Q_N a_6605_3239# 6.1e-19
C67 check[1] a_8803_4112# 4.26e-19
C68 x69.Q_N a_10794_3239# 8.64e-20
C69 a_9872_3521# x69.Q_N 2.02e-20
C70 a_12265_5083# x36.Q_N 2.02e-20
C71 check[2] a_8384_4086# 6.25e-20
C72 x5.X a_7562_4478# 1.85e-19
C73 VDD a_11629_4386# 0.59f
C74 sel_bit[0] a_2788_5674# 3.68e-19
C75 x7.X a_3504_2340# 0.00285f
C76 VDD a_9151_3213# 0.353f
C77 check[2] a_11088_2366# 0.00327f
C78 check[0] a_4926_4296# 0.00111f
C79 check[4] a_10776_4086# 0.00416f
C80 eob x7.X 0.0869f
C81 x30.Q_N a_8288_2340# 2.02e-19
C82 a_9237_2340# a_9374_2732# 0.00907f
C83 D[4] a_9577_2366# 7.47e-20
C84 a_10628_3239# a_11088_2366# 1.89e-19
C85 a_10794_3239# a_10775_2340# 3.73e-19
C86 check[4] a_8402_3239# 1.83e-21
C87 x4.X a_7562_4112# 6.4e-19
C88 x4.A x7.X 1.17e-19
C89 a_6985_4112# a_7186_4112# 3.34e-19
C90 check[2] a_4855_4775# 2.07e-19
C91 a_8289_4086# a_8697_4112# 4.37e-19
C92 a_897_4112# a_1511_4112# 9.05e-20
C93 x4.X a_7246_3213# 0.115f
C94 VDD a_8938_2340# 0.177f
C95 a_5992_4086# a_6605_3239# 1.16e-20
C96 x45.Q_N a_6198_3239# 7.37e-20
C97 a_8237_4801# a_8858_4775# 0.117f
C98 x36.Q_N a_11331_4086# 1.3e-22
C99 a_10680_2340# a_11628_2640# 9.65e-21
C100 a_2061_2340# x51.Q_N 1.07e-19
C101 a_2265_2340# a_2533_2550# 0.205f
C102 a_10795_4801# a_11543_3213# 2.05e-21
C103 a_11250_4775# a_11075_3605# 1.33e-23
C104 a_11076_5167# a_11249_3213# 3.52e-21
C105 eob a_1207_2340# 7.14e-20
C106 a_4367_3213# a_4585_3239# 3.73e-19
C107 a_4680_3239# a_4213_3239# 0.00316f
C108 check[1] a_7481_5083# 4.45e-19
C109 VDD a_1976_4775# 0.489f
C110 a_1061_4801# a_897_4112# 0.00384f
C111 x4.X a_6844_2640# 0.00904f
C112 VDD a_12047_2648# 0.00984f
C113 x7.X D[2] 0.0211f
C114 x48.Q a_4318_5083# 4.61e-19
C115 a_4971_4801# a_4658_4086# 7.76e-20
C116 x4.A a_1207_2340# 7.71e-20
C117 x7.X x60.Q_N 3.61e-19
C118 a_4453_4386# a_3452_3239# 6.5e-20
C119 a_4155_4086# a_3618_3239# 1.07e-20
C120 x45.Q_N a_7049_2340# 1.11e-19
C121 a_3913_4112# a_4073_3213# 0.00148f
C122 a_6291_3605# D[0] 3.23e-21
C123 a_6759_3213# a_7953_3239# 6.04e-19
C124 VDD a_4155_4086# 0.348f
C125 VDD a_12048_4394# 0.00984f
C126 x4.X a_9953_2732# 1.17e-19
C127 x4.X a_12146_3239# 5.65e-19
C128 a_3453_4801# a_3807_4801# 0.0662f
C129 x4.X a_4073_3213# 0.00798f
C130 a_3619_4801# a_4681_4801# 0.137f
C131 a_3900_5167# a_4368_4775# 0.0633f
C132 x4.X a_11761_3239# 4.96e-19
C133 x30.Q_N a_6846_4086# 0.0258f
C134 a_11089_4112# a_11630_4086# 0.125f
C135 a_11331_4086# a_11629_4386# 0.137f
C136 a_9377_4112# x39.Q_N 2.88e-20
C137 x5.X a_9152_4775# 0.00142f
C138 a_2853_5648# a_3373_5674# 0.394f
C139 check[1] a_3258_5648# 0.0414f
C140 x45.Q_N a_4367_3213# 3.74e-20
C141 a_5845_4801# a_8591_4801# 3.65e-21
C142 a_6011_4801# a_6291_3605# 8.52e-21
C143 a_6292_5167# a_6010_3239# 1.65e-21
C144 a_6466_4775# a_6465_3213# 2.59e-19
C145 a_7073_4801# a_8403_4801# 4e-20
C146 a_6760_4775# a_5844_3239# 9.66e-21
C147 check[1] sel_bit[1] 0.26f
C148 x33.Q_N x39.Q_N 2.41e-20
C149 check[5] a_9237_2340# 7.28e-22
C150 D[0] a_6304_2366# 1.92e-21
C151 a_8683_3605# a_9151_3213# 0.0633f
C152 a_3912_2366# x57.Q_N 8.28e-21
C153 a_8402_3239# a_9464_3239# 0.137f
C154 a_8236_3239# a_8590_3239# 0.0708f
C155 a_4453_2340# a_6845_2340# 0.00176f
C156 x27.Q_N x75.Q_N 0.02f
C157 a_10795_4801# a_11857_4801# 0.137f
C158 x36.Q_N a_11194_2366# 0.0102f
C159 a_11076_5167# a_11544_4775# 0.0633f
C160 a_10629_4801# a_10983_4801# 0.0665f
C161 x48.Q_N a_4113_4394# 2.02e-20
C162 a_4453_4386# a_4872_4394# 2.46e-19
C163 a_3913_4112# a_5372_4112# 1.65e-21
C164 a_4658_4086# a_4591_4478# 9.46e-19
C165 a_929_3238# x7.X 0.225f
C166 x27.Q_N a_3913_4112# 1.32e-21
C167 a_8237_4801# x42.Q_N 3.67e-20
C168 a_9465_4801# a_8697_4112# 3.76e-19
C169 a_9152_4775# a_9237_4386# 7.46e-19
C170 a_7186_4112# a_7246_3213# 4.45e-20
C171 a_8591_4801# a_8384_4086# 3.44e-19
C172 a_3373_5674# a_3671_5674# 0.00489f
C173 a_6844_2640# D[4] 0.00557f
C174 a_6845_2340# a_7763_2366# 0.0708f
C175 a_7049_2340# a_7561_2732# 6.69e-20
C176 x36.Q_N a_11195_4112# 2.89e-22
C177 a_8683_3605# a_8938_2340# 2.41e-20
C178 a_8236_3239# a_9441_2340# 4.77e-19
C179 a_8402_3239# a_9237_2340# 6.38e-20
C180 a_9151_3213# a_8696_2366# 3.36e-20
C181 a_8857_3213# a_9236_2640# 2.68e-19
C182 a_4367_3213# a_4452_2640# 5.32e-19
C183 a_4680_3239# a_3912_2366# 2.17e-19
C184 a_8997_3239# D[1] 1.13e-20
C185 a_3806_3239# a_3599_2340# 2.02e-19
C186 x4.X a_5372_4112# 0.00623f
C187 x33.Q_N a_9709_2550# 0.181f
C188 a_5992_4086# a_6846_4086# 0.0492f
C189 a_6305_4112# a_6845_4386# 0.139f
C190 x4.X x27.Q_N 0.425f
C191 VDD a_7953_3239# 0.19f
C192 a_2853_5648# eob 0.00163f
C193 VDD a_4925_2550# 0.174f
C194 check[2] D[3] 0.194f
C195 x4.X x36.Q_N 0.278f
C196 a_929_3238# a_1207_2340# 0.00346f
C197 a_5845_4801# a_6931_5083# 0.00907f
C198 a_6011_4801# a_6710_5083# 2.46e-19
C199 a_10628_3239# D[3] 5.2e-19
C200 D[1] a_10680_2340# 0.00635f
C201 a_8288_2340# x60.Q_N 0.178f
C202 a_8383_2340# a_9236_2640# 0.0264f
C203 a_8696_2366# a_8938_2340# 0.124f
C204 a_9639_4775# a_10983_4801# 8.26e-21
C205 x33.Q_N a_11768_2366# 2.75e-20
C206 a_12030_3213# a_11942_3605# 7.71e-20
C207 a_11543_3213# a_11389_3239# 0.00943f
C208 a_11075_3605# a_11183_3239# 0.00812f
C209 a_11249_3213# a_11761_3239# 9.75e-19
C210 a_11856_3239# a_11714_3521# 0.00412f
C211 a_10628_3239# x66.Q_N 1.07e-19
C212 VDD a_5845_4801# 0.81f
C213 x4.X a_2533_2550# 5.96e-19
C214 VDD a_11075_3605# 0.176f
C215 a_4794_4112# a_3912_2366# 1.26e-20
C216 x39.Q_N a_9954_4112# 2.57e-20
C217 a_11630_4086# a_11767_4478# 0.00907f
C218 VDD a_12147_4801# 0.0101f
C219 check[2] check[4] 0.347f
C220 a_1520_2366# a_1996_2732# 0.00133f
C221 x27.Q_N a_4657_2340# 0.179f
C222 a_9709_2550# a_9953_2366# 0.00812f
C223 check[4] a_10628_3239# 0.00655f
C224 a_10629_4801# D[1] 1.99e-20
C225 a_3452_3239# a_5561_3239# 1.03e-19
C226 check[2] a_2883_5674# 0.0516f
C227 a_2389_5648# a_2969_6040# 0.00342f
C228 a_1338_5674# sel_bit[1] 0.0467f
C229 VDD a_8384_4086# 0.716f
C230 x5.X a_4591_4478# 1.55e-19
C231 check[1] a_9709_2550# 2.04e-19
C232 x4.X a_11629_4386# 0.0479f
C233 x4.X a_9151_3213# 0.111f
C234 a_9442_4086# x42.Q_N 0.00116f
C235 a_1508_5167# a_1976_4775# 0.0627f
C236 VDD a_11088_2366# 0.348f
C237 a_5089_5083# a_5845_4801# 4.06e-20
C238 a_2979_2366# a_2777_2366# 3.67e-19
C239 a_4074_4775# a_4367_3213# 7.57e-21
C240 x5.X a_11390_4801# 9.46e-19
C241 a_3453_4801# a_4680_3239# 4.76e-21
C242 a_3504_2340# a_3599_2340# 0.0968f
C243 a_1996_2366# a_2401_2366# 2.46e-21
C244 x20.Q_N a_1112_2340# 4.68e-19
C245 x20.Q_N a_4367_3213# 1.25e-21
C246 check[4] a_9376_2366# 9.3e-20
C247 a_2061_2340# x54.Q_N 2.94e-19
C248 a_7246_3213# a_7072_3239# 0.197f
C249 a_5844_3239# a_6709_3521# 0.00276f
C250 a_8403_4801# a_9370_4801# 0.00126f
C251 a_8237_4801# a_9873_5083# 1.25e-19
C252 a_9152_4775# a_9551_5167# 0.00133f
C253 a_8684_5167# a_8998_4801# 0.0258f
C254 a_6759_3213# a_6198_3239# 3.79e-20
C255 a_6291_3605# a_6375_3605# 0.00972f
C256 reset x3.A 0.00364f
C257 x36.Q_N a_11249_3213# 5.36e-19
C258 x48.Q a_2993_5674# 1.96e-19
C259 VDD a_4855_4775# 0.723f
C260 a_6305_4112# a_7264_4394# 1.21e-20
C261 a_6547_4086# a_6411_4112# 0.0282f
C262 a_6845_4386# a_6983_4478# 1.09e-19
C263 a_9442_4086# x7.X 4.39e-21
C264 x4.X a_8938_2340# 0.00706f
C265 x5.X a_7954_4801# 0.0293f
C266 VDD a_12031_4775# 0.709f
C267 x7.X a_12101_2550# 0.00818f
C268 a_6466_4775# check[5] 1.71e-20
C269 check[0] a_5562_4801# 0.0162f
C270 D[0] a_8857_3213# 8.87e-20
C271 a_7246_3213# a_6845_2340# 8.72e-19
C272 a_7072_3239# a_6844_2640# 1.11e-20
C273 check[1] a_4926_4296# 1.97e-22
C274 a_6759_3213# a_7049_2340# 0.00144f
C275 check[4] a_11250_4775# 6.31e-19
C276 x72.Q_N D[0] 2.5e-19
C277 x36.Q_N a_10775_2340# 0.142f
C278 a_1061_4801# a_1415_4801# 0.0708f
C279 x4.X a_1976_4775# 0.0979f
C280 a_1227_4801# a_2289_4801# 0.137f
C281 sel_bit[1] a_3453_4801# 0.00123f
C282 a_3505_4086# a_4454_4086# 1.03e-19
C283 a_3600_4086# a_4453_4386# 0.0264f
C284 a_3913_4112# a_4155_4086# 0.124f
C285 a_2883_5674# x20.Q_N 5.75e-20
C286 x4.X a_12047_2648# 2.86e-19
C287 check[2] a_11834_4086# 1.08e-19
C288 a_4368_4775# x27.Q_N 0.00773f
C289 a_3807_4801# a_4008_4801# 3.67e-19
C290 a_4855_4775# a_5089_5083# 0.00945f
C291 a_4681_4801# a_4586_4801# 0.00276f
C292 x5.X a_8236_3239# 9.93e-20
C293 check[6] a_4388_2366# 2.11e-20
C294 a_11834_4086# a_10628_3239# 0.00195f
C295 a_11630_4086# a_10794_3239# 6.04e-20
C296 a_11089_4112# a_11543_3213# 3.33e-20
C297 a_11331_4086# a_11075_3605# 1.7e-20
C298 a_11629_4386# a_11249_3213# 0.0015f
C299 D[0] a_8383_2340# 0.00127f
C300 x30.Q_N a_6010_3239# 4.02e-19
C301 a_5991_2340# x57.Q_N 0.124f
C302 a_9464_3239# a_10628_3239# 6.38e-20
C303 a_9151_3213# a_11249_3213# 4.53e-20
C304 a_6844_2640# a_6845_2340# 0.781f
C305 a_9638_3213# a_10794_3239# 1.69e-19
C306 a_6304_2366# a_7317_2550# 0.0633f
C307 a_6546_2340# a_7049_2340# 0.00187f
C308 a_4367_3213# a_6759_3213# 3.6e-20
C309 a_4854_3213# a_6291_3605# 7.98e-21
C310 a_9464_3239# a_9369_3239# 0.00276f
C311 a_9151_3213# x69.Q_N 0.00553f
C312 a_9638_3213# a_9872_3521# 0.00945f
C313 a_8590_3239# a_8791_3239# 3.67e-19
C314 a_1062_5674# a_1061_4801# 0.00165f
C315 x4.X a_4155_4086# 0.00873f
C316 a_11544_4775# x36.Q_N 0.0059f
C317 a_12031_4775# a_12265_5083# 0.00945f
C318 a_10983_4801# a_11184_4801# 3.67e-19
C319 a_11857_4801# a_11762_4801# 0.00276f
C320 VDD a_9173_4478# 0.00371f
C321 x4.X a_12048_4394# 8.47e-19
C322 a_4454_4086# x45.Q_N 3.85e-19
C323 a_9237_4386# a_9578_4112# 0.00118f
C324 VDD a_7182_4801# 7.87e-19
C325 a_8939_4086# a_10776_4086# 1.86e-21
C326 x42.Q_N a_10156_4112# 8.23e-20
C327 VDD a_6198_3239# 0.109f
C328 a_9238_4086# a_9377_4112# 2.56e-19
C329 check[2] a_9237_2340# 6.22e-19
C330 a_9237_4386# a_8236_3239# 6.5e-20
C331 x7.X x77.Y 0.00119f
C332 check[6] a_6199_4801# 0.165f
C333 a_8697_4112# a_8857_3213# 0.00148f
C334 a_8939_4086# a_8402_3239# 1.07e-20
C335 x33.Q_N a_9238_4086# 0.026f
C336 a_5561_3239# D[5] 0.00127f
C337 D[4] a_8938_2340# 1.94e-19
C338 a_9638_3213# a_9577_2366# 1.2e-20
C339 reset a_653_3238# 1.96e-19
C340 check[1] x27.D 1.12e-20
C341 eob a_1616_4801# 4.1e-19
C342 x33.Q_N a_11833_2340# 8.49e-21
C343 a_10156_4112# x7.X 5.5e-20
C344 check[0] a_3876_6040# 2.26e-19
C345 a_3170_4801# a_1511_4112# 5.42e-19
C346 x7.X a_4388_2732# 1.8e-19
C347 VDD a_7049_2340# 0.304f
C348 a_6305_4112# a_5844_3239# 2.21e-19
C349 a_5992_4086# a_6010_3239# 3.48e-19
C350 x48.Q_N a_3599_2340# 9.38e-21
C351 a_4453_4386# a_4453_2340# 7.25e-19
C352 a_4454_4086# a_4452_2640# 7.02e-19
C353 check[0] a_6305_4112# 0.00126f
C354 a_3600_4086# x54.Q_N 2.32e-20
C355 a_8697_4112# a_8383_2340# 5.05e-21
C356 a_9953_2732# a_10155_2366# 8.94e-19
C357 a_10983_4801# a_10776_4086# 3.44e-19
C358 a_11544_4775# a_11629_4386# 7.46e-19
C359 a_10629_4801# x39.Q_N 3.68e-20
C360 a_11857_4801# a_11089_4112# 3.76e-19
C361 a_9236_2640# a_9577_2366# 0.00118f
C362 a_9237_2340# a_9376_2366# 2.56e-19
C363 a_8938_2340# a_10775_2340# 1.86e-21
C364 a_8696_2366# a_11088_2366# 4.59e-21
C365 a_12146_3239# a_11965_3239# 4.11e-20
C366 a_3452_3239# a_4854_3213# 0.0492f
C367 a_4073_3213# a_3899_3605# 0.205f
C368 a_3618_3239# a_4367_3213# 0.139f
C369 check[1] a_6760_4775# 0.00254f
C370 x33.Q_N a_9755_4801# 3.78e-19
C371 a_1061_4801# a_3170_4801# 1.03e-19
C372 x5.A a_1338_5674# 0.3f
C373 a_1062_5674# a_2389_5648# 2.65e-20
C374 check[2] a_4454_4086# 2.36e-20
C375 x5.X a_1511_4112# 2.24e-19
C376 x4.X a_7953_3239# 0.00272f
C377 check[6] x7.X 0.0236f
C378 x4.X a_4925_2550# 0.00127f
C379 x5.X a_11289_4394# 4.41e-19
C380 VDD D[3] 0.221f
C381 VDD a_1112_2340# 0.226f
C382 VDD a_4367_3213# 0.356f
C383 VDD x66.Q_N 0.0716f
C384 a_4539_5083# check[6] 1.43e-21
C385 check[3] x7.X 0.0244f
C386 a_11195_4112# a_11075_3605# 1.12e-20
C387 x27.Q_N a_6845_2340# 6.49e-21
C388 a_11628_2640# a_11564_2732# 2.13e-19
C389 a_11629_2340# a_11288_2648# 1.25e-19
C390 a_11088_2366# a_11194_2366# 0.0552f
C391 a_11330_2340# a_11766_2732# 0.00412f
C392 x77.Y a_4018_2366# 6.03e-20
C393 check[1] a_9238_4086# 2.12e-19
C394 x5.X a_1061_4801# 0.265f
C395 a_11715_5083# check[3] 9.55e-19
C396 x4.X a_5845_4801# 0.00422f
C397 x5.X a_7318_4296# 6.4e-19
C398 x4.X a_11075_3605# 0.0178f
C399 a_7247_4775# a_6846_4086# 0.00169f
C400 a_2463_4775# a_3900_5167# 7.98e-21
C401 a_6466_4775# x45.Q_N 2.19e-19
C402 a_6760_4775# a_7050_4086# 0.00268f
C403 a_7073_4801# a_6845_4386# 1.96e-20
C404 VDD check[4] 0.5f
C405 x4.X a_12147_4801# 0.00557f
C406 a_2289_4801# x20.Q_N 8.79e-19
C407 a_8803_4112# a_8402_3239# 4.04e-21
C408 x27.Q_N a_6606_4801# 1.93e-20
C409 a_11195_4112# a_11088_2366# 8.38e-21
C410 x27.Q_N a_3899_3605# 0.00192f
C411 a_4855_4775# x75.Q_N 4.45e-20
C412 a_4453_2340# x54.Q_N 1.07e-19
C413 a_4657_2340# a_4925_2550# 0.205f
C414 VDD a_2883_5674# 0.172f
C415 x36.Q_N a_10155_2366# 1.34e-20
C416 a_8998_4801# x33.Q_N 4.01e-20
C417 VDD a_4389_4112# 9.51e-19
C418 x36.Q_N a_11965_3239# 1.68e-19
C419 x4.X a_8384_4086# 0.101f
C420 a_2389_5648# a_3170_4801# 1.39e-19
C421 a_4368_4775# a_4155_4086# 3.72e-19
C422 a_4855_4775# a_3913_4112# 0.00161f
C423 a_6547_4086# x42.Q_N 7.23e-21
C424 a_4074_4775# a_4454_4086# 0.00336f
C425 a_3619_4801# a_4658_4086# 0.00221f
C426 x4.X a_11088_2366# 0.112f
C427 x20.Q_N a_4454_4086# 1.21e-19
C428 check[0] a_6983_4478# 6.27e-20
C429 x48.Q check[0] 0.0102f
C430 x45.Q_N x75.Q 9.42e-21
C431 check[6] a_4018_2366# 1.17e-19
C432 a_7481_5083# check[5] 1.93e-21
C433 x30.Q_N a_7954_4801# 0.182f
C434 a_7953_3239# D[4] 0.00127f
C435 D[5] a_7317_2550# 1.96e-20
C436 a_8402_3239# D[1] 5.69e-21
C437 D[7] a_2061_2340# 1.85e-19
C438 a_1227_4801# a_3807_4801# 3.07e-21
C439 a_2389_5648# x5.X 0.00105f
C440 x4.X a_4855_4775# 0.102f
C441 sel_bit[0] a_2853_5648# 1.09f
C442 check[2] a_6466_4775# 1.08e-19
C443 sel_bit[1] x3.A 1.43e-20
C444 x4.X a_12031_4775# 0.0991f
C445 clk_sar reset 1.31e-20
C446 x30.Q_N a_8236_3239# 8.92e-20
C447 x39.Q_N a_11942_3605# 3.64e-19
C448 a_6845_2340# a_8938_2340# 6.38e-20
C449 a_7317_2550# a_8383_2340# 7.98e-21
C450 a_5561_3239# a_4453_2340# 4.83e-19
C451 a_10794_3239# a_11543_3213# 0.139f
C452 a_10628_3239# a_12030_3213# 0.0492f
C453 a_7049_2340# a_8696_2366# 8.4e-21
C454 a_11249_3213# a_11075_3605# 0.205f
C455 x30.Q_N a_6977_3239# 4.04e-19
C456 check[2] a_8939_4086# 5.79e-20
C457 x5.X a_8289_4086# 0.0767f
C458 VDD a_11834_4086# 0.487f
C459 x27.D a_3453_4801# 0.412f
C460 a_3170_4801# a_3619_4801# 6.24e-19
C461 VDD a_9464_3239# 0.18f
C462 check[2] a_11628_2640# 3.14e-19
C463 x42.Q_N a_9101_3521# 0.00136f
C464 x30.Q_N a_6984_2366# 0.00473f
C465 a_9237_2340# a_9655_2648# 0.00276f
C466 a_9236_2640# a_9953_2732# 4.45e-20
C467 a_8696_2366# D[3] 1.61e-20
C468 a_11249_3213# a_11088_2366# 0.0014f
C469 a_11075_3605# a_10775_2340# 3.9e-20
C470 a_10628_3239# a_11628_2640# 6.01e-20
C471 check[1] a_5562_4801# 3.76e-20
C472 x4.X a_9173_4478# 2.12e-19
C473 x5.X a_3619_4801# 0.0076f
C474 a_7764_4112# a_9238_4086# 3.65e-21
C475 a_8289_4086# a_9237_4386# 9.65e-21
C476 x5.X a_2697_5083# 3.53e-19
C477 x4.X a_6198_3239# 0.00604f
C478 x7.X a_6504_2648# 1.52e-19
C479 x4.X a_7182_4801# 2.39e-19
C480 VDD a_9237_2340# 0.784f
C481 a_4368_4775# a_5845_4801# 1.72e-19
C482 x5.X a_10795_4801# 0.0203f
C483 x45.Q_N a_4970_3239# 9.58e-21
C484 a_1520_2366# a_1996_2366# 2.87e-21
C485 D[3] a_11194_2366# 5.39e-19
C486 a_8237_4801# a_9152_4775# 0.125f
C487 a_8403_4801# a_8684_5167# 0.155f
C488 a_10775_2340# a_11088_2366# 0.273f
C489 check[4] a_8696_2366# 1.1e-20
C490 x36.Q_N a_11630_4086# 0.0255f
C491 a_11857_4801# a_10794_3239# 6.75e-21
C492 x77.Y a_3599_2340# 2.75e-19
C493 a_11544_4775# a_12147_4801# 0.0552f
C494 a_4367_3213# x75.Q_N 0.00553f
C495 eob a_1762_2340# 2.19e-19
C496 a_4854_3213# a_5088_3521# 0.00945f
C497 a_4680_3239# a_4585_3239# 0.00276f
C498 a_3806_3239# a_4007_3239# 3.67e-19
C499 VDD a_2289_4801# 0.203f
C500 x48.Q a_4389_4478# 3.17e-19
C501 check[6] a_6846_4086# 2.07e-22
C502 VDD a_12547_2366# 0.109f
C503 x4.X a_7049_2340# 0.00149f
C504 x48.Q a_4767_5167# 1.31e-19
C505 x4.A a_1762_2340# 3.45e-19
C506 a_4454_4086# a_3618_3239# 6.04e-20
C507 a_3913_4112# a_4367_3213# 3.33e-20
C508 a_4658_4086# a_3452_3239# 0.00195f
C509 a_4453_4386# a_4073_3213# 0.0015f
C510 a_4155_4086# a_3899_3605# 1.7e-20
C511 a_3599_2340# a_4388_2732# 7.71e-20
C512 a_3912_2366# a_4112_2648# 0.00185f
C513 a_5844_3239# a_5896_2340# 4.5e-19
C514 a_7246_3213# D[0] 0.0116f
C515 check[0] a_5896_2340# 0.028f
C516 a_4970_3239# a_4452_2640# 5.05e-21
C517 VDD a_4454_4086# 0.809f
C518 x36.Q_N a_9236_2640# 0.00112f
C519 check[2] a_8803_4112# 1.27e-20
C520 VDD a_12548_4112# 0.109f
C521 x4.X a_6400_4801# 8.46e-20
C522 x4.X D[3] 5.34e-19
C523 x4.X a_1112_2340# 0.0104f
C524 a_4074_4775# a_3807_4801# 6.99e-20
C525 a_3619_4801# a_3984_5167# 4.45e-20
C526 a_4368_4775# a_4855_4775# 0.273f
C527 x4.X a_4367_3213# 0.112f
C528 x5.X a_9465_4801# 0.00117f
C529 x4.X x66.Q_N 0.00462f
C530 x20.Q_N a_3807_4801# 1.92e-19
C531 check[2] a_9323_5083# 4.69e-19
C532 a_11089_4112# a_12102_4296# 0.0633f
C533 a_10776_4086# x39.Q_N 0.155f
C534 a_11629_4386# a_11630_4086# 0.782f
C535 a_11331_4086# a_11834_4086# 0.00187f
C536 x30.Q_N a_7318_4296# 5.71e-19
C537 x45.Q_N a_4680_3239# 1.74e-21
C538 check[6] a_3599_2340# 2.38e-20
C539 a_6466_4775# a_6759_3213# 7.57e-21
C540 a_5845_4801# a_7072_3239# 4.76e-21
C541 check[1] a_6305_4112# 0.00312f
C542 D[0] a_6844_2640# 6.76e-19
C543 a_7953_3239# a_6845_2340# 4.83e-19
C544 a_4452_2640# x57.Q_N 1.53e-19
C545 a_8857_3213# a_8590_3239# 6.99e-20
C546 a_9151_3213# a_9638_3213# 0.273f
C547 a_8402_3239# a_8767_3605# 4.45e-20
C548 a_11250_4775# a_10983_4801# 6.99e-20
C549 sel_bit[1] a_3505_4086# 1.09e-19
C550 a_11544_4775# a_12031_4775# 0.273f
C551 a_10795_4801# a_11160_5167# 4.45e-20
C552 a_4454_4086# a_5170_4478# 0.0018f
C553 a_4453_4386# a_5372_4112# 0.162f
C554 a_4658_4086# a_4872_4394# 0.0104f
C555 a_3913_4112# a_4389_4112# 2.87e-21
C556 a_8384_4086# a_8897_4394# 0.00945f
C557 x4.X check[4] 0.037f
C558 comparator_out x7.X 0.0433f
C559 x27.Q_N a_4453_4386# 0.0318f
C560 check[2] D[1] 0.171f
C561 a_9465_4801# a_9237_4386# 1.96e-20
C562 a_9639_4775# a_9238_4086# 0.00169f
C563 a_8858_4775# x42.Q_N 2.19e-19
C564 a_9152_4775# a_9442_4086# 0.00268f
C565 a_7317_2550# a_7763_2366# 0.0367f
C566 a_10345_3239# a_10794_3239# 3.74e-19
C567 D[1] a_10628_3239# 0.348f
C568 sel_bit[1] a_1227_4801# 3.53e-20
C569 x75.Q a_6759_3213# 9.18e-20
C570 a_9151_3213# a_9236_2640# 5.32e-19
C571 a_9464_3239# a_8696_2366# 2.17e-19
C572 a_8590_3239# a_8383_2340# 2.02e-19
C573 a_9369_3239# D[1] 1.36e-20
C574 a_4680_3239# a_4452_2640# 1.11e-20
C575 a_4367_3213# a_4657_2340# 0.00144f
C576 a_4854_3213# a_4453_2340# 8.72e-19
C577 x4.X a_4389_4112# 3.84e-19
C578 a_6305_4112# a_7050_4086# 0.199f
C579 a_5992_4086# a_7318_4296# 4.7e-22
C580 a_6547_4086# a_6846_4086# 0.0334f
C581 a_4794_4112# x45.Q_N 5.94e-20
C582 x5.X a_6710_5083# 3.44e-19
C583 a_6466_4775# a_6931_5083# 9.46e-19
C584 a_6011_4801# a_7159_5167# 2.13e-19
C585 x5.X a_3452_3239# 3.24e-20
C586 a_5845_4801# a_6606_4801# 6.04e-20
C587 check[0] a_4318_5083# 1.54e-19
C588 eob a_1511_4112# 0.0585f
C589 a_8938_2340# a_9236_2640# 0.137f
C590 a_11543_3213# a_12146_3239# 0.0552f
C591 a_8696_2366# a_9237_2340# 0.125f
C592 a_9639_4775# a_9755_4801# 0.0397f
C593 a_9152_4775# a_9574_4801# 2.87e-21
C594 a_11856_3239# a_11389_3239# 0.00316f
C595 a_11543_3213# a_11761_3239# 3.73e-19
C596 VDD a_6466_4775# 0.488f
C597 x4.A a_1511_4112# 0.619f
C598 a_3453_4801# a_5562_4801# 1.03e-19
C599 VDD a_12030_3213# 0.568f
C600 VDD reset 0.161f
C601 a_11089_4112# a_11565_4112# 2.87e-21
C602 a_11629_4386# a_12346_4478# 4.45e-20
C603 eob a_1061_4801# 0.514f
C604 a_11630_4086# a_12048_4394# 0.00276f
C605 a_7954_4801# a_8237_4801# 8.18e-19
C606 a_2061_2340# a_1720_2648# 1.25e-19
C607 x42.Q_N a_9573_3239# 7.87e-19
C608 a_1520_2366# a_1626_2366# 0.0552f
C609 a_1762_2340# a_2198_2732# 0.00412f
C610 a_2060_2640# a_1996_2732# 2.13e-19
C611 x27.Q_N x54.Q_N 4.08e-19
C612 check[1] a_6983_4478# 9.03e-21
C613 D[3] a_10775_2340# 0.0131f
C614 a_10155_2366# a_11088_2366# 3.42e-20
C615 x30.Q_N a_9172_2366# 1.14e-20
C616 check[2] a_3258_5648# 0.0201f
C617 check[1] x48.Q 0.0512f
C618 a_2389_5648# a_3373_5674# 0.176f
C619 x77.Y a_6010_3239# 0.00188f
C620 a_10629_4801# a_12738_4801# 9.94e-20
C621 check[4] x69.Q_N 0.00316f
C622 a_1061_4801# x4.A 0.00353f
C623 check[2] sel_bit[1] 0.393f
C624 x5.X a_4872_4394# 1.11e-19
C625 VDD a_8939_4086# 0.34f
C626 clk_sar sel_bit[1] 0.329f
C627 x4.X a_11834_4086# 0.00986f
C628 a_5845_4801# a_5897_4086# 6.04e-19
C629 a_1976_4775# a_2463_4775# 0.271f
C630 a_6199_4801# x7.X 1.97e-20
C631 VDD x75.Q 0.216f
C632 x4.X a_9464_3239# 0.00475f
C633 VDD a_11628_2640# 0.269f
C634 x27.Q_N a_6011_4801# 1.48e-19
C635 x5.X a_11762_4801# 2.61e-19
C636 a_4368_4775# a_4367_3213# 0.00121f
C637 a_8237_4801# a_8236_3239# 6.9e-19
C638 a_8403_4801# x33.Q_N 2.97e-20
C639 a_7363_4801# a_7182_4801# 4.11e-20
C640 a_9465_4801# a_9551_5167# 0.00976f
C641 check[4] a_10775_2340# 7.18e-21
C642 a_6465_3213# a_6709_3521# 0.0104f
C643 a_6010_3239# a_6930_3521# 1.09e-19
C644 x77.Y a_4793_2366# 5.33e-22
C645 x48.Q a_3877_5674# 4.02e-19
C646 x36.Q_N a_11543_3213# 0.00494f
C647 VDD a_3807_4801# 0.117f
C648 x36.Q_N a_11966_4801# 7.29e-21
C649 a_6845_4386# a_7264_4394# 2.46e-19
C650 x45.Q_N a_6505_4394# 2.02e-20
C651 a_6305_4112# a_7764_4112# 1.65e-21
C652 a_7050_4086# a_6983_4478# 9.46e-19
C653 x42.Q_N x7.X 0.00133f
C654 x4.X a_9237_2340# 0.00274f
C655 VDD a_10983_4801# 0.109f
C656 a_6760_4775# check[5] 0.00406f
C657 a_7247_4775# a_7954_4801# 0.0968f
C658 check[6] a_6010_3239# 9.27e-20
C659 a_4018_2366# a_4388_2366# 4.11e-20
C660 a_2389_5648# eob 0.222f
C661 x27.Q_N a_5561_3239# 0.00748f
C662 D[0] a_9151_3213# 1.24e-19
C663 a_7246_3213# a_7317_2550# 1.66e-21
C664 a_7072_3239# a_7049_2340# 1.03e-19
C665 check[4] a_11544_4775# 0.00302f
C666 x36.Q_N a_11330_2340# 0.16f
C667 x4.X a_2289_4801# 0.167f
C668 a_1061_4801# a_1926_5083# 0.00276f
C669 a_1227_4801# a_1592_5167# 4.45e-20
C670 a_1682_4775# a_1415_4801# 6.99e-20
C671 sel_bit[1] x20.Q_N 3.57e-20
C672 a_4155_4086# a_4453_4386# 0.137f
C673 a_3913_4112# a_4454_4086# 0.125f
C674 x5.X a_11089_4112# 0.00571f
C675 check[2] x39.Q_N 0.0223f
C676 x4.X a_12547_2366# 5.99e-20
C677 a_4681_4801# x27.Q_N 5.04e-19
C678 x5.X D[5] 3.43e-19
C679 check[5] a_9238_4086# 6.24e-22
C680 check[6] a_4793_2366# 4.42e-19
C681 a_11629_4386# a_11543_3213# 5.72e-19
C682 a_11089_4112# a_11856_3239# 2.16e-19
C683 a_10776_4086# a_10982_3239# 2.44e-19
C684 x39.Q_N a_10628_3239# 0.0434f
C685 a_6606_4801# a_7182_4801# 2.46e-21
C686 x30.Q_N a_6291_3605# 0.00193f
C687 a_9151_3213# a_11543_3213# 3.6e-20
C688 a_6845_2340# a_7049_2340# 0.117f
C689 a_6844_2640# a_7317_2550# 0.145f
C690 a_6546_2340# x57.Q_N 9.58e-21
C691 a_9638_3213# a_11075_3605# 7.98e-21
C692 x4.X a_4454_4086# 0.0468f
C693 x33.Q_N a_9754_3239# 0.00342f
C694 a_9464_3239# x69.Q_N 9.58e-21
C695 x5.A a_1227_4801# 6.27e-21
C696 a_11857_4801# x36.Q_N 8.57e-20
C697 check[1] a_8403_4801# 0.00119f
C698 VDD a_8803_4112# 0.00996f
C699 x4.X a_12548_4112# 0.00434f
C700 a_4926_4296# x45.Q_N 1.43e-19
C701 VDD a_4970_3239# 0.00144f
C702 VDD a_9323_5083# 0.0163f
C703 a_9238_4086# a_10776_4086# 2.98e-19
C704 a_9442_4086# a_9578_4112# 0.07f
C705 x42.Q_N a_9173_4112# 0.00139f
C706 x7.X a_1207_2340# 8.03e-19
C707 a_9237_4386# a_11089_4112# 9.95e-20
C708 check[6] a_4971_4801# 8.4e-20
C709 a_9238_4086# a_8402_3239# 6.04e-20
C710 a_8697_4112# a_9151_3213# 3.33e-20
C711 a_9237_4386# a_8857_3213# 0.0015f
C712 a_8939_4086# a_8683_3605# 1.7e-20
C713 a_9442_4086# a_8236_3239# 0.00195f
C714 a_11089_4112# a_11629_2340# 1.4e-21
C715 a_11331_4086# a_11628_2640# 4.75e-21
C716 x33.Q_N a_9710_4296# 5.71e-19
C717 D[4] a_9237_2340# 1.09e-19
C718 eob a_3619_4801# 9.05e-22
C719 x30.Q_N a_6304_2366# 0.0928f
C720 a_10628_3239# a_12737_3239# 1.03e-19
C721 check[5] a_9755_4801# 1.85e-20
C722 a_4214_4801# x77.Y 1.91e-20
C723 eob a_2697_5083# 4.29e-19
C724 D[1] a_11183_3239# 1.22e-19
C725 x33.Q_N x63.Q_N 7.78e-20
C726 x27.D a_3505_4086# 5.09e-21
C727 VDD D[1] 0.3f
C728 VDD x57.Q_N 0.0716f
C729 check[0] a_6845_4386# 1.56e-19
C730 check[2] a_11768_2366# 3.3e-19
C731 a_6547_4086# a_6010_3239# 1.07e-20
C732 a_6305_4112# a_6465_3213# 0.00148f
C733 a_6845_4386# a_5844_3239# 6.5e-20
C734 a_4926_4296# a_4452_2640# 6.02e-22
C735 a_4453_4386# a_4925_2550# 6.45e-21
C736 a_12031_4775# a_11630_4086# 0.00169f
C737 a_11250_4775# x39.Q_N 2.02e-19
C738 a_11857_4801# a_11629_4386# 1.96e-20
C739 a_11544_4775# a_11834_4086# 0.00268f
C740 x30.Q_N a_8802_2366# 9.32e-20
C741 a_9441_2340# a_9577_2366# 0.07f
C742 a_9236_2640# a_11088_2366# 1.89e-19
C743 a_9237_2340# a_10775_2340# 0.00116f
C744 a_3618_3239# a_4680_3239# 0.137f
C745 a_3452_3239# a_3806_3239# 0.0662f
C746 check[1] a_7073_4801# 0.00111f
C747 a_3899_3605# a_4367_3213# 0.0632f
C748 a_1227_4801# x27.D 4.24e-20
C749 a_12264_3521# x66.Q_N 2.02e-20
C750 check[2] a_4926_4296# 2.18e-22
C751 x5.A check[2] 6.94e-20
C752 x5.X a_3600_4086# 1.13e-19
C753 clk_sar x5.A 0.00353f
C754 check[2] a_11769_4112# 3.17e-20
C755 x5.X a_11767_4478# 4e-19
C756 x48.Q a_3453_4801# 0.0505f
C757 VDD a_7481_5083# 0.00506f
C758 VDD a_4680_3239# 0.183f
C759 x7.X a_8288_2340# 7.84e-19
C760 a_6305_4112# a_5991_2340# 5.05e-21
C761 D[6] a_1996_2366# 3.71e-20
C762 check[5] a_8998_4801# 2.15e-19
C763 a_11629_2340# a_11766_2732# 0.00907f
C764 check[4] a_10155_2366# 0.00335f
C765 check[1] a_9710_4296# 3.53e-20
C766 x5.X a_1682_4775# 0.00288f
C767 x75.Q_N x75.Q 2.81e-20
C768 a_11390_4801# check[3] 1.02e-20
C769 x4.X a_6466_4775# 9.39e-19
C770 x4.X a_12030_3213# 0.116f
C771 a_6760_4775# x45.Q_N 9.66e-21
C772 a_7247_4775# a_7318_4296# 2.97e-21
C773 a_7073_4801# a_7050_4086# 2.59e-19
C774 a_9710_4296# a_9954_4112# 0.00812f
C775 a_5372_4112# a_4854_3213# 2.07e-19
C776 a_8803_4112# a_8683_3605# 1.12e-20
C777 x27.Q_N a_6978_4801# 1.15e-20
C778 a_3912_2366# a_5896_2340# 1.34e-20
C779 VDD a_3258_5648# 0.116f
C780 a_3599_2340# a_4388_2366# 4.2e-20
C781 x27.Q_N a_4854_3213# 0.0125f
C782 a_7953_3239# D[0] 0.0968f
C783 a_10346_4801# check[4] 0.13f
C784 VDD sel_bit[1] 0.38f
C785 a_7246_3213# a_8590_3239# 8.26e-21
C786 a_9370_4801# x33.Q_N 4.03e-20
C787 VDD a_4794_4112# 0.0336f
C788 x4.X a_8939_4086# 0.00731f
C789 check[2] x27.D 1.63e-20
C790 a_4368_4775# a_4454_4086# 4.63e-19
C791 a_4855_4775# a_4453_4386# 6.17e-19
C792 a_6846_4086# x42.Q_N 2.42e-19
C793 x4.X x75.Q 8.71e-19
C794 x4.X a_11628_2640# 0.00712f
C795 a_8237_4801# a_8289_4086# 6.04e-19
C796 a_6411_4112# a_6010_3239# 4.04e-21
C797 x5.X a_4453_2340# 2.59e-20
C798 check[0] a_7264_4394# 1.47e-20
C799 a_8803_4112# a_8696_2366# 8.38e-21
C800 a_3452_3239# a_3504_2340# 4.5e-19
C801 a_2784_5996# a_2883_5674# 0.00134f
C802 a_9151_3213# a_10345_3239# 6.04e-19
C803 a_8683_3605# D[1] 3.23e-21
C804 a_1112_2340# x51.Q_N 0.178f
C805 D[7] a_2533_2550# 6.45e-20
C806 eob a_3452_3239# 3.51e-19
C807 x4.X a_3807_4801# 2.51e-19
C808 a_6846_4086# x7.X 3.21e-20
C809 check[2] a_6760_4775# 1.3e-19
C810 x4.X a_10983_4801# 2.36e-19
C811 check[2] a_10982_3239# 0.00707f
C812 a_5845_4801# a_6011_4801# 0.751f
C813 sel_bit[0] a_1511_4112# 3.42e-19
C814 x20.Q_N a_1996_2732# 3.64e-19
C815 a_8237_4801# a_10795_4801# 2.9e-21
C816 a_8403_4801# a_10629_4801# 4e-20
C817 x30.Q_N D[5] 0.00272f
C818 D[1] a_8696_2366# 1.64e-21
C819 a_10628_3239# a_10982_3239# 0.0708f
C820 x30.Q_N x72.Q_N 0.0201f
C821 a_6845_2340# a_9237_2340# 0.00176f
C822 a_11075_3605# a_11543_3213# 0.0633f
C823 a_6304_2366# x60.Q_N 5.09e-21
C824 a_10794_3239# a_11856_3239# 0.137f
C825 a_12147_4801# a_11543_3213# 1.05e-20
C826 a_12147_4801# a_11966_4801# 4.11e-20
C827 VDD x39.Q_N 0.458f
C828 check[2] a_9238_4086# 0.439f
C829 sel_bit[0] a_1061_4801# 4.66e-20
C830 check[5] a_6305_4112# 7.68e-22
C831 x27.D a_4074_4775# 6.07e-19
C832 VDD a_8767_3605# 0.0042f
C833 x7.X a_3599_2340# 0.00328f
C834 x20.Q_N x27.D 0.0032f
C835 x48.Q a_4790_4801# 6.64e-20
C836 check[2] a_11833_2340# 4.61e-19
C837 check[4] a_11630_4086# 1.46e-21
C838 x42.Q_N a_9550_3605# 3.64e-19
C839 a_9236_2640# D[3] 0.00531f
C840 x30.Q_N a_8383_2340# 1.64e-19
C841 check[4] a_9638_3213# 0.00527f
C842 a_9237_2340# a_10155_2366# 0.0708f
C843 a_9441_2340# a_9953_2732# 6.69e-20
C844 a_11543_3213# a_11088_2366# 3.36e-20
C845 a_11249_3213# a_11628_2640# 2.68e-19
C846 a_10628_3239# a_11833_2340# 4.77e-19
C847 a_11075_3605# a_11330_2340# 2.41e-20
C848 a_10794_3239# a_11629_2340# 6.38e-20
C849 a_11389_3239# D[2] 1.3e-20
C850 VDD a_6505_4394# 0.00506f
C851 x4.X a_8803_4112# 0.00332f
C852 check[2] a_2579_4801# 1.13e-21
C853 a_8384_4086# a_8697_4112# 0.272f
C854 x5.X a_3900_5167# 1.6e-19
C855 x4.X a_4970_3239# 5.69e-19
C856 VDD a_12737_3239# 0.189f
C857 x7.X a_6982_2732# 9.43e-19
C858 VDD a_9709_2550# 0.172f
C859 a_4855_4775# a_6011_4801# 1.83e-19
C860 a_4681_4801# a_5845_4801# 6.38e-20
C861 x5.X a_11076_5167# 0.00471f
C862 x45.Q_N a_6709_3521# 0.00136f
C863 a_1626_2366# D[6] 3.23e-20
C864 a_8237_4801# a_9465_4801# 0.0334f
C865 a_8403_4801# a_9639_4775# 0.0264f
C866 a_8858_4775# a_9152_4775# 0.199f
C867 check[3] a_11289_4394# 1.21e-21
C868 a_1520_2366# a_2401_2366# 0.00943f
C869 check[0] a_5844_3239# 0.051f
C870 a_1762_2340# a_2200_2366# 0.00276f
C871 a_2061_2340# a_3504_2340# 8.18e-19
C872 x36.Q_N a_12102_4296# 1.85e-19
C873 a_12031_4775# a_11543_3213# 1.08e-22
C874 check[4] a_9236_2640# 0.0285f
C875 a_11544_4775# a_12030_3213# 1.06e-20
C876 a_10775_2340# a_11628_2640# 0.0264f
C877 a_10680_2340# x63.Q_N 0.178f
C878 a_11088_2366# a_11330_2340# 0.124f
C879 x77.Y a_4154_2340# 0.00178f
C880 a_12031_4775# a_11966_4801# 4.2e-20
C881 a_11857_4801# a_12147_4801# 0.0282f
C882 a_5372_4112# a_5170_4112# 3.67e-19
C883 eob a_2061_2340# 0.00216f
C884 a_4680_3239# x75.Q_N 9.58e-21
C885 VDD a_1592_5167# 0.00558f
C886 x4.X D[1] 0.0011f
C887 VDD a_11768_2366# 6.2e-19
C888 x4.X x57.Q_N 0.00786f
C889 x48.Q a_4008_4801# 3.94e-19
C890 a_2389_5648# sel_bit[0] 0.137f
C891 a_4453_4386# a_4367_3213# 5.72e-19
C892 a_3600_4086# a_3806_3239# 2.44e-19
C893 a_3913_4112# a_4680_3239# 2.16e-19
C894 a_4855_4775# a_5561_3239# 4.94e-20
C895 a_4154_2340# a_4388_2732# 0.00976f
C896 a_3912_2366# a_4590_2732# 0.00652f
C897 a_3599_2340# a_4018_2366# 0.0397f
C898 a_4970_3239# a_4657_2340# 3.49e-20
C899 VDD x5.A 0.181f
C900 VDD a_4926_4296# 0.319f
C901 sel_bit[1] a_1508_5167# 5.1e-20
C902 a_2883_5674# a_2463_4775# 6.31e-19
C903 VDD a_11769_4112# 0.00445f
C904 x4.X a_4680_3239# 0.0059f
C905 a_3900_5167# a_3984_5167# 0.00972f
C906 a_4855_4775# a_4681_4801# 0.197f
C907 a_3453_4801# a_4318_5083# 0.00276f
C908 a_11331_4086# x39.Q_N 0.029f
C909 a_11630_4086# a_11834_4086# 0.117f
C910 x5.X a_8768_5167# 4.18e-19
C911 a_11629_4386# a_12102_4296# 0.155f
C912 x20.Q_N a_2579_4801# 0.00429f
C913 check[6] a_4154_2340# 1.2e-19
C914 a_5371_2366# a_5169_2366# 3.67e-19
C915 a_7247_4775# a_9465_4801# 1.86e-21
C916 a_6760_4775# a_6759_3213# 0.00121f
C917 a_5896_2340# a_5991_2340# 0.0968f
C918 a_4388_2366# a_4793_2366# 2.46e-21
C919 check[1] a_6845_4386# 0.163f
C920 a_3373_5674# a_3600_4086# 2.25e-20
C921 a_9638_3213# a_9464_3239# 0.197f
C922 a_9151_3213# a_8590_3239# 3.79e-20
C923 a_8236_3239# a_9101_3521# 0.00276f
C924 a_8683_3605# a_8767_3605# 0.00972f
C925 a_11544_4775# a_10983_4801# 3.29e-21
C926 a_11076_5167# a_11160_5167# 0.00972f
C927 a_12031_4775# a_11857_4801# 0.197f
C928 a_10629_4801# a_11494_5083# 0.00276f
C929 x36.Q_N a_11564_2366# 9.42e-19
C930 a_4926_4296# a_5170_4478# 0.00972f
C931 a_3913_4112# a_4794_4112# 0.00943f
C932 a_4454_4086# a_5897_4086# 3.23e-19
C933 a_4155_4086# a_4593_4112# 0.00276f
C934 a_4658_4086# a_5372_4112# 6.99e-20
C935 VDD a_1996_2732# 0.00483f
C936 a_8697_4112# a_9173_4478# 0.00133f
C937 check[2] a_5562_4801# 4.53e-20
C938 a_9465_4801# a_9442_4086# 2.59e-19
C939 a_9639_4775# a_9710_4296# 2.97e-21
C940 a_9152_4775# x42.Q_N 9.8e-21
C941 sel_bit[0] a_3619_4801# 8.15e-19
C942 a_10681_4086# a_10680_2340# 1.07e-20
C943 a_3619_4801# x77.Y 5.26e-21
C944 a_3258_5648# x4.X 3.57e-21
C945 x30.Q_N a_4453_2340# 1.57e-19
C946 sel_bit[1] x4.X 2.14e-19
C947 D[1] a_11249_3213# 8.77e-20
C948 a_9151_3213# a_9441_2340# 0.00144f
C949 a_9464_3239# a_9236_2640# 1.11e-20
C950 a_9638_3213# a_9237_2340# 8.72e-19
C951 x69.Q_N D[1] 2.5e-19
C952 a_4680_3239# a_4657_2340# 1.03e-19
C953 x4.X a_4794_4112# 0.00375f
C954 a_4854_3213# a_4925_2550# 1.66e-21
C955 VDD x27.D 0.294f
C956 a_6305_4112# x45.Q_N 0.093f
C957 a_6845_4386# a_7050_4086# 0.153f
C958 x7.X a_6010_3239# 0.149f
C959 x7.X a_2979_2366# 0.157f
C960 a_3600_4086# a_3504_2340# 2.97e-20
C961 x5.X a_7159_5167# 1.05e-19
C962 a_6011_4801# a_6400_4801# 0.0019f
C963 a_6466_4775# a_6606_4801# 0.07f
C964 a_10629_4801# a_10681_4086# 6.04e-19
C965 a_5845_4801# a_6978_4801# 2.56e-19
C966 a_6760_4775# a_6931_5083# 0.00652f
C967 x39.Q_N a_11194_2366# 5e-20
C968 check[0] a_4767_5167# 1.92e-19
C969 eob a_3600_4086# 4.72e-22
C970 x30.Q_N a_7763_2366# 0.0318f
C971 D[1] a_10775_2340# 0.00122f
C972 a_8938_2340# a_9441_2340# 0.00187f
C973 a_12030_3213# a_11965_3239# 4.2e-20
C974 a_9236_2640# a_9237_2340# 0.781f
C975 a_9465_4801# a_9574_4801# 0.00707f
C976 a_8383_2340# x60.Q_N 0.124f
C977 a_11856_3239# a_12146_3239# 0.0282f
C978 a_8696_2366# a_9709_2550# 0.0633f
C979 a_11856_3239# a_11761_3239# 0.00276f
C980 a_10982_3239# a_11183_3239# 3.67e-19
C981 a_12030_3213# a_12264_3521# 0.00945f
C982 a_11543_3213# x66.Q_N 0.00553f
C983 VDD a_6760_4775# 0.449f
C984 a_3619_4801# check[6] 5.82e-21
C985 VDD a_10982_3239# 0.109f
C986 x39.Q_N a_11195_4112# 0.0451f
C987 a_11834_4086# a_12346_4478# 6.69e-20
C988 a_11630_4086# a_12548_4112# 0.0708f
C989 a_11331_4086# a_11769_4112# 0.00276f
C990 a_11089_4112# a_11970_4112# 0.00943f
C991 eob a_1682_4775# 0.0484f
C992 check[5] a_8403_4801# 0.162f
C993 a_2061_2340# a_2198_2732# 0.00907f
C994 check[1] a_7264_4394# 6.91e-21
C995 check[4] a_11543_3213# 8.39e-21
C996 D[3] a_11330_2340# 1.99e-19
C997 a_2389_5648# a_2788_5674# 2.97e-20
C998 a_4367_3213# a_5561_3239# 6.04e-19
C999 a_10795_4801# check[3] 8.42e-19
C1000 check[4] a_11966_4801# 9.01e-21
C1001 a_1682_4775# x4.A 0.00205f
C1002 x5.X a_5372_4112# 9.6e-19
C1003 VDD a_9238_4086# 0.805f
C1004 check[2] a_6305_4112# 1.74e-20
C1005 x4.X x39.Q_N 0.253f
C1006 x48.Q a_3505_4086# 0.0868f
C1007 x4.X a_8767_3605# 9.07e-19
C1008 a_1508_5167# a_1592_5167# 0.00972f
C1009 VDD a_11833_2340# 0.304f
C1010 a_2463_4775# a_2289_4801# 0.197f
C1011 x5.X x27.Q_N 0.00103f
C1012 x7.X a_9172_2732# 1.81e-19
C1013 x27.Q_N a_6292_5167# 5.48e-20
C1014 x45.Q_N a_7181_3239# 7.87e-19
C1015 check[4] a_8697_4112# 3.77e-22
C1016 x5.X x36.Q_N 0.00489f
C1017 a_4855_4775# a_4854_3213# 0.00237f
C1018 a_8403_4801# a_8402_3239# 1.39e-19
C1019 a_3504_2340# a_4453_2340# 1.03e-19
C1020 a_12345_2732# a_12547_2366# 8.94e-19
C1021 a_6759_3213# a_6709_3521# 1.21e-20
C1022 a_6198_3239# a_6375_3605# 8.94e-19
C1023 a_9152_4775# a_9873_5083# 0.00185f
C1024 a_8684_5167# x33.Q_N 1.74e-20
C1025 a_6010_3239# a_6605_3239# 0.00118f
C1026 x4.X a_6505_4394# 1.75e-19
C1027 x36.Q_N a_11856_3239# 0.00293f
C1028 x48.Q a_1227_4801# 5.44e-21
C1029 a_6305_4112# a_6781_4112# 2.87e-21
C1030 a_6845_4386# a_7764_4112# 0.162f
C1031 a_7050_4086# a_7264_4394# 0.0104f
C1032 a_6846_4086# a_7562_4478# 0.0018f
C1033 VDD a_2579_4801# 0.0073f
C1034 x4.X a_12737_3239# 0.00277f
C1035 x4.X a_9709_2550# 0.00146f
C1036 VDD a_9755_4801# 0.0101f
C1037 a_5897_4086# x75.Q 0.00123f
C1038 a_7073_4801# check[5] 6.72e-20
C1039 a_4452_2640# a_5169_2366# 0.00105f
C1040 check[0] a_6780_2366# 1.28e-19
C1041 D[0] a_9464_3239# 3.72e-20
C1042 check[4] a_11857_4801# 4.17e-20
C1043 x77.Y a_3452_3239# 0.51f
C1044 x36.Q_N a_11629_2340# 0.0468f
C1045 a_1682_4775# a_1926_5083# 0.0104f
C1046 a_1227_4801# a_2147_5083# 1.09e-19
C1047 a_3600_4086# x48.Q_N 0.124f
C1048 a_3913_4112# a_4926_4296# 0.0633f
C1049 a_4453_4386# a_4454_4086# 0.75f
C1050 a_4155_4086# a_4658_4086# 0.00187f
C1051 x5.X a_11629_4386# 0.00326f
C1052 a_12346_4478# a_12548_4112# 8.94e-19
C1053 check[6] a_6304_2366# 2.39e-20
C1054 a_11834_4086# a_11543_3213# 0.0014f
C1055 x39.Q_N a_11249_3213# 0.194f
C1056 a_11630_4086# a_12030_3213# 7.94e-19
C1057 x30.Q_N a_7246_3213# 0.0127f
C1058 a_7247_4775# x72.Q_N 4.45e-20
C1059 a_12147_4801# a_12102_4296# 1.9e-20
C1060 D[0] a_9237_2340# 1.09e-20
C1061 a_6845_2340# x57.Q_N 1.07e-19
C1062 a_4854_3213# a_6198_3239# 8.26e-21
C1063 a_7049_2340# a_7317_2550# 0.205f
C1064 x4.X a_4926_4296# 0.0211f
C1065 check[1] a_5844_3239# 2.07e-22
C1066 VDD a_9954_4478# 0.0042f
C1067 check[1] check[0] 0.0116f
C1068 x4.X a_11769_4112# 6.71e-19
C1069 VDD a_4112_2648# 0.00555f
C1070 check[2] x48.Q 0.0879f
C1071 VDD a_6709_3521# 0.00984f
C1072 VDD a_8998_4801# 0.0332f
C1073 a_1508_5167# x27.D 4.66e-22
C1074 x7.X a_1762_2340# 1.88e-19
C1075 a_9238_4086# a_11331_4086# 1.67e-21
C1076 a_9710_4296# a_10776_4086# 7.98e-21
C1077 a_1976_4775# a_3170_4801# 6.04e-19
C1078 x42.Q_N a_9578_4112# 0.00172f
C1079 a_9237_4386# a_9151_3213# 5.72e-19
C1080 a_8384_4086# a_8590_3239# 2.44e-19
C1081 x42.Q_N a_8236_3239# 0.0435f
C1082 a_8697_4112# a_9464_3239# 2.16e-19
C1083 check[6] a_6710_5083# 2.57e-21
C1084 x20.Q_N a_1996_2366# 7.87e-19
C1085 check[6] a_3452_3239# 1.79e-20
C1086 a_11630_4086# a_11628_2640# 7.02e-19
C1087 a_10776_4086# x63.Q_N 2.32e-20
C1088 x39.Q_N a_10775_2340# 2.2e-19
C1089 a_11629_4386# a_11629_2340# 7.25e-19
C1090 x30.Q_N a_6844_2640# 0.57f
C1091 a_10345_3239# D[3] 0.00127f
C1092 D[1] a_11965_3239# 1.23e-20
C1093 D[4] a_9709_2550# 1.83e-20
C1094 a_10794_3239# D[2] 5.71e-21
C1095 x4.X a_1996_2732# 4.32e-19
C1096 VDD a_5562_4801# 0.192f
C1097 check[0] a_3877_5674# 0.00787f
C1098 x5.X a_1976_4775# 0.00314f
C1099 x7.X a_5169_2732# 8.25e-19
C1100 x7.X a_8236_3239# 0.147f
C1101 VDD a_12738_4801# 0.177f
C1102 a_6845_4386# a_6465_3213# 0.0015f
C1103 a_6547_4086# a_6291_3605# 1.7e-20
C1104 a_6305_4112# a_6759_3213# 3.33e-20
C1105 a_6846_4086# a_6010_3239# 6.04e-20
C1106 a_7050_4086# a_5844_3239# 0.00195f
C1107 check[2] a_12345_2366# 2.05e-20
C1108 check[0] a_7050_4086# 1.2e-19
C1109 a_4658_4086# a_4925_2550# 2.22e-22
C1110 a_8697_4112# a_9237_2340# 1.4e-21
C1111 a_8939_4086# a_9236_2640# 4.75e-21
C1112 a_11544_4775# x39.Q_N 9.93e-21
C1113 a_11857_4801# a_11834_4086# 2.59e-19
C1114 x27.Q_N a_4789_3239# 1.68e-19
C1115 a_12031_4775# a_12102_4296# 2.97e-21
C1116 a_1207_2340# a_1762_2340# 0.197f
C1117 check[4] a_10345_3239# 0.0274f
C1118 a_9709_2550# a_10775_2340# 7.98e-21
C1119 a_9237_2340# a_11330_2340# 6.38e-20
C1120 a_9441_2340# a_11088_2366# 7.2e-21
C1121 a_1112_2340# D[7] 0.0786f
C1122 a_3618_3239# a_3983_3605# 4.45e-20
C1123 a_4073_3213# a_3806_3239# 6.99e-20
C1124 a_4367_3213# a_4854_3213# 0.273f
C1125 a_3452_3239# a_4317_3521# 0.00276f
C1126 x4.X x27.D 0.00252f
C1127 x5.X a_4155_4086# 7.39e-20
C1128 x48.Q a_4074_4775# 0.00395f
C1129 x5.X a_12048_4394# 1.32e-19
C1130 VDD a_3983_3605# 0.00494f
C1131 x48.Q x20.Q_N 0.0441f
C1132 a_2979_2366# a_3599_2340# 8.26e-21
C1133 a_2533_2550# a_2777_2366# 0.00812f
C1134 D[6] a_2401_2366# 5.27e-19
C1135 check[5] a_9370_4801# 7.95e-20
C1136 check[0] a_3912_2366# 2.06e-21
C1137 a_11629_2340# a_12047_2648# 0.00276f
C1138 a_11088_2366# a_11564_2366# 2.87e-21
C1139 a_11628_2640# a_12345_2732# 4.45e-20
C1140 a_11762_4801# check[3] 7.79e-21
C1141 x4.X a_6760_4775# 0.104f
C1142 x4.X a_10982_3239# 0.00531f
C1143 x7.X a_11288_2648# 1.53e-19
C1144 a_2463_4775# a_3807_4801# 8.26e-21
C1145 check[2] a_8403_4801# 4.08e-19
C1146 a_10681_4086# a_10776_4086# 0.0968f
C1147 a_9173_4112# a_9578_4112# 2.46e-21
C1148 a_4454_4086# a_5561_3239# 4.72e-19
C1149 a_1822_4801# a_2194_4801# 3.34e-19
C1150 x27.Q_N x30.Q_N 2.3e-20
C1151 check[0] a_6410_2366# 0.00226f
C1152 a_4452_2640# a_5896_2340# 6.96e-19
C1153 a_4154_2340# a_4388_2366# 0.00707f
C1154 VDD a_3876_6040# 0.00865f
C1155 a_3912_2366# a_4592_2366# 3.73e-19
C1156 a_7246_3213# a_7362_3239# 0.0397f
C1157 a_6759_3213# a_7181_3239# 2.87e-21
C1158 a_6605_3239# a_6977_3239# 3.34e-19
C1159 VDD a_6305_4112# 0.448f
C1160 a_1511_4112# x7.X 8.67e-19
C1161 x4.X a_9238_4086# 0.0468f
C1162 a_7318_4296# x42.Q_N 8.46e-20
C1163 a_4855_4775# a_4658_4086# 4.44e-19
C1164 a_4368_4775# a_4926_4296# 2.85e-19
C1165 x4.X a_11833_2340# 0.00145f
C1166 x5.X a_7953_3239# 0.00125f
C1167 a_6411_4112# a_6291_3605# 1.12e-20
C1168 check[6] D[5] 0.141f
C1169 a_5991_2340# a_6780_2732# 7.71e-20
C1170 a_6304_2366# a_6504_2648# 0.00185f
C1171 check[3] a_11089_4112# 0.0033f
C1172 a_9638_3213# D[1] 0.0115f
C1173 a_8236_3239# a_8288_2340# 4.5e-19
C1174 a_7362_3239# a_6844_2640# 5.05e-21
C1175 a_2883_5674# a_2969_6040# 0.0136f
C1176 x77.Y a_5088_3521# 8.16e-21
C1177 a_5372_4112# a_5992_4086# 8.26e-21
C1178 x4.X a_2579_4801# 0.0171f
C1179 VDD a_1996_2366# 4.24e-19
C1180 check[2] a_7073_4801# 4.32e-20
C1181 x5.X a_5845_4801# 0.27f
C1182 x4.X a_9755_4801# 0.00557f
C1183 a_1511_4112# a_1207_2340# 1.58e-19
C1184 a_6411_4112# a_6304_2366# 8.38e-21
C1185 a_6011_4801# a_6466_4775# 0.153f
C1186 sel_bit[0] a_3600_4086# 3.59e-19
C1187 a_5845_4801# a_6292_5167# 0.15f
C1188 x20.Q_N a_1626_2366# 0.00967f
C1189 a_3600_4086# x77.Y 1.36e-19
C1190 check[0] a_3453_4801# 0.00279f
C1191 x5.X a_12147_4801# 2.09e-19
C1192 x39.Q_N a_11965_3239# 7.87e-19
C1193 x30.Q_N a_9151_3213# 8.28e-21
C1194 x33.Q_N a_9953_2366# 0.00224f
C1195 x39.Q_N a_12264_3521# 2.75e-19
C1196 a_11249_3213# a_10982_3239# 6.99e-20
C1197 a_10345_3239# a_9237_2340# 4.83e-19
C1198 a_11543_3213# a_12030_3213# 0.273f
C1199 a_10794_3239# a_11159_3605# 4.45e-20
C1200 D[1] a_9236_2640# 5.41e-19
C1201 check[1] a_9377_4112# 3.4e-20
C1202 a_6844_2640# x60.Q_N 1.38e-19
C1203 check[1] x33.Q_N 0.0011f
C1204 check[2] a_9710_4296# 0.00118f
C1205 x5.X a_8384_4086# 0.0202f
C1206 VDD a_5169_2366# 4e-20
C1207 sel_bit[0] a_1682_4775# 3.83e-20
C1208 x27.D a_4368_4775# 0.00307f
C1209 check[5] a_6845_4386# 0.0306f
C1210 x7.X a_4154_2340# 0.00109f
C1211 a_7954_4801# a_6846_4086# 6.67e-19
C1212 check[2] x63.Q_N 0.0121f
C1213 x48.Q a_3618_3239# 2.51e-19
C1214 x27.Q_N a_3504_2340# 3.7e-19
C1215 x30.Q_N a_8938_2340# 5.93e-20
C1216 D[2] a_12146_3239# 9.48e-20
C1217 a_9709_2550# a_10155_2366# 0.0367f
C1218 a_10982_3239# a_10775_2340# 2.02e-19
C1219 a_11761_3239# D[2] 1.36e-20
C1220 a_11856_3239# a_11088_2366# 2.17e-19
C1221 a_11543_3213# a_11628_2640# 5.32e-19
C1222 VDD a_6983_4478# 0.0163f
C1223 x4.X a_9954_4478# 9.15e-19
C1224 VDD x48.Q 0.638f
C1225 x4.X a_4112_2648# 0.00102f
C1226 a_8289_4086# x42.Q_N 0.18f
C1227 x5.X a_4855_4775# 0.00928f
C1228 a_8697_4112# a_8939_4086# 0.124f
C1229 a_8384_4086# a_9237_4386# 0.0264f
C1230 x4.X a_8998_4801# 7.25e-19
C1231 x4.X a_6709_3521# 2.91e-19
C1232 x7.X a_7263_2648# 6.92e-19
C1233 a_4855_4775# a_6292_5167# 7.98e-21
C1234 x5.X a_12031_4775# 0.00483f
C1235 x45.Q_N a_7158_3605# 3.63e-19
C1236 a_5844_3239# a_6465_3213# 0.117f
C1237 a_8684_5167# a_9639_4775# 4.7e-22
C1238 a_8237_4801# a_8768_5167# 0.0018f
C1239 a_8403_4801# a_8591_4801# 0.162f
C1240 a_1520_2366# a_3912_2366# 6.12e-21
C1241 a_2060_2640# a_2401_2366# 0.00118f
C1242 a_2061_2340# a_2200_2366# 2.56e-19
C1243 a_1762_2340# a_3599_2340# 1.86e-21
C1244 a_8858_4775# a_9465_4801# 0.00187f
C1245 D[3] a_11564_2366# 3.38e-20
C1246 a_5561_3239# x75.Q 0.0955f
C1247 check[4] a_9441_2340# 7.03e-20
C1248 x77.Y a_4453_2340# 3.65e-20
C1249 a_12031_4775# a_11856_3239# 1.33e-23
C1250 a_11088_2366# a_11629_2340# 0.125f
C1251 a_11330_2340# a_11628_2640# 0.137f
C1252 a_11857_4801# a_12030_3213# 4.82e-21
C1253 check[1] a_9953_2366# 2.06e-20
C1254 eob a_2533_2550# 4.21e-20
C1255 a_8289_4086# x7.X 2.05e-21
C1256 x4.X a_5562_4801# 0.00612f
C1257 x48.Q a_5170_4478# 5.12e-20
C1258 VDD a_2147_5083# 0.0199f
C1259 x4.X a_12738_4801# 0.00262f
C1260 x48.Q a_5089_5083# 1.17e-19
C1261 a_4658_4086# a_4367_3213# 0.0014f
C1262 a_4454_4086# a_4854_3213# 7.94e-19
C1263 a_4452_2640# a_4590_2732# 1.09e-19
C1264 D[6] a_4592_2366# 3.35e-19
C1265 a_4154_2340# a_4018_2366# 0.0282f
C1266 a_3912_2366# a_4871_2648# 1.21e-20
C1267 a_2853_5648# a_1511_4112# 6.37e-19
C1268 a_5844_3239# a_5991_2340# 8.35e-19
C1269 check[0] a_5991_2340# 0.0146f
C1270 check[1] a_9954_4112# 5.77e-22
C1271 x36.Q_N D[2] 0.00122f
C1272 sel_bit[1] a_2463_4775# 5.3e-20
C1273 check[2] a_10681_4086# 0.126f
C1274 x5.X a_9173_4478# 3.15e-19
C1275 x4.X a_3983_3605# 0.00103f
C1276 a_4074_4775# a_4318_5083# 0.0104f
C1277 a_3619_4801# a_4539_5083# 1.09e-19
C1278 a_10795_4801# x7.X 2.89e-21
C1279 x5.X a_7182_4801# 5.34e-20
C1280 a_11630_4086# x39.Q_N 0.00117f
C1281 a_11834_4086# a_12102_4296# 0.205f
C1282 a_10681_4086# a_10628_3239# 5.06e-19
C1283 check[6] a_4453_2340# 0.0409f
C1284 x39.Q_N a_9638_3213# 3.76e-21
C1285 a_7247_4775# a_7246_3213# 0.00237f
C1286 a_6760_4775# a_7363_4801# 0.0552f
C1287 check[1] a_7050_4086# 7.72e-19
C1288 a_8857_3213# a_9101_3521# 0.0104f
C1289 a_8402_3239# a_9322_3521# 1.09e-19
C1290 x33.Q_N a_8997_3239# 6.08e-19
C1291 a_11250_4775# a_11494_5083# 0.0104f
C1292 x36.Q_N a_11969_2366# 0.0403f
C1293 a_10795_4801# a_11715_5083# 1.09e-19
C1294 a_4453_4386# a_4794_4112# 0.00118f
C1295 a_4155_4086# a_5992_4086# 1.86e-21
C1296 a_4454_4086# a_4593_4112# 2.56e-19
C1297 VDD a_1626_2366# 0.00785f
C1298 a_8939_4086# a_9375_4478# 0.00412f
C1299 a_8697_4112# a_8803_4112# 0.051f
C1300 a_9238_4086# a_8897_4394# 1.25e-19
C1301 VDD a_8403_4801# 0.593f
C1302 a_9237_4386# a_9173_4478# 2.13e-19
C1303 a_11630_4086# a_12737_3239# 4.72e-19
C1304 sel_bit[0] a_3900_5167# 2.68e-19
C1305 a_3900_5167# x77.Y 7.98e-21
C1306 a_6410_2366# a_6780_2366# 4.11e-20
C1307 x30.Q_N a_7953_3239# 0.00834f
C1308 reset a_897_4112# 0.00119f
C1309 a_621_4112# x3.A 0.129f
C1310 D[1] a_11543_3213# 1.24e-19
C1311 a_9464_3239# a_9441_2340# 1.03e-19
C1312 x33.Q_N a_10680_2340# 1.87e-19
C1313 a_9638_3213# a_9709_2550# 1.66e-21
C1314 eob a_1976_4775# 0.0525f
C1315 check[3] a_10794_3239# 1.56e-21
C1316 x4.X a_6305_4112# 0.11f
C1317 a_6845_4386# x45.Q_N 0.00117f
C1318 a_6846_4086# a_7318_4296# 0.15f
C1319 VDD a_5896_2340# 0.189f
C1320 x7.X a_6291_3605# 0.00113f
C1321 check[0] a_4019_4112# 1.03e-20
C1322 x5.X D[3] 3.43e-19
C1323 x5.X a_6400_4801# 2.84e-19
C1324 a_8289_4086# a_8288_2340# 1.07e-20
C1325 a_7247_4775# a_7159_5167# 7.71e-20
C1326 a_6292_5167# a_6400_4801# 0.00812f
C1327 a_6760_4775# a_6606_4801# 0.00943f
C1328 a_5845_4801# x30.Q_N 2.24e-19
C1329 a_7073_4801# a_6931_5083# 0.00412f
C1330 a_6466_4775# a_6978_4801# 9.75e-19
C1331 a_2389_5648# a_2853_5648# 0.202f
C1332 a_8938_2340# x60.Q_N 9.58e-21
C1333 a_9237_2340# a_9441_2340# 0.117f
C1334 a_9236_2640# a_9709_2550# 0.145f
C1335 x33.Q_N a_10629_4801# 7.17e-19
C1336 a_11856_3239# x66.Q_N 9.58e-21
C1337 VDD a_7073_4801# 0.343f
C1338 VDD a_9754_3239# 4.88e-19
C1339 a_3900_5167# check[6] 1.4e-21
C1340 x7.X a_6304_2366# 0.00689f
C1341 a_4368_4775# a_5562_4801# 6.04e-19
C1342 a_11630_4086# a_11769_4112# 2.56e-19
C1343 a_12102_4296# a_12548_4112# 0.0367f
C1344 x42.Q_N a_8802_2366# 4.74e-20
C1345 a_11629_4386# a_11970_4112# 0.00118f
C1346 x5.X check[4] 0.167f
C1347 a_2060_2640# a_2777_2732# 4.45e-20
C1348 check[5] a_8684_5167# 0.00124f
C1349 check[5] a_5844_3239# 1.81e-20
C1350 a_1520_2366# D[6] 6.36e-20
C1351 a_2061_2340# a_2479_2648# 0.00276f
C1352 check[1] a_7764_4112# 0.165f
C1353 D[3] a_11629_2340# 1.1e-19
C1354 a_12146_3239# a_12101_2550# 1.01e-20
C1355 check[2] a_2993_5674# 0.0021f
C1356 a_4854_3213# x75.Q 0.0108f
C1357 a_11076_5167# check[3] 5.35e-19
C1358 a_11544_4775# a_12738_4801# 6.04e-19
C1359 check[2] a_6845_4386# 1.41e-20
C1360 VDD a_9710_4296# 0.317f
C1361 x48.Q a_3913_4112# 8.72e-19
C1362 a_5845_4801# a_5992_4086# 0.00159f
C1363 x4.X a_7181_3239# 1.05e-19
C1364 VDD x63.Q_N 0.0716f
C1365 a_1976_4775# a_1926_5083# 1.21e-20
C1366 x7.X a_3452_3239# 6.64e-19
C1367 a_10346_4801# a_9238_4086# 6.67e-19
C1368 check[4] a_9237_4386# 0.028f
C1369 a_8684_5167# a_8402_3239# 1.65e-21
C1370 a_8858_4775# a_8857_3213# 2.59e-19
C1371 a_9152_4775# a_8236_3239# 9.66e-21
C1372 a_5844_3239# a_8402_3239# 2.9e-21
C1373 a_3599_2340# a_4154_2340# 0.197f
C1374 a_6010_3239# a_8236_3239# 4e-20
C1375 a_8403_4801# a_8683_3605# 8.52e-21
C1376 a_6010_3239# a_6977_3239# 0.00126f
C1377 a_9639_4775# x33.Q_N 0.126f
C1378 a_5844_3239# a_7480_3521# 1.25e-19
C1379 a_621_4112# a_653_3238# 6.51e-19
C1380 a_6759_3213# a_7158_3605# 0.00133f
C1381 check[1] a_3453_4801# 9.29e-20
C1382 a_6291_3605# a_6605_3239# 0.0258f
C1383 a_2853_5648# a_3619_4801# 3.82e-19
C1384 check[4] a_11629_2340# 1.57e-21
C1385 x4.X a_6983_4478# 0.00114f
C1386 x48.Q x4.X 0.188f
C1387 VDD a_4318_5083# 0.0104f
C1388 a_7050_4086# a_7764_4112# 6.99e-20
C1389 a_6547_4086# a_6985_4112# 0.00276f
C1390 a_7318_4296# a_7562_4478# 0.00972f
C1391 a_6305_4112# a_7186_4112# 0.00943f
C1392 a_6846_4086# a_8289_4086# 3.23e-19
C1393 VDD a_11494_5083# 0.00984f
C1394 a_4453_2340# a_6504_2648# 4.06e-20
C1395 check[0] a_7185_2366# 4.21e-19
C1396 x77.Y a_4073_3213# 0.201f
C1397 x36.Q_N a_12101_2550# 0.181f
C1398 a_1227_4801# a_1822_4801# 0.00118f
C1399 a_4454_4086# a_4658_4086# 0.117f
C1400 a_4453_4386# a_4926_4296# 0.155f
C1401 a_4155_4086# x48.Q_N 9.58e-21
C1402 x5.X a_11834_4086# 3.65e-19
C1403 a_12102_4296# a_12030_3213# 3.74e-20
C1404 a_11834_4086# a_11856_3239# 4.33e-20
C1405 x39.Q_N a_11543_3213# 0.0983f
C1406 a_6304_2366# a_8288_2340# 8.55e-21
C1407 a_10345_3239# D[1] 0.0968f
C1408 a_5991_2340# a_6780_2366# 4.2e-20
C1409 x30.Q_N a_7182_4801# 7.02e-20
C1410 a_9638_3213# a_10982_3239# 8.26e-21
C1411 a_4367_3213# a_4789_3239# 2.87e-21
C1412 a_4854_3213# a_4970_3239# 0.0397f
C1413 VDD a_10681_4086# 0.189f
C1414 x4.X a_12346_4112# 6.38e-19
C1415 VDD a_4590_2732# 0.0172f
C1416 a_1511_4112# a_2979_2366# 3.09e-20
C1417 x7.X a_2061_2340# 0.188f
C1418 VDD a_7158_3605# 0.00371f
C1419 VDD a_9370_4801# 0.00445f
C1420 a_8697_4112# x39.Q_N 1.05e-20
C1421 a_9238_4086# a_11630_4086# 1.37e-19
C1422 a_2463_4775# x27.D 0.00431f
C1423 x5.X a_9237_2340# 2.59e-20
C1424 x42.Q_N a_8857_3213# 0.194f
C1425 a_9442_4086# a_9151_3213# 0.0014f
C1426 a_9238_4086# a_9638_3213# 7.94e-19
C1427 x20.Q_N a_2401_2366# 0.0313f
C1428 x39.Q_N a_11330_2340# 0.0018f
C1429 a_12102_4296# a_11628_2640# 6.02e-22
C1430 a_11629_4386# a_12101_2550# 6.45e-21
C1431 x27.Q_N x77.Y 0.00357f
C1432 a_11543_3213# a_12737_3239# 6.04e-19
C1433 x30.Q_N a_7049_2340# 0.179f
C1434 a_11075_3605# D[2] 3.24e-21
C1435 x4.X a_1626_2366# 3.78e-20
C1436 a_11089_4112# x7.X 2.29e-20
C1437 x4.X a_8403_4801# 0.005f
C1438 x5.X a_2289_4801# 0.00166f
C1439 x7.X D[5] 0.00123f
C1440 x7.X a_8857_3213# 4.83e-19
C1441 a_5992_4086# a_6198_3239# 2.44e-19
C1442 x45.Q_N a_5844_3239# 0.0434f
C1443 a_6305_4112# a_7072_3239# 2.16e-19
C1444 a_6845_4386# a_6759_3213# 5.72e-19
C1445 x7.X x72.Q_N 1.49e-19
C1446 check[0] x45.Q_N 0.0173f
C1447 a_9238_4086# a_9236_2640# 7.02e-19
C1448 a_8384_4086# x60.Q_N 2.32e-20
C1449 x42.Q_N a_8383_2340# 2.17e-19
C1450 a_9237_4386# a_9237_2340# 7.25e-19
C1451 a_1207_2340# a_2061_2340# 0.0492f
C1452 a_1520_2366# a_2060_2640# 0.139f
C1453 a_6400_4801# x30.Q_N 3.71e-20
C1454 D[2] a_11088_2366# 5.92e-20
C1455 a_8696_2366# x63.Q_N 4.29e-21
C1456 a_9237_2340# a_11629_2340# 0.00176f
C1457 a_3899_3605# a_3983_3605# 0.00972f
C1458 a_4073_3213# a_4317_3521# 0.0104f
C1459 a_3618_3239# a_4538_3521# 1.09e-19
C1460 a_4854_3213# a_4680_3239# 0.197f
C1461 x33.Q_N a_11184_4801# 3.99e-20
C1462 x5.X a_4454_4086# 0.258f
C1463 sel_bit[1] a_897_4112# 1.46e-20
C1464 check[6] a_5372_4112# 0.00256f
C1465 x4.X a_5896_2340# 0.00507f
C1466 x48.Q a_4368_4775# 0.0017f
C1467 x5.X a_12548_4112# 5.39e-19
C1468 x7.X a_8383_2340# 0.00434f
C1469 a_6547_4086# a_6844_2640# 4.75e-21
C1470 a_6305_4112# a_6845_2340# 1.4e-21
C1471 VDD a_4538_3521# 0.0174f
C1472 x27.Q_N check[6] 0.934f
C1473 clk_sar a_621_4112# 9.27e-21
C1474 D[6] a_3912_2366# 0.00221f
C1475 a_11330_2340# a_11768_2366# 0.00276f
C1476 a_11833_2340# a_12345_2732# 6.69e-20
C1477 a_11088_2366# a_11969_2366# 0.00943f
C1478 check[5] x33.Q_N 3.66e-21
C1479 a_11629_2340# a_12547_2366# 0.0708f
C1480 check[0] a_4452_2640# 2.1e-19
C1481 x36.Q_N check[3] 1.17f
C1482 x4.X a_7073_4801# 0.00316f
C1483 x4.X a_9754_3239# 5.61e-19
C1484 x7.X a_11766_2732# 9.47e-19
C1485 check[2] a_8684_5167# 1.92e-19
C1486 a_1976_4775# a_2398_4801# 2.87e-21
C1487 a_2463_4775# a_2579_4801# 0.0397f
C1488 check[2] check[0] 0.872f
C1489 a_1822_4801# x20.Q_N 1.36e-19
C1490 a_4794_4112# a_4854_3213# 4.45e-20
C1491 a_5845_4801# a_8237_4801# 0.00176f
C1492 a_6465_3213# a_6410_2366# 5.71e-21
C1493 a_11970_4112# a_11088_2366# 1.26e-20
C1494 check[5] a_6780_2366# 2.23e-20
C1495 a_3912_2366# a_5991_2340# 1.15e-20
C1496 a_4154_2340# a_4793_2366# 0.00316f
C1497 a_4452_2640# a_4592_2366# 0.00126f
C1498 VDD a_2993_5674# 4.34e-19
C1499 a_7072_3239# a_7181_3239# 0.00707f
C1500 x33.Q_N a_8402_3239# 3.88e-19
C1501 VDD a_6845_4386# 0.59f
C1502 a_3600_4086# a_4113_4394# 0.00945f
C1503 x4.X a_9710_4296# 0.021f
C1504 a_3600_4086# x7.X 4.69e-20
C1505 a_4681_4801# a_4926_4296# 3.59e-20
C1506 x4.X x63.Q_N 0.00782f
C1507 a_8237_4801# a_8384_4086# 0.00159f
C1508 check[0] a_6781_4112# 9.63e-22
C1509 a_7247_4775# a_7953_3239# 4.94e-20
C1510 a_3648_5972# a_3258_5648# 8.72e-19
C1511 sel_bit[0] a_1976_4775# 1.72e-19
C1512 a_6304_2366# a_6982_2732# 0.00652f
C1513 a_5991_2340# a_6410_2366# 0.0397f
C1514 a_6546_2340# a_6780_2732# 0.00976f
C1515 check[3] a_11629_4386# 0.138f
C1516 a_2883_5674# a_3373_5674# 4.47e-19
C1517 a_12031_4775# a_11970_4112# 1.79e-20
C1518 a_12738_4801# a_11630_4086# 6.67e-19
C1519 a_3452_3239# a_3599_2340# 8.35e-19
C1520 a_7362_3239# a_7049_2340# 3.49e-20
C1521 check[1] check[5] 0.343f
C1522 a_5897_4086# a_6305_4112# 4.37e-19
C1523 a_4593_4112# a_4794_4112# 3.34e-19
C1524 VDD a_2401_2366# 0.00631f
C1525 x5.X a_6466_4775# 0.00314f
C1526 a_1511_4112# a_1762_2340# 4.16e-20
C1527 a_5845_4801# a_7247_4775# 0.0492f
C1528 a_6466_4775# a_6292_5167# 0.205f
C1529 a_6011_4801# a_6760_4775# 0.139f
C1530 x20.Q_N a_2777_2732# 8.48e-19
C1531 a_4155_4086# x77.Y 0.00176f
C1532 check[0] a_4074_4775# 5.86e-19
C1533 a_7763_2366# a_7561_2366# 3.67e-19
C1534 a_6780_2366# a_7185_2366# 2.46e-21
C1535 a_8288_2340# a_8383_2340# 0.0968f
C1536 a_9152_4775# a_10795_4801# 8.44e-20
C1537 a_9639_4775# a_10629_4801# 0.00116f
C1538 a_11543_3213# a_10982_3239# 3.79e-20
C1539 a_10628_3239# a_11493_3521# 0.00276f
C1540 a_12030_3213# a_11856_3239# 0.197f
C1541 a_11075_3605# a_11159_3605# 0.00972f
C1542 check[1] a_8402_3239# 0.0363f
C1543 VDD a_6780_2732# 0.00371f
C1544 x5.X a_8939_4086# 0.00115f
C1545 a_4019_4112# a_3912_2366# 8.38e-21
C1546 x7.X a_4453_2340# 0.181f
C1547 x27.D a_4681_4801# 2.31e-21
C1548 VDD a_9322_3521# 0.0163f
C1549 a_4658_4086# a_4970_3239# 5.48e-21
C1550 x5.X x75.Q 0.0011f
C1551 x42.Q_N a_10794_3239# 9.16e-19
C1552 eob a_2883_5674# 6.72e-19
C1553 x42.Q_N a_9872_3521# 2.75e-19
C1554 x30.Q_N a_9237_2340# 8.11e-21
C1555 a_12030_3213# a_11629_2340# 8.72e-19
C1556 a_11856_3239# a_11628_2640# 1.11e-20
C1557 a_11543_3213# a_11833_2340# 0.00144f
C1558 x66.Q_N D[2] 2.25e-19
C1559 VDD a_7264_4394# 0.00984f
C1560 x4.X a_10681_4086# 0.0036f
C1561 x4.X a_4590_2732# 9.81e-19
C1562 a_8939_4086# a_9237_4386# 0.137f
C1563 a_8697_4112# a_9238_4086# 0.125f
C1564 a_6985_4112# x42.Q_N 1.96e-20
C1565 x5.X a_3807_4801# 5.48e-19
C1566 x7.X a_7763_2366# 0.155f
C1567 x5.A a_897_4112# 5.71e-20
C1568 x4.X a_7158_3605# 4.4e-19
C1569 x4.X a_9370_4801# 5.55e-19
C1570 x7.X a_10794_3239# 0.148f
C1571 x42.Q_N a_9577_2366# 5.33e-22
C1572 x5.X a_10983_4801# 0.00551f
C1573 check[3] a_12048_4394# 5.14e-21
C1574 a_2061_2340# a_3599_2340# 0.00116f
C1575 a_6010_3239# a_6291_3605# 0.155f
C1576 a_5844_3239# a_6759_3213# 0.126f
C1577 a_9152_4775# a_9465_4801# 0.124f
C1578 D[3] a_11969_2366# 7.69e-20
C1579 a_8684_5167# a_8591_4801# 0.0367f
C1580 a_8858_4775# a_8768_5167# 6.69e-20
C1581 a_8403_4801# a_7363_4801# 4.14e-20
C1582 a_2060_2640# a_3912_2366# 1.9e-19
C1583 a_2265_2340# a_2401_2366# 0.07f
C1584 check[0] a_6759_3213# 1.67e-20
C1585 a_11628_2640# a_11629_2340# 0.781f
C1586 a_11330_2340# a_11833_2340# 0.00187f
C1587 a_11088_2366# a_12101_2550# 0.0633f
C1588 a_10775_2340# x63.Q_N 0.124f
C1589 x77.Y a_4925_2550# 0.00196f
C1590 a_4213_3239# a_4585_3239# 3.34e-19
C1591 VDD a_1822_4801# 0.00544f
C1592 a_929_3238# a_1112_2340# 0.00185f
C1593 a_4658_4086# a_4680_3239# 4.33e-20
C1594 a_4926_4296# a_4854_3213# 3.74e-20
C1595 check[5] a_6410_2366# 1.31e-19
C1596 a_3912_2366# a_5371_2366# 9.06e-21
C1597 x54.Q_N a_4112_2648# 2.02e-20
C1598 a_4657_2340# a_4590_2732# 9.46e-19
C1599 a_4452_2640# a_4871_2648# 2.46e-19
C1600 a_6010_3239# a_6304_2366# 5.94e-19
C1601 a_2853_5648# a_3600_4086# 2.47e-19
C1602 a_6465_3213# a_5991_2340# 2.5e-19
C1603 check[0] a_6546_2340# 0.00104f
C1604 x20.Q_N a_4389_4478# 3.31e-21
C1605 check[2] a_9377_4112# 6.45e-20
C1606 a_4368_4775# a_4318_5083# 1.21e-20
C1607 a_3619_4801# a_4214_4801# 0.00118f
C1608 VDD a_621_4112# 0.256f
C1609 a_3807_4801# a_3984_5167# 8.94e-19
C1610 x4.X a_4538_3521# 0.00211f
C1611 check[5] a_7764_4112# 0.00263f
C1612 check[2] x33.Q_N 0.0366f
C1613 a_12102_4296# x39.Q_N 0.00244f
C1614 x5.X a_9323_5083# 5.14e-19
C1615 check[6] a_4925_2550# 9.23e-19
C1616 a_7073_4801# a_7363_4801# 0.0282f
C1617 a_7247_4775# a_7182_4801# 4.2e-20
C1618 a_5896_2340# a_6845_2340# 1.03e-19
C1619 check[1] x45.Q_N 0.00102f
C1620 a_3618_3239# a_5844_3239# 4e-20
C1621 a_3452_3239# a_6010_3239# 2.9e-21
C1622 a_8590_3239# a_8767_3605# 8.94e-19
C1623 a_8402_3239# a_8997_3239# 0.00118f
C1624 a_9151_3213# a_9101_3521# 1.21e-20
C1625 x33.Q_N a_10628_3239# 8.92e-20
C1626 a_1061_4801# a_1511_4112# 0.00351f
C1627 a_10983_4801# a_11160_5167# 8.94e-19
C1628 a_11544_4775# a_11494_5083# 1.21e-20
C1629 a_10795_4801# a_11390_4801# 0.00118f
C1630 x33.Q_N a_9369_3239# 4.04e-19
C1631 a_1062_5674# sel_bit[1] 0.0392f
C1632 a_4453_4386# a_6305_4112# 8.96e-20
C1633 a_4658_4086# a_4794_4112# 0.07f
C1634 a_4454_4086# a_5992_4086# 2.98e-19
C1635 VDD a_2777_2732# 0.00561f
C1636 x42.Q_N a_7562_4112# 2.85e-21
C1637 VDD a_5844_3239# 0.791f
C1638 VDD check[0] 0.685f
C1639 a_9238_4086# a_9375_4478# 0.00907f
C1640 VDD a_8684_5167# 0.317f
C1641 check[6] a_5845_4801# 0.416f
C1642 x5.X D[1] 0.00133f
C1643 a_5562_4801# a_6011_4801# 4.06e-19
C1644 a_8289_4086# a_8236_3239# 5.06e-19
C1645 a_10776_4086# a_10680_2340# 2.97e-20
C1646 a_10681_4086# a_10775_2340# 1.57e-20
C1647 x42.Q_N a_7246_3213# 3.76e-21
C1648 x20.Q_N a_1520_2366# 0.0983f
C1649 a_6844_2640# a_7561_2366# 0.00105f
C1650 a_8237_4801# check[4] 8.28e-20
C1651 a_8403_4801# a_10346_4801# 9.65e-21
C1652 D[1] a_11856_3239# 3.54e-20
C1653 x33.Q_N a_9376_2366# 0.00473f
C1654 eob a_2289_4801# 0.0076f
C1655 x4.X a_6845_4386# 0.048f
C1656 check[3] a_12147_4801# 2.59e-19
C1657 a_7050_4086# x45.Q_N 0.00116f
C1658 VDD a_4592_2366# 0.00111f
C1659 x7.X a_7246_3213# 0.00381f
C1660 a_3600_4086# a_3599_2340# 5.27e-19
C1661 a_9238_4086# a_10345_3239# 4.72e-19
C1662 a_7073_4801# a_6606_4801# 0.00316f
C1663 a_10629_4801# a_10776_4086# 0.00159f
C1664 a_6466_4775# x30.Q_N 1.17e-19
C1665 a_5562_4801# a_5561_3239# 9.85e-20
C1666 a_6760_4775# a_6978_4801# 3.73e-19
C1667 check[2] check[1] 2.29f
C1668 check[0] a_5089_5083# 4.43e-19
C1669 D[1] a_11629_2340# 1.09e-20
C1670 a_9441_2340# a_9709_2550# 0.205f
C1671 a_9237_2340# x60.Q_N 1.07e-19
C1672 check[3] a_11088_2366# 1.09e-20
C1673 x33.Q_N a_11250_4775# 4.4e-20
C1674 a_3258_5648# a_3170_4801# 0.00133f
C1675 a_2389_5648# a_1511_4112# 0.00132f
C1676 sel_bit[1] a_3170_4801# 1.85e-19
C1677 VDD a_8896_2648# 0.00506f
C1678 check[2] a_9954_4112# 1.28e-19
C1679 VDD a_6376_5167# 0.0042f
C1680 a_5897_4086# a_5896_2340# 1.07e-20
C1681 x48.Q a_2463_4775# 9e-19
C1682 x7.X a_6844_2640# 0.108f
C1683 a_4855_4775# check[6] 0.0103f
C1684 VDD a_11493_3521# 0.00984f
C1685 x39.Q_N a_11565_4112# 0.0014f
C1686 a_11834_4086# a_11970_4112# 0.07f
C1687 x27.Q_N a_4388_2366# 9.43e-19
C1688 a_2265_2340# a_2777_2732# 6.69e-20
C1689 a_2060_2640# D[6] 0.00655f
C1690 a_2061_2340# a_2979_2366# 0.0708f
C1691 check[5] a_9639_4775# 2.58e-20
C1692 D[2] a_12547_2366# 6.35e-19
C1693 check[1] a_6781_4112# 1.37e-20
C1694 D[3] a_12101_2550# 1.91e-20
C1695 x5.X a_3258_5648# 0.00256f
C1696 a_1338_5674# a_1227_4801# 0.00258f
C1697 check[2] a_3877_5674# 8.16e-20
C1698 x77.Y a_6198_3239# 1.34e-20
C1699 x5.X sel_bit[1] 0.117f
C1700 a_12031_4775# check[3] 0.0678f
C1701 check[1] a_9376_2366# 3.33e-19
C1702 check[2] a_7050_4086# 4.4e-21
C1703 a_4926_4296# a_5170_4112# 0.00812f
C1704 x4.X a_6780_2732# 4.32e-19
C1705 x48.Q a_4453_4386# 1.14e-19
C1706 a_6466_4775# a_5992_4086# 4.54e-19
C1707 a_6011_4801# a_6305_4112# 9.06e-19
C1708 x7.X a_9953_2732# 8.29e-19
C1709 x4.X a_9322_3521# 9.99e-19
C1710 a_1415_4801# a_1592_5167# 8.94e-19
C1711 a_1976_4775# a_2375_5167# 0.00133f
C1712 x45.Q_N a_6410_2366# 4.18e-20
C1713 a_1508_5167# a_1822_4801# 0.0258f
C1714 x7.X a_4073_3213# 3.96e-19
C1715 x27.Q_N a_6199_4801# 3.25e-20
C1716 check[5] a_5991_2340# 2.6e-20
C1717 a_3599_2340# a_4453_2340# 0.0492f
C1718 a_3912_2366# a_4452_2640# 0.139f
C1719 a_8858_4775# a_9151_3213# 7.57e-21
C1720 a_8237_4801# a_9464_3239# 4.76e-21
C1721 check[1] a_4074_4775# 5.89e-20
C1722 a_8591_4801# x33.Q_N 4.33e-22
C1723 a_7072_3239# a_7158_3605# 0.00976f
C1724 a_6010_3239# x72.Q_N 5.46e-21
C1725 a_4970_3239# a_4789_3239# 4.11e-20
C1726 VDD a_4389_4478# 0.00402f
C1727 check[1] x20.Q_N 8.16e-19
C1728 x4.X a_7264_4394# 8.47e-19
C1729 VDD a_4767_5167# 0.00394f
C1730 a_3453_4801# a_3505_4086# 6.04e-19
C1731 a_6845_4386# a_7186_4112# 0.00118f
C1732 a_6846_4086# a_6985_4112# 2.56e-19
C1733 a_6547_4086# a_8384_4086# 1.86e-21
C1734 x45.Q_N a_7764_4112# 8.17e-20
C1735 x5.A a_1415_4801# 7.19e-20
C1736 VDD a_11943_5167# 0.00371f
C1737 check[6] a_7182_4801# 1.13e-20
C1738 a_5371_2366# a_5991_2340# 8.26e-21
C1739 a_4452_2640# a_6410_2366# 2.44e-20
C1740 D[0] a_7181_3239# 9.28e-21
C1741 a_1227_4801# a_3453_4801# 5.24e-20
C1742 x77.Y a_4367_3213# 0.106f
C1743 a_1061_4801# a_3619_4801# 2.9e-21
C1744 a_5372_4112# x7.X 4.39e-20
C1745 a_1338_5674# check[2] 2.03e-19
C1746 a_1227_4801# a_2194_4801# 0.00126f
C1747 a_1061_4801# a_2697_5083# 1.25e-19
C1748 x4.X a_1822_4801# 0.0326f
C1749 a_1062_5674# x5.A 0.129f
C1750 clk_sar a_1338_5674# 0.00117f
C1751 eob reset 3.99e-19
C1752 a_4454_4086# x48.Q_N 1.07e-19
C1753 a_4658_4086# a_4926_4296# 0.205f
C1754 x27.Q_N x7.X 0.272f
C1755 VDD a_1520_2366# 0.402f
C1756 x5.X x39.Q_N 0.00647f
C1757 a_4214_4801# a_4586_4801# 3.34e-19
C1758 x36.Q_N x7.X 0.267f
C1759 reset x4.A 0.00101f
C1760 x39.Q_N a_11856_3239# 0.162f
C1761 a_4073_3213# a_4018_2366# 5.71e-21
C1762 a_6844_2640# a_8288_2340# 6.58e-19
C1763 a_6546_2340# a_6780_2366# 0.00707f
C1764 a_6304_2366# a_6984_2366# 3.73e-19
C1765 a_9638_3213# a_9754_3239# 0.0397f
C1766 a_9151_3213# a_9573_3239# 2.87e-21
C1767 a_4680_3239# a_4789_3239# 0.00707f
C1768 x75.Q_N a_5844_3239# 2.94e-19
C1769 check[0] x75.Q_N 4.68e-20
C1770 a_8997_3239# a_9369_3239# 3.34e-19
C1771 a_11390_4801# a_11762_4801# 3.34e-19
C1772 check[1] a_6759_3213# 2.39e-20
C1773 x5.X a_6505_4394# 5.63e-19
C1774 VDD a_9377_4112# 0.00445f
C1775 VDD a_4871_2648# 0.0102f
C1776 sel_bit[0] a_2883_5674# 0.0666f
C1777 x4.X a_621_4112# 9.87e-20
C1778 VDD x33.Q_N 0.446f
C1779 check[2] a_10680_2340# 0.027f
C1780 x7.X a_2533_2550# 0.00698f
C1781 a_9237_4386# x39.Q_N 2.03e-19
C1782 check[0] a_3913_4112# 0.00318f
C1783 x5.X a_12737_3239# 0.00125f
C1784 check[4] a_10156_4112# 0.00259f
C1785 x42.Q_N a_9151_3213# 0.0983f
C1786 check[6] a_6400_4801# 1.18e-19
C1787 a_9710_4296# a_9638_3213# 3.74e-20
C1788 a_9442_4086# a_9464_3239# 4.33e-20
C1789 x20.Q_N a_3912_2366# 1.17e-19
C1790 a_5562_4801# a_4854_3213# 3.19e-20
C1791 a_8696_2366# a_8896_2648# 0.00185f
C1792 a_8383_2340# a_9172_2732# 7.71e-20
C1793 check[6] a_4367_3213# 1.13e-19
C1794 x39.Q_N a_11629_2340# 3.65e-20
C1795 a_11834_4086# a_12101_2550# 2.22e-22
C1796 a_10628_3239# a_10680_2340# 4.5e-19
C1797 x30.Q_N x57.Q_N 4.08e-19
C1798 a_12030_3213# D[2] 0.00376f
C1799 a_9754_3239# a_9236_2640# 5.05e-21
C1800 check[3] x66.Q_N 0.00297f
C1801 check[2] a_3453_4801# 9.66e-20
C1802 x4.X a_8684_5167# 0.00132f
C1803 x4.X a_5844_3239# 0.0457f
C1804 x5.X a_1592_5167# 4.22e-19
C1805 check[0] x4.X 0.245f
C1806 a_11629_4386# x7.X 2.51e-20
C1807 check[2] a_10629_4801# 0.00307f
C1808 x7.X a_9151_3213# 7.47e-19
C1809 a_6846_4086# a_7246_3213# 7.94e-19
C1810 a_7363_4801# a_6845_4386# 8.84e-21
C1811 a_7050_4086# a_6759_3213# 0.0014f
C1812 x45.Q_N a_6465_3213# 0.194f
C1813 x27.Q_N a_4018_2366# 0.0102f
C1814 a_9237_4386# a_9709_2550# 6.45e-21
C1815 a_9710_4296# a_9236_2640# 6.02e-22
C1816 x42.Q_N a_8938_2340# 0.00179f
C1817 a_7481_5083# x30.Q_N 2.02e-20
C1818 a_1207_2340# a_2533_2550# 4.7e-22
C1819 a_1762_2340# a_2061_2340# 0.0334f
C1820 a_1520_2366# a_2265_2340# 0.199f
C1821 D[2] a_11628_2640# 0.00729f
C1822 a_12030_3213# a_11969_2366# 1.2e-20
C1823 a_12737_3239# a_11629_2340# 4.83e-19
C1824 a_10629_4801# a_10628_3239# 6.9e-19
C1825 a_9236_2640# x63.Q_N 1.48e-19
C1826 check[4] check[3] 9.63e-20
C1827 a_3618_3239# a_4213_3239# 0.00118f
C1828 check[1] a_6931_5083# 4.8e-19
C1829 a_4367_3213# a_4317_3521# 1.21e-20
C1830 x5.A x5.X 0.00522f
C1831 x5.X a_4926_4296# 5.33e-19
C1832 x48.Q a_4681_4801# 0.00128f
C1833 x7.X a_8938_2340# 0.00103f
C1834 a_6846_4086# a_6844_2640# 7.02e-19
C1835 a_5992_4086# x57.Q_N 2.32e-20
C1836 VDD a_4213_3239# 0.00187f
C1837 x45.Q_N a_5991_2340# 2.01e-19
C1838 a_6845_4386# a_6845_2340# 7.25e-19
C1839 VDD check[1] 0.762f
C1840 check[5] a_8402_3239# 1.82e-19
C1841 a_2979_2366# a_4453_2340# 3.65e-21
C1842 x3.A a_653_3238# 1.87e-19
C1843 D[6] a_4452_2640# 1.85e-19
C1844 a_11970_4112# a_12030_3213# 4.45e-20
C1845 a_11629_2340# a_11768_2366# 2.56e-19
C1846 a_11628_2640# a_11969_2366# 0.00118f
C1847 a_12101_2550# a_12547_2366# 0.0367f
C1848 x4.X a_8896_2648# 0.00102f
C1849 a_3453_4801# a_4074_4775# 0.117f
C1850 a_3170_4801# x27.D 0.0749f
C1851 x7.X a_12047_2648# 6.95e-19
C1852 a_2289_4801# a_2398_4801# 0.00707f
C1853 check[2] a_9639_4775# 0.0119f
C1854 x20.Q_N a_3453_4801# 0.00252f
C1855 x4.X a_11493_3521# 2.91e-19
C1856 a_10681_4086# a_11630_4086# 7e-20
C1857 a_2194_4801# x20.Q_N 1.61e-19
C1858 check[5] a_7185_2366# 4.92e-19
C1859 VDD a_3877_5674# 3.02e-19
C1860 a_4452_2640# a_5991_2340# 3.67e-19
C1861 a_4657_2340# a_4592_2366# 9.75e-19
C1862 a_4453_2340# a_4793_2366# 6.04e-20
C1863 a_8236_3239# a_8857_3213# 0.117f
C1864 x72.Q_N a_8236_3239# 2.94e-19
C1865 a_10629_4801# a_11250_4775# 0.117f
C1866 x33.Q_N a_8683_3605# 0.00192f
C1867 VDD a_7050_4086# 0.487f
C1868 a_3913_4112# a_4389_4478# 0.00133f
C1869 x5.X x27.D 0.151f
C1870 a_4214_4801# a_3600_4086# 1.08e-19
C1871 a_8858_4775# a_8384_4086# 4.54e-19
C1872 a_8403_4801# a_8697_4112# 9.06e-19
C1873 check[0] a_7186_4112# 3.6e-20
C1874 a_3258_5648# a_3373_5674# 0.18f
C1875 a_6844_2640# a_6982_2732# 1.09e-19
C1876 a_2883_5674# a_2788_5674# 0.00133f
C1877 a_6304_2366# a_7263_2648# 1.21e-20
C1878 D[5] a_6984_2366# 8.02e-20
C1879 a_6546_2340# a_6410_2366# 0.0282f
C1880 sel_bit[1] a_3373_5674# 0.0439f
C1881 D[7] a_1996_2366# 1.53e-19
C1882 a_8236_3239# a_8383_2340# 8.35e-19
C1883 check[3] a_11834_4086# 8.07e-19
C1884 x4.X a_4389_4478# 2.12e-19
C1885 a_3618_3239# a_3912_2366# 5.94e-19
C1886 a_4073_3213# a_3599_2340# 2.5e-19
C1887 D[0] a_9754_3239# 1.61e-20
C1888 x33.Q_N a_8696_2366# 0.0928f
C1889 a_5372_4112# a_6846_4086# 3.65e-21
C1890 a_5897_4086# a_6845_4386# 9.02e-21
C1891 x5.X a_6760_4775# 0.00141f
C1892 VDD a_3912_2366# 0.359f
C1893 x27.Q_N a_6846_4086# 1.92e-21
C1894 a_1511_4112# a_2061_2340# 0.00155f
C1895 a_6011_4801# a_7073_4801# 0.137f
C1896 a_5845_4801# a_6199_4801# 0.0663f
C1897 a_6292_5167# a_6760_4775# 0.0633f
C1898 check[0] a_4368_4775# 0.00265f
C1899 x20.Q_N D[6] 0.00261f
C1900 a_4454_4086# x77.Y 2.63e-20
C1901 a_8237_4801# a_10983_4801# 3.65e-21
C1902 a_9465_4801# a_10795_4801# 2.57e-20
C1903 x33.Q_N a_11194_2366# 8.7e-20
C1904 a_10794_3239# a_11714_3521# 1.09e-19
C1905 a_11249_3213# a_11493_3521# 0.0104f
C1906 VDD a_1338_5674# 0.386f
C1907 check[1] a_8683_3605# 8.21e-20
C1908 x5.X a_9238_4086# 0.261f
C1909 x4.X a_1520_2366# 0.112f
C1910 VDD a_6410_2366# 4.84e-19
C1911 x7.X a_7953_3239# 0.00109f
C1912 check[5] x45.Q_N 5.14e-20
C1913 x7.X a_4925_2550# 0.0087f
C1914 a_10776_4086# a_11565_4478# 7.71e-20
C1915 a_11089_4112# a_11289_4394# 0.00185f
C1916 VDD a_8997_3239# 5.47e-21
C1917 eob a_3258_5648# 3.1e-19
C1918 eob sel_bit[1] 0.317f
C1919 x27.Q_N a_3599_2340# 0.142f
C1920 a_8802_2366# a_9172_2366# 4.11e-20
C1921 a_12030_3213# a_12101_2550# 1.66e-21
C1922 a_11856_3239# a_11833_2340# 1.03e-19
C1923 check[3] a_12547_2366# 0.00323f
C1924 VDD a_7764_4112# 0.109f
C1925 sel_bit[1] x4.A 8.64e-21
C1926 x4.X a_9377_4112# 6.75e-19
C1927 check[1] a_8696_2366# 0.0033f
C1928 x4.X a_4871_2648# 2.86e-19
C1929 check[6] a_4454_4086# 0.0339f
C1930 x4.X x33.Q_N 0.421f
C1931 a_8384_4086# x42.Q_N 0.154f
C1932 a_8697_4112# a_9710_4296# 0.0633f
C1933 a_8939_4086# a_9442_4086# 0.00187f
C1934 VDD a_10680_2340# 0.189f
C1935 a_9237_4386# a_9238_4086# 0.75f
C1936 x4.X a_6399_3239# 6.32e-19
C1937 a_4855_4775# a_6199_4801# 8.26e-21
C1938 clk_sar x3.A 1.29e-20
C1939 x7.X a_11075_3605# 0.0011f
C1940 x45.Q_N a_8402_3239# 9.58e-19
C1941 x5.X a_9755_4801# 2.07e-19
C1942 a_3453_4801# a_3618_3239# 8.16e-19
C1943 a_3619_4801# a_3452_3239# 9.04e-19
C1944 x45.Q_N a_7480_3521# 2.75e-19
C1945 a_8403_4801# a_9102_5083# 2.46e-19
C1946 a_8237_4801# a_9323_5083# 0.00907f
C1947 a_5844_3239# a_7072_3239# 0.0334f
C1948 a_6465_3213# a_6759_3213# 0.199f
C1949 a_2061_2340# a_4154_2340# 6.38e-20
C1950 a_2533_2550# a_3599_2340# 7.98e-21
C1951 check[3] a_12548_4112# 0.159f
C1952 a_6010_3239# a_7246_3213# 0.0264f
C1953 a_2265_2340# a_3912_2366# 9.6e-21
C1954 a_2853_5648# a_1976_4775# 1.02e-19
C1955 a_11629_2340# a_11833_2340# 0.117f
C1956 a_11628_2640# a_12101_2550# 0.145f
C1957 a_11330_2340# x63.Q_N 9.58e-21
C1958 x48.Q a_3648_5972# 0.00114f
C1959 VDD a_3453_4801# 0.841f
C1960 a_5992_4086# a_6505_4394# 0.00945f
C1961 a_8384_4086# x7.X 0.00194f
C1962 VDD a_2194_4801# 0.00214f
C1963 check[2] check[5] 7.25e-20
C1964 VDD a_10629_4801# 0.81f
C1965 x7.X a_11088_2366# 0.00716f
C1966 x45.Q_N a_7185_2366# 5.33e-22
C1967 a_9755_4801# a_9237_4386# 8.84e-21
C1968 a_4657_2340# a_4871_2648# 0.0104f
C1969 a_4452_2640# a_5371_2366# 0.159f
C1970 a_4453_2340# a_5169_2732# 0.0018f
C1971 check[1] a_3913_4112# 9.87e-21
C1972 a_6291_3605# a_6304_2366# 1.71e-19
C1973 a_5844_3239# a_6845_2340# 6.52e-20
C1974 a_6465_3213# a_6546_2340# 4.18e-20
C1975 a_6759_3213# a_5991_2340# 9.06e-19
C1976 a_6010_3239# a_6844_2640# 4.04e-20
C1977 check[0] a_6845_2340# 1.9e-19
C1978 sel_bit[0] reset 8.49e-21
C1979 a_4074_4775# a_4019_4112# 8.14e-21
C1980 check[2] a_10776_4086# 0.0128f
C1981 x5.X a_9954_4478# 1.64e-19
C1982 a_4368_4775# a_4767_5167# 0.00133f
C1983 x4.X a_4213_3239# 0.00268f
C1984 a_3453_4801# a_5089_5083# 1.25e-19
C1985 a_3619_4801# a_4586_4801# 0.00126f
C1986 a_3900_5167# a_4214_4801# 0.0258f
C1987 x5.X a_8998_4801# 9.4e-19
C1988 x20.Q_N a_4008_4801# 9.98e-20
C1989 check[1] x4.X 0.262f
C1990 a_10776_4086# a_10628_3239# 8.29e-19
C1991 a_7481_5083# a_8237_4801# 4.06e-20
C1992 D[7] a_1626_2366# 0.00202f
C1993 a_8402_3239# a_10628_3239# 4e-20
C1994 a_5991_2340# a_6546_2340# 0.197f
C1995 a_8236_3239# a_10794_3239# 2.9e-21
C1996 x33.Q_N D[4] 0.00278f
C1997 a_8236_3239# a_9872_3521# 1.25e-19
C1998 a_8683_3605# a_8997_3239# 0.0258f
C1999 a_8402_3239# a_9369_3239# 0.00126f
C2000 a_9151_3213# a_9550_3605# 0.00133f
C2001 a_1682_4775# a_1511_4112# 0.00416f
C2002 a_10629_4801# a_12265_5083# 1.25e-19
C2003 a_10795_4801# a_11762_4801# 0.00126f
C2004 x77.Y x75.Q 3.59e-19
C2005 a_11076_5167# a_11390_4801# 0.0258f
C2006 a_11544_4775# a_11943_5167# 0.00133f
C2007 x33.Q_N x69.Q_N 0.02f
C2008 x4.X a_9954_4112# 6.39e-19
C2009 a_4454_4086# a_6547_4086# 1.67e-21
C2010 a_4926_4296# a_5992_4086# 7.98e-21
C2011 VDD D[6] 0.28f
C2012 VDD a_6465_3213# 0.308f
C2013 VDD a_9639_4775# 0.72f
C2014 x5.X a_5562_4801# 0.0294f
C2015 a_8384_4086# a_9173_4112# 4.2e-20
C2016 a_9237_4386# a_9954_4478# 4.45e-20
C2017 a_9238_4086# a_9656_4394# 0.00276f
C2018 check[6] a_6466_4775# 6.88e-19
C2019 x5.X a_12738_4801# 0.0161f
C2020 sel_bit[0] a_3807_4801# 7.41e-20
C2021 x20.Q_N a_2060_2640# 0.351f
C2022 x39.Q_N D[2] 0.00168f
C2023 a_8858_4775# check[4] 9.03e-21
C2024 a_3877_5674# x4.X 4.83e-20
C2025 a_6845_2340# a_8896_2648# 4.06e-20
C2026 a_1061_4801# a_1682_4775# 0.113f
C2027 eob a_1592_5167# 5.68e-19
C2028 x33.Q_N a_10775_2340# 1.5e-19
C2029 x4.X a_7050_4086# 0.00987f
C2030 check[3] a_12030_3213# 0.00748f
C2031 a_1338_5674# a_1508_5167# 3.38e-19
C2032 VDD a_5991_2340# 0.561f
C2033 a_5897_4086# a_5844_3239# 5.06e-19
C2034 check[0] a_5897_4086# 0.116f
C2035 a_4155_4086# a_3599_2340# 1.3e-22
C2036 a_3913_4112# a_3912_2366# 1.8e-19
C2037 x7.X a_6198_3239# 0.158f
C2038 a_8289_4086# a_8383_2340# 1.57e-20
C2039 a_8384_4086# a_8288_2340# 2.97e-20
C2040 a_6760_4775# x30.Q_N 0.00766f
C2041 a_6199_4801# a_6400_4801# 3.67e-19
C2042 x27.Q_N a_6010_3239# 7.07e-20
C2043 x27.Q_N a_2979_2366# 1.34e-20
C2044 a_7247_4775# a_7481_5083# 0.00945f
C2045 check[6] x75.Q 0.0149f
C2046 a_7073_4801# a_6978_4801# 0.00276f
C2047 a_11250_4775# a_10776_4086# 4.54e-19
C2048 a_10795_4801# a_11089_4112# 9.06e-19
C2049 x39.Q_N a_11969_2366# 5.33e-22
C2050 x5.A eob 0.00158f
C2051 a_8383_2340# a_9172_2366# 4.2e-20
C2052 a_8696_2366# a_10680_2340# 7.33e-21
C2053 a_12737_3239# D[2] 0.0747f
C2054 x33.Q_N a_11544_4775# 1.35e-20
C2055 check[3] a_11628_2640# 0.0274f
C2056 a_3373_5674# x27.D 5.58e-20
C2057 check[1] D[4] 0.194f
C2058 x5.A x4.A 5.06e-21
C2059 VDD a_4790_4801# 9.01e-19
C2060 x4.X a_3912_2366# 0.105f
C2061 VDD a_9374_2732# 0.0163f
C2062 VDD a_11942_3605# 0.00371f
C2063 a_6846_4086# a_7953_3239# 4.72e-19
C2064 x7.X a_7049_2340# 0.00589f
C2065 x30.Q_N a_9238_4086# 1.91e-21
C2066 x39.Q_N a_11970_4112# 0.00173f
C2067 a_12102_4296# a_12346_4112# 0.00812f
C2068 x27.Q_N a_4793_2366# 0.0404f
C2069 check[5] a_8591_4801# 0.165f
C2070 a_2265_2340# D[6] 1.59e-19
C2071 a_7954_4801# a_7246_3213# 3.19e-20
C2072 a_2533_2550# a_2979_2366# 0.0367f
C2073 check[5] a_6759_3213# 1.11e-19
C2074 check[1] a_7186_4112# 2.11e-19
C2075 eob a_1996_2732# 4.16e-20
C2076 a_1338_5674# x4.X 4.31e-21
C2077 x77.Y a_4970_3239# 0.00967f
C2078 a_10983_4801# check[3] 1.14e-19
C2079 check[2] x45.Q_N 2.88e-21
C2080 x5.X a_6305_4112# 0.00598f
C2081 x4.X a_6410_2366# 3.78e-20
C2082 x48.Q a_4658_4086# 3.93e-19
C2083 a_6466_4775# a_6547_4086# 8.83e-20
C2084 a_5845_4801# a_6846_4086# 1.15e-19
C2085 a_6011_4801# a_6845_4386# 7.24e-20
C2086 a_6760_4775# a_5992_4086# 0.0018f
C2087 a_6292_5167# a_6305_4112# 2.81e-19
C2088 x4.X a_8997_3239# 0.00265f
C2089 a_2289_4801# a_2375_5167# 0.00976f
C2090 x7.X D[3] 0.00125f
C2091 x7.X a_1112_2340# 6.44e-19
C2092 a_4019_4112# a_3618_3239# 4.04e-21
C2093 x7.X a_4367_3213# 5.5e-19
C2094 x7.X x66.Q_N 2.08e-20
C2095 check[4] x42.Q_N 6.27e-20
C2096 x27.Q_N a_4971_4801# 0.00139f
C2097 check[5] a_6546_2340# 1.34e-19
C2098 a_4154_2340# a_4453_2340# 0.0334f
C2099 a_7246_3213# a_8236_3239# 0.00116f
C2100 a_9152_4775# a_9151_3213# 0.00121f
C2101 a_3599_2340# a_4925_2550# 4.7e-22
C2102 a_6759_3213# a_8402_3239# 1.98e-19
C2103 a_11768_2366# a_11969_2366# 3.34e-19
C2104 a_3912_2366# a_4657_2340# 0.199f
C2105 check[1] a_4368_4775# 1.09e-19
C2106 eob x27.D 4.69e-19
C2107 a_6759_3213# a_7480_3521# 0.00185f
C2108 VDD a_4019_4112# 0.0124f
C2109 x4.X a_7764_4112# 0.00621f
C2110 a_6845_4386# a_8697_4112# 1.34e-19
C2111 a_3619_4801# a_3600_4086# 6.63e-19
C2112 a_7050_4086# a_7186_4112# 0.07f
C2113 x45.Q_N a_6781_4112# 0.00138f
C2114 a_6846_4086# a_8384_4086# 2.98e-19
C2115 a_3453_4801# a_3913_4112# 3.05e-19
C2116 VDD a_4008_4801# 2.82e-19
C2117 VDD x3.A 0.204f
C2118 x4.X a_10680_2340# 0.00342f
C2119 x20.Q_N a_3505_4086# 0.00428f
C2120 check[4] x7.X 0.0222f
C2121 D[5] a_6304_2366# 8.64e-19
C2122 a_1112_2340# a_1207_2340# 0.0968f
C2123 x33.Q_N a_6845_2340# 1.52e-19
C2124 x77.Y a_4680_3239# 0.16f
C2125 x4.X a_3453_4801# 0.00472f
C2126 a_1227_4801# x20.Q_N 1.52e-19
C2127 x4.X a_2194_4801# 0.00509f
C2128 VDD check[5] 0.493f
C2129 VDD a_2060_2640# 0.329f
C2130 x4.X a_10629_4801# 0.00428f
C2131 x48.Q a_3170_4801# 0.00244f
C2132 check[2] a_10628_3239# 0.0451f
C2133 a_4214_4801# x27.Q_N 1.45e-19
C2134 a_11769_4112# a_11970_4112# 3.34e-19
C2135 a_8857_3213# a_8802_2366# 5.71e-21
C2136 x39.Q_N a_11159_3605# 8.48e-19
C2137 check[1] a_8897_4394# 9.73e-20
C2138 a_6546_2340# a_7185_2366# 0.00316f
C2139 a_6304_2366# a_8383_2340# 7.3e-21
C2140 a_6844_2640# a_6984_2366# 0.00126f
C2141 x33.Q_N a_10155_2366# 0.032f
C2142 a_9464_3239# a_9573_3239# 0.00707f
C2143 a_11390_4801# x36.Q_N 4.02e-20
C2144 VDD a_10776_4086# 0.716f
C2145 x5.X a_6983_4478# 7.44e-19
C2146 x5.X x48.Q 0.203f
C2147 sel_bit[0] a_3258_5648# 0.0205f
C2148 VDD a_5371_2366# 0.109f
C2149 VDD a_8402_3239# 0.275f
C2150 a_6466_4775# a_6411_4112# 8.14e-21
C2151 sel_bit[0] sel_bit[1] 0.428f
C2152 VDD a_7480_3521# 0.00506f
C2153 a_1926_5083# x27.D 3.95e-22
C2154 a_9442_4086# x39.Q_N 3.43e-20
C2155 check[0] a_4453_4386# 0.164f
C2156 a_4794_4112# x77.Y 7.13e-20
C2157 x42.Q_N a_9464_3239# 0.162f
C2158 a_8383_2340# a_8802_2366# 0.0397f
C2159 x39.Q_N a_12101_2550# 0.00196f
C2160 a_8938_2340# a_9172_2732# 0.00976f
C2161 a_8696_2366# a_9374_2732# 0.00652f
C2162 x33.Q_N a_10346_4801# 0.184f
C2163 a_9754_3239# a_9441_2340# 3.49e-20
C2164 check[1] a_6845_2340# 6.25e-19
C2165 check[2] a_4074_4775# 1.07e-19
C2166 x4.X D[6] 0.00589f
C2167 a_7318_4296# a_7562_4112# 0.00812f
C2168 x4.X a_6465_3213# 0.00499f
C2169 x4.X a_9639_4775# 0.103f
C2170 VDD a_653_3238# 0.268f
C2171 x5.X a_2147_5083# 4.05e-19
C2172 check[2] x20.Q_N 4.28e-20
C2173 a_11834_4086# x7.X 4.39e-21
C2174 x27.D x48.Q_N 8.11e-20
C2175 a_7050_4086# a_7072_3239# 4.33e-20
C2176 a_7363_4801# a_7050_4086# 7.76e-20
C2177 a_7318_4296# a_7246_3213# 3.74e-20
C2178 x7.X a_9464_3239# 1.93e-19
C2179 x45.Q_N a_6759_3213# 0.0983f
C2180 x42.Q_N a_9237_2340# 3.65e-20
C2181 a_9442_4086# a_9709_2550# 2.22e-22
C2182 a_10155_2366# a_9953_2366# 3.67e-19
C2183 a_10795_4801# a_10794_3239# 1.39e-19
C2184 a_10680_2340# a_10775_2340# 0.0968f
C2185 a_2060_2640# a_2265_2340# 0.153f
C2186 a_9172_2366# a_9577_2366# 2.46e-21
C2187 a_1520_2366# x51.Q_N 0.00553f
C2188 D[2] a_11833_2340# 4.68e-20
C2189 a_3899_3605# a_4213_3239# 0.0258f
C2190 a_3806_3239# a_3983_3605# 8.94e-19
C2191 a_3618_3239# a_4585_3239# 0.00126f
C2192 a_4367_3213# a_4766_3605# 0.00133f
C2193 a_3452_3239# a_5088_3521# 1.25e-19
C2194 x4.X a_5991_2340# 0.111f
C2195 VDD a_11564_2732# 0.00371f
C2196 x48.Q a_3984_5167# 5.76e-19
C2197 VDD a_4585_3239# 0.00112f
C2198 a_3600_4086# a_3452_3239# 8.29e-19
C2199 x7.X a_9237_2340# 0.184f
C2200 a_6845_4386# a_7317_2550# 6.45e-21
C2201 a_7318_4296# a_6844_2640# 6.02e-22
C2202 x45.Q_N a_6546_2340# 0.0018f
C2203 x27.Q_N a_6984_2366# 2.64e-20
C2204 D[6] a_4657_2340# 2.71e-19
C2205 a_5844_3239# D[0] 7.04e-20
C2206 a_6010_3239# a_7953_3239# 1e-20
C2207 reset comparator_out 0.00121f
C2208 a_11833_2340# a_11969_2366# 0.07f
C2209 VDD a_3505_4086# 0.212f
C2210 VDD a_11565_4478# 0.00371f
C2211 x4.X a_4790_4801# 2.39e-19
C2212 x4.X a_9374_2732# 9.81e-19
C2213 a_3453_4801# a_4368_4775# 0.125f
C2214 a_3619_4801# a_3900_5167# 0.155f
C2215 x4.X a_11942_3605# 4.4e-19
C2216 x5.X a_8403_4801# 0.0201f
C2217 x7.X a_12547_2366# 0.155f
C2218 x20.Q_N a_4074_4775# 8.63e-20
C2219 a_10156_4112# x39.Q_N 8.08e-20
C2220 x30.Q_N a_6305_4112# 1.32e-21
C2221 a_10776_4086# a_11331_4086# 0.197f
C2222 a_6760_4775# a_8237_4801# 1.67e-19
C2223 a_6011_4801# a_5844_3239# 9.04e-19
C2224 a_5845_4801# a_6010_3239# 8.16e-19
C2225 a_2853_5648# a_2883_5674# 0.224f
C2226 check[0] a_6011_4801# 4.88e-19
C2227 check[1] a_5897_4086# 1.24e-21
C2228 x33.Q_N a_11630_4086# 1.91e-21
C2229 check[5] a_8696_2366# 2.42e-20
C2230 a_8402_3239# a_8683_3605# 0.155f
C2231 a_8236_3239# a_9151_3213# 0.126f
C2232 a_4925_2550# a_4793_2366# 0.0258f
C2233 a_4452_2640# a_6546_2340# 4.11e-20
C2234 a_4453_2340# a_6304_2366# 3.16e-19
C2235 VDD a_1227_4801# 0.34f
C2236 x27.Q_N a_4007_3239# 6.74e-20
C2237 a_9639_4775# x69.Q_N 4.45e-20
C2238 a_10629_4801# a_11544_4775# 0.125f
C2239 x33.Q_N a_9638_3213# 0.0126f
C2240 a_10795_4801# a_11076_5167# 0.155f
C2241 a_4155_4086# a_4591_4478# 0.00412f
C2242 a_3913_4112# a_4019_4112# 0.0552f
C2243 a_4453_4386# a_4389_4478# 2.13e-19
C2244 VDD x45.Q_N 0.458f
C2245 a_4454_4086# a_4113_4394# 1.25e-19
C2246 a_4454_4086# x7.X 3.22e-20
C2247 a_12548_4112# x7.X 4.04e-20
C2248 a_8858_4775# a_8939_4086# 8.83e-20
C2249 a_8684_5167# a_8697_4112# 2.81e-19
C2250 a_9152_4775# a_8384_4086# 0.0018f
C2251 a_8403_4801# a_9237_4386# 7.24e-20
C2252 a_8237_4801# a_9238_4086# 1.15e-19
C2253 a_3373_5674# a_3876_6040# 0.00336f
C2254 a_6844_2640# a_7263_2648# 2.46e-19
C2255 check[3] x39.Q_N 1.04e-19
C2256 a_7049_2340# a_6982_2732# 9.46e-19
C2257 a_6304_2366# a_7763_2366# 5.76e-21
C2258 sel_bit[1] a_2788_5674# 2.36e-19
C2259 x57.Q_N a_6504_2648# 2.02e-20
C2260 check[0] a_5561_3239# 0.0043f
C2261 a_8857_3213# a_8383_2340# 2.5e-19
C2262 D[7] a_2401_2366# 4.38e-19
C2263 a_5561_3239# a_5844_3239# 8.18e-19
C2264 a_8402_3239# a_8696_2366# 5.94e-19
C2265 x4.X a_4019_4112# 0.00642f
C2266 a_3618_3239# a_4452_2640# 4.04e-20
C2267 a_4073_3213# a_4154_2340# 4.18e-20
C2268 a_3452_3239# a_4453_2340# 6.52e-20
C2269 a_4367_3213# a_3599_2340# 9.06e-19
C2270 a_3899_3605# a_3912_2366# 1.71e-19
C2271 x33.Q_N a_9236_2640# 0.572f
C2272 a_5992_4086# a_6305_4112# 0.272f
C2273 x4.X a_4008_4801# 8.46e-20
C2274 x4.X x3.A 2.12e-20
C2275 VDD a_4452_2640# 0.273f
C2276 x5.X a_7073_4801# 0.00115f
C2277 a_1511_4112# a_2533_2550# 6.53e-19
C2278 x4.X a_11184_4801# 8.46e-20
C2279 a_6760_4775# a_7247_4775# 0.273f
C2280 a_6011_4801# a_6376_5167# 4.45e-20
C2281 x5.A sel_bit[0] 0.0387f
C2282 a_6466_4775# a_6199_4801# 6.99e-20
C2283 check[0] a_4681_4801# 0.00122f
C2284 a_4926_4296# x77.Y 0.00166f
C2285 a_8288_2340# a_9237_2340# 1.03e-19
C2286 x30.Q_N a_7181_3239# 1.68e-19
C2287 check[3] a_12737_3239# 0.0275f
C2288 a_10794_3239# a_11389_3239# 0.00118f
C2289 a_11543_3213# a_11493_3521# 1.21e-20
C2290 a_10982_3239# a_11159_3605# 8.94e-19
C2291 VDD check[2] 0.713f
C2292 VDD clk_sar 0.114f
C2293 x4.X check[5] 0.0317f
C2294 x4.X a_2060_2640# 0.00821f
C2295 x5.X a_9710_4296# 6.08e-19
C2296 VDD a_7561_2732# 0.0042f
C2297 VDD a_10628_3239# 0.791f
C2298 VDD a_9369_3239# 6.2e-19
C2299 a_11089_4112# a_11767_4478# 0.00652f
C2300 a_11331_4086# a_11565_4478# 0.00976f
C2301 a_10776_4086# a_11195_4112# 0.0397f
C2302 x27.Q_N a_4154_2340# 0.16f
C2303 a_9236_2640# a_9953_2366# 0.00105f
C2304 check[3] a_11768_2366# 9.26e-20
C2305 VDD a_6781_4112# 3.56e-19
C2306 x4.X a_10776_4086# 0.1f
C2307 check[1] a_9236_2640# 3.18e-19
C2308 x4.X a_5371_2366# 8.28e-20
C2309 x4.X a_8402_3239# 0.0429f
C2310 a_9237_4386# a_9710_4296# 0.155f
C2311 a_8939_4086# x42.Q_N 0.0287f
C2312 VDD a_9376_2366# 6.2e-19
C2313 a_9238_4086# a_9442_4086# 0.117f
C2314 x4.X a_7480_3521# 0.00103f
C2315 x7.X a_12030_3213# 0.00336f
C2316 a_4368_4775# a_4790_4801# 2.87e-21
C2317 a_4855_4775# a_4971_4801# 0.0397f
C2318 a_8858_4775# a_8803_4112# 8.14e-21
C2319 x3.A x7.A 0.00115f
C2320 a_3619_4801# a_4073_3213# 3.18e-21
C2321 a_3900_5167# a_3452_3239# 8.3e-21
C2322 x5.X a_11494_5083# 3.98e-19
C2323 sel_bit[0] x27.D 0.00108f
C2324 a_7954_4801# a_7953_3239# 9.85e-20
C2325 x20.Q_N a_3618_3239# 0.0017f
C2326 a_621_4112# a_897_4112# 0.00202f
C2327 a_8403_4801# a_9551_5167# 2.13e-19
C2328 a_8858_4775# a_9323_5083# 9.46e-19
C2329 a_8237_4801# a_8998_4801# 6.04e-20
C2330 a_6291_3605# a_7246_3213# 4.7e-22
C2331 a_6010_3239# a_6198_3239# 0.163f
C2332 a_6465_3213# a_7072_3239# 0.00187f
C2333 a_5844_3239# a_6375_3605# 0.0018f
C2334 a_1520_2366# x54.Q_N 5.89e-21
C2335 a_2061_2340# a_4453_2340# 0.00176f
C2336 check[1] a_2463_4775# 0.00193f
C2337 a_11629_2340# x63.Q_N 1.07e-19
C2338 a_11833_2340# a_12101_2550# 0.205f
C2339 eob a_1996_2366# 1.64e-21
C2340 x48.Q a_3373_5674# 0.0679f
C2341 a_6305_4112# a_6781_4478# 0.00133f
C2342 VDD a_4074_4775# 0.494f
C2343 a_1976_4775# a_1511_4112# 0.00824f
C2344 VDD x20.Q_N 1.29f
C2345 x4.X a_653_3238# 5.14e-19
C2346 VDD a_11250_4775# 0.488f
C2347 x7.X x75.Q 0.00133f
C2348 x7.X a_11628_2640# 0.108f
C2349 a_5845_4801# a_7954_4801# 1.03e-19
C2350 a_9755_4801# a_9442_4086# 7.76e-20
C2351 check[5] D[4] 0.00424f
C2352 a_7953_3239# a_8236_3239# 8.18e-19
C2353 a_4453_2340# D[5] 0.338f
C2354 check[1] a_4453_4386# 1.28e-20
C2355 a_4657_2340# a_5371_2366# 6.99e-20
C2356 a_4925_2550# a_5169_2732# 0.00972f
C2357 a_7246_3213# a_6304_2366# 8.4e-19
C2358 x33.Q_N D[0] 1.28e-20
C2359 a_6010_3239# a_7049_2340# 0.00154f
C2360 check[0] a_7317_2550# 1.78e-19
C2361 a_6759_3213# a_6546_2340# 2.17e-19
C2362 a_10346_4801# a_10629_4801# 8.18e-19
C2363 a_6465_3213# a_6845_2340# 0.00199f
C2364 a_1061_4801# a_1976_4775# 0.117f
C2365 a_1227_4801# a_1508_5167# 0.151f
C2366 a_3505_4086# a_3913_4112# 6.04e-19
C2367 x4.X a_11564_2732# 4.32e-19
C2368 x5.X a_10681_4086# 0.0752f
C2369 check[2] a_11331_4086# 3.82e-19
C2370 a_4681_4801# a_4767_5167# 0.00976f
C2371 a_2579_4801# a_2398_4801# 4.11e-20
C2372 x4.X a_4585_3239# 5e-19
C2373 a_3619_4801# x27.Q_N 1.18e-19
C2374 a_10983_4801# x7.X 1.78e-20
C2375 x5.X a_9370_4801# 2.59e-19
C2376 a_10776_4086# a_11249_3213# 2.45e-19
C2377 a_11089_4112# a_10794_3239# 4.9e-19
C2378 x45.Q_N x75.Q_N 6.77e-21
C2379 x30.Q_N a_8403_4801# 2.26e-19
C2380 a_5991_2340# a_6845_2340# 0.0492f
C2381 a_6304_2366# a_6844_2640# 0.139f
C2382 a_4367_3213# a_6010_3239# 2.89e-19
C2383 eob x48.Q 0.0102f
C2384 a_4854_3213# a_5844_3239# 0.00116f
C2385 check[0] a_4854_3213# 0.00313f
C2386 a_9464_3239# a_9550_3605# 0.00976f
C2387 x33.Q_N a_11543_3213# 8.28e-21
C2388 a_8402_3239# x69.Q_N 4.5e-21
C2389 a_7362_3239# a_7181_3239# 4.11e-20
C2390 x4.X a_3505_4086# 0.0122f
C2391 a_11857_4801# a_11943_5167# 0.00976f
C2392 a_10795_4801# x36.Q_N 2.98e-20
C2393 a_9755_4801# a_9574_4801# 4.11e-20
C2394 x4.X a_11565_4478# 2.12e-19
C2395 a_4454_4086# a_6846_4086# 1.37e-19
C2396 a_3913_4112# x45.Q_N 1.22e-20
C2397 x48.Q x4.A 1.09e-20
C2398 a_8939_4086# a_9173_4112# 0.00707f
C2399 VDD a_6759_3213# 0.353f
C2400 a_9238_4086# a_10156_4112# 0.0663f
C2401 VDD a_8591_4801# 0.109f
C2402 a_9237_4386# a_10681_4086# 3.59e-19
C2403 x42.Q_N a_8803_4112# 0.0446f
C2404 a_8697_4112# a_9377_4112# 3.73e-19
C2405 a_9442_4086# a_9954_4478# 6.69e-20
C2406 check[2] a_8696_2366# 1.08e-21
C2407 check[6] a_6760_4775# 0.00308f
C2408 a_8384_4086# a_8236_3239# 8.29e-19
C2409 x33.Q_N a_8697_4112# 7.32e-22
C2410 a_653_3238# x7.A 0.129f
C2411 x20.Q_N a_2265_2340# 0.194f
C2412 a_10776_4086# a_10775_2340# 5.27e-19
C2413 x30.Q_N a_5896_2340# 3.7e-19
C2414 a_1227_4801# x4.X 0.311f
C2415 a_7763_2366# a_8383_2340# 8.26e-21
C2416 a_9152_4775# check[4] 0.00456f
C2417 a_9639_4775# a_10346_4801# 0.0968f
C2418 a_6844_2640# a_8802_2366# 1.71e-20
C2419 D[1] a_9573_3239# 9.28e-21
C2420 eob a_2147_5083# 0.00298f
C2421 x33.Q_N a_11330_2340# 5.36e-20
C2422 x4.X x45.Q_N 0.252f
C2423 check[1] D[0] 0.169f
C2424 a_2389_5648# a_1976_4775# 1.09e-19
C2425 VDD a_6546_2340# 0.177f
C2426 check[2] a_11194_2366# 0.00242f
C2427 check[0] a_4593_4112# 5.07e-20
C2428 a_4453_4386# a_3912_2366# 1.93e-22
C2429 x42.Q_N D[1] 0.00176f
C2430 a_10795_4801# a_11629_4386# 7.24e-20
C2431 a_7073_4801# x30.Q_N 4.49e-19
C2432 a_11076_5167# a_11089_4112# 2.81e-19
C2433 a_11250_4775# a_11331_4086# 8.83e-20
C2434 a_11544_4775# a_10776_4086# 0.0018f
C2435 a_10629_4801# a_11630_4086# 1.15e-19
C2436 a_4971_4801# a_4367_3213# 1.05e-20
C2437 a_9236_2640# a_10680_2340# 6.83e-19
C2438 a_8696_2366# a_9376_2366# 3.73e-19
C2439 a_8938_2340# a_9172_2366# 0.00707f
C2440 a_3452_3239# a_4073_3213# 0.115f
C2441 x33.Q_N a_11857_4801# 1.75e-20
C2442 a_8998_4801# a_9574_4801# 2.46e-21
C2443 check[3] a_11833_2340# 6.99e-20
C2444 check[1] a_6011_4801# 4e-19
C2445 a_11389_3239# a_11761_3239# 3.34e-19
C2446 check[2] a_3913_4112# 1.35e-20
C2447 x4.X a_4452_2640# 0.00799f
C2448 VDD a_6931_5083# 0.0163f
C2449 check[2] a_11195_4112# 4.22e-19
C2450 VDD a_9655_2648# 0.00984f
C2451 a_5992_4086# a_5896_2340# 2.97e-20
C2452 a_5897_4086# a_5991_2340# 1.57e-20
C2453 x7.X D[1] 0.025f
C2454 VDD a_3618_3239# 0.291f
C2455 x7.X x57.Q_N 2.04e-19
C2456 x27.Q_N a_6304_2366# 8.23e-20
C2457 check[5] a_7363_4801# 8.69e-20
C2458 a_10775_2340# a_11564_2732# 7.71e-20
C2459 a_11088_2366# a_11288_2648# 0.00185f
C2460 check[1] a_8697_4112# 0.00119f
C2461 check[2] x4.X 0.258f
C2462 x5.X a_6845_4386# 0.0101f
C2463 x4.X a_7561_2732# 1.17e-19
C2464 x48.Q x48.Q_N 0.00314f
C2465 x4.X a_10628_3239# 0.0456f
C2466 a_6760_4775# a_6547_4086# 3.72e-19
C2467 a_7247_4775# a_6305_4112# 0.00161f
C2468 a_9954_4478# a_10156_4112# 8.94e-19
C2469 a_6011_4801# a_7050_4086# 0.00221f
C2470 a_8803_4112# a_9173_4112# 4.11e-20
C2471 a_6466_4775# a_6846_4086# 0.00336f
C2472 a_1976_4775# a_3619_4801# 2.05e-19
C2473 a_2463_4775# a_3453_4801# 0.00116f
C2474 x4.X a_9369_3239# 4.91e-19
C2475 a_1508_5167# x20.Q_N 9.58e-20
C2476 a_1976_4775# a_2697_5083# 0.00185f
C2477 a_4019_4112# a_3899_3605# 1.12e-20
C2478 x7.X a_4680_3239# 1.77e-19
C2479 check[5] a_6845_2340# 0.0379f
C2480 a_4214_4801# a_4367_3213# 1.61e-20
C2481 x27.Q_N a_3452_3239# 2.63e-19
C2482 a_7072_3239# a_8402_3239# 3.9e-20
C2483 a_9639_4775# a_9638_3213# 0.00237f
C2484 a_6759_3213# a_8683_3605# 4.38e-20
C2485 a_5844_3239# a_8590_3239# 3.65e-21
C2486 a_3912_2366# x54.Q_N 0.00553f
C2487 a_4452_2640# a_4657_2340# 0.153f
C2488 check[1] a_4681_4801# 3.58e-20
C2489 a_7246_3213# x72.Q_N 0.124f
C2490 a_2853_5648# a_3807_4801# 1.57e-19
C2491 VDD a_5170_4478# 0.00436f
C2492 x4.X a_6781_4112# 8.67e-20
C2493 x36.Q_N a_11389_3239# 6.11e-19
C2494 a_7318_4296# a_8384_4086# 7.98e-21
C2495 a_3453_4801# a_4453_4386# 9.86e-20
C2496 a_3900_5167# a_3600_4086# 4.9e-20
C2497 a_4074_4775# a_3913_4112# 0.0025f
C2498 a_6846_4086# a_8939_4086# 1.67e-21
C2499 x45.Q_N a_7186_4112# 0.00171f
C2500 VDD a_5089_5083# 0.00529f
C2501 x20.Q_N a_3913_4112# 7.65e-19
C2502 check[0] a_5170_4112# 8.39e-20
C2503 VDD a_12265_5083# 0.00506f
C2504 a_6606_4801# check[5] 1.24e-20
C2505 a_11250_4775# a_11195_4112# 8.14e-21
C2506 D[7] a_1520_2366# 0.00164f
C2507 D[5] a_6844_2640# 4.09e-20
C2508 a_5371_2366# a_6845_2340# 3.65e-21
C2509 x33.Q_N a_10345_3239# 0.0101f
C2510 D[0] a_8997_3239# 1.6e-19
C2511 check[4] a_11390_4801# 1.64e-19
C2512 x4.X a_4074_4775# 0.00101f
C2513 x4.X x20.Q_N 0.274f
C2514 x4.X a_11250_4775# 9.45e-19
C2515 VDD a_2265_2340# 0.326f
C2516 a_5562_4801# check[6] 0.133f
C2517 a_4586_4801# x27.Q_N 1.61e-19
C2518 check[2] x69.Q_N 4.68e-20
C2519 a_10628_3239# a_11249_3213# 0.117f
C2520 a_7049_2340# a_6984_2366# 9.75e-19
C2521 a_6845_2340# a_7185_2366# 6.04e-20
C2522 a_6844_2640# a_8383_2340# 3.42e-19
C2523 check[1] a_9375_4478# 6.38e-20
C2524 x69.Q_N a_10628_3239# 2.94e-19
C2525 x75.Q_N a_6759_3213# 2.97e-20
C2526 a_12738_4801# check[3] 0.175f
C2527 a_11762_4801# x36.Q_N 4.04e-20
C2528 VDD a_11331_4086# 0.34f
C2529 x5.X a_7264_4394# 3.07e-19
C2530 sel_bit[0] a_3876_6040# 0.00262f
C2531 VDD a_8683_3605# 0.176f
C2532 check[2] a_10775_2340# 0.0128f
C2533 check[0] a_4658_4086# 7.37e-19
C2534 x42.Q_N a_8767_3605# 8.48e-19
C2535 x27.Q_N a_2061_2340# 1.55e-19
C2536 a_9236_2640# a_9374_2732# 1.09e-19
C2537 a_10628_3239# a_10775_2340# 8.35e-19
C2538 check[4] a_8236_3239# 1.94e-20
C2539 a_8696_2366# a_9655_2648# 1.21e-20
C2540 a_8938_2340# a_8802_2366# 0.0282f
C2541 D[4] a_9376_2366# 7.47e-20
C2542 a_6781_4112# a_7186_4112# 2.46e-21
C2543 a_8289_4086# a_8384_4086# 0.0968f
C2544 check[2] a_4368_4775# 1.3e-19
C2545 x4.X a_8591_4801# 2.37e-19
C2546 x39.Q_N x7.X 6.03e-19
C2547 x4.X a_6759_3213# 0.111f
C2548 VDD a_8696_2366# 0.348f
C2549 a_3619_4801# a_5845_4801# 4e-20
C2550 a_3453_4801# a_6011_4801# 2.9e-21
C2551 x45.Q_N a_7072_3239# 0.162f
C2552 x27.Q_N D[5] 0.00536f
C2553 x42.Q_N a_9709_2550# 0.00196f
C2554 a_8237_4801# a_8403_4801# 0.751f
C2555 x36.Q_N a_11089_4112# 1.39e-22
C2556 a_2061_2340# a_2533_2550# 0.15f
C2557 a_2060_2640# x51.Q_N 4.18e-21
C2558 a_10795_4801# a_11075_3605# 8.52e-21
C2559 a_11250_4775# a_11249_3213# 2.59e-19
C2560 a_11544_4775# a_10628_3239# 9.66e-21
C2561 a_11076_5167# a_10794_3239# 1.65e-21
C2562 a_3618_3239# x75.Q_N 1.93e-21
C2563 a_4680_3239# a_4766_3605# 0.00976f
C2564 VDD a_1508_5167# 0.197f
C2565 VDD a_11194_2366# 4.84e-19
C2566 x4.X a_6546_2340# 0.00704f
C2567 x7.X a_12737_3239# 1.9e-19
C2568 x7.X a_9709_2550# 0.00825f
C2569 x45.Q_N a_6845_2340# 3.65e-20
C2570 a_3600_4086# a_4073_3213# 2.45e-19
C2571 a_7050_4086# a_7317_2550# 2.22e-22
C2572 VDD x75.Q_N 0.0719f
C2573 a_3913_4112# a_3618_3239# 4.9e-19
C2574 a_6465_3213# D[0] 1.23e-20
C2575 D[6] x54.Q_N 0.00317f
C2576 a_12101_2550# a_12345_2366# 0.00812f
C2577 VDD a_3913_4112# 0.46f
C2578 VDD a_11195_4112# 0.00996f
C2579 x4.X a_9655_2648# 2.86e-19
C2580 a_3453_4801# a_4681_4801# 0.0334f
C2581 a_3619_4801# a_4855_4775# 0.0265f
C2582 x4.X a_3618_3239# 0.0489f
C2583 a_4074_4775# a_4368_4775# 0.199f
C2584 x4.X a_11183_3239# 6.32e-19
C2585 a_10776_4086# a_11630_4086# 0.0492f
C2586 x30.Q_N a_6845_4386# 0.0327f
C2587 x5.X a_5844_3239# 8.91e-20
C2588 x5.X a_8684_5167# 0.00465f
C2589 a_6606_4801# x45.Q_N 2.3e-19
C2590 x20.Q_N a_4368_4775# 3e-20
C2591 a_11089_4112# a_11629_4386# 0.139f
C2592 a_2853_5648# a_3258_5648# 0.0197f
C2593 x5.X check[0] 0.789f
C2594 a_2853_5648# sel_bit[1] 0.0368f
C2595 sel_bit[0] x48.Q 0.0566f
C2596 a_7073_4801# a_8237_4801# 6.38e-20
C2597 a_6292_5167# a_5844_3239# 8.3e-21
C2598 a_6011_4801# a_6465_3213# 3.18e-21
C2599 a_7247_4775# a_8403_4801# 2.64e-19
C2600 x48.Q x77.Y 6.96e-20
C2601 a_7246_3213# a_7763_2366# 2.38e-19
C2602 a_4925_2550# a_6304_2366# 9.52e-21
C2603 a_8236_3239# a_9464_3239# 0.0334f
C2604 a_4452_2640# a_6845_2340# 2.9e-21
C2605 a_8402_3239# a_9638_3213# 0.0264f
C2606 a_4453_2340# a_6844_2640# 4e-20
C2607 a_8857_3213# a_9151_3213# 0.199f
C2608 VDD x4.X 5.73f
C2609 x72.Q_N a_9151_3213# 2.97e-20
C2610 a_10795_4801# a_12031_4775# 0.0264f
C2611 a_10629_4801# a_11857_4801# 0.0334f
C2612 a_11250_4775# a_11544_4775# 0.199f
C2613 a_2883_5674# a_1511_4112# 1.46e-20
C2614 a_4454_4086# a_4591_4478# 0.00907f
C2615 a_8858_4775# a_9238_4086# 0.00336f
C2616 check[6] a_5169_2366# 5.24e-20
C2617 a_8403_4801# a_9442_4086# 0.00221f
C2618 a_9639_4775# a_8697_4112# 0.00161f
C2619 a_9152_4775# a_8939_4086# 3.72e-19
C2620 a_3258_5648# a_3671_5674# 3.58e-19
C2621 a_6845_2340# a_7561_2732# 0.0018f
C2622 a_6844_2640# a_7763_2366# 0.159f
C2623 a_7049_2340# a_7263_2648# 0.0104f
C2624 x75.Q a_6010_3239# 0.00207f
C2625 a_8402_3239# a_9236_2640# 4.04e-20
C2626 a_9151_3213# a_8383_2340# 9.06e-19
C2627 a_8683_3605# a_8696_2366# 1.71e-19
C2628 a_8857_3213# a_8938_2340# 4.18e-20
C2629 a_8236_3239# a_9237_2340# 6.52e-20
C2630 a_3618_3239# a_4657_2340# 0.00154f
C2631 a_4854_3213# a_3912_2366# 8.4e-19
C2632 a_4367_3213# a_4154_2340# 2.17e-19
C2633 a_4073_3213# a_4453_2340# 0.00199f
C2634 x33.Q_N a_9441_2340# 0.179f
C2635 x4.X a_5170_4478# 9.15e-19
C2636 a_5897_4086# x45.Q_N 0.182f
C2637 a_5992_4086# a_6845_4386# 0.0264f
C2638 a_6305_4112# a_6547_4086# 0.124f
C2639 VDD a_4657_2340# 0.307f
C2640 x5.X a_6376_5167# 4.16e-19
C2641 a_6292_5167# a_6376_5167# 0.00972f
C2642 a_7247_4775# a_7073_4801# 0.197f
C2643 a_6760_4775# a_6199_4801# 8.23e-22
C2644 a_5845_4801# a_6710_5083# 0.00276f
C2645 a_8383_2340# a_8938_2340# 0.197f
C2646 x33.Q_N a_11564_2366# 1e-20
C2647 a_9639_4775# a_11857_4801# 1.86e-21
C2648 a_10794_3239# a_11761_3239# 0.00126f
C2649 a_11075_3605# a_11389_3239# 0.0258f
C2650 a_10628_3239# a_12264_3521# 1.25e-19
C2651 a_11543_3213# a_11942_3605# 0.00133f
C2652 check[1] a_8590_3239# 0.00666f
C2653 VDD x7.A 0.213f
C2654 VDD D[4] 0.221f
C2655 x4.X a_2265_2340# 0.00118f
C2656 VDD a_11249_3213# 0.308f
C2657 a_11089_4112# a_12048_4394# 1.21e-20
C2658 VDD x69.Q_N 0.0716f
C2659 check[2] a_10346_4801# 0.0147f
C2660 a_11629_4386# a_11767_4478# 1.09e-19
C2661 a_11331_4086# a_11195_4112# 0.0282f
C2662 x27.D a_4539_5083# 3.01e-21
C2663 eob a_2993_5674# 9.62e-20
C2664 a_1207_2340# a_1996_2732# 7.71e-20
C2665 a_1520_2366# a_1720_2648# 0.00185f
C2666 x42.Q_N a_10982_3239# 1.34e-20
C2667 a_9442_4086# a_9754_3239# 5.48e-21
C2668 x27.Q_N a_4453_2340# 0.0462f
C2669 a_9237_2340# a_11288_2648# 4.06e-20
C2670 check[3] a_12345_2366# 5.09e-20
C2671 a_2389_5648# a_2883_5674# 0.169f
C2672 check[2] a_2784_5996# 6.63e-19
C2673 VDD a_7186_4112# 0.0326f
C2674 x5.X a_4389_4478# 4.04e-20
C2675 check[2] a_5897_4086# 1.35e-21
C2676 check[1] a_9441_2340# 4.56e-19
C2677 x4.X a_11331_4086# 0.00706f
C2678 x4.X a_8683_3605# 0.0177f
C2679 a_9238_4086# x42.Q_N 0.00114f
C2680 a_9442_4086# a_9710_4296# 0.205f
C2681 VDD a_10775_2340# 0.561f
C2682 x7.X a_10982_3239# 0.157f
C2683 a_4681_4801# a_4790_4801# 0.00707f
C2684 x5.X a_11943_5167# 1.78e-19
C2685 a_3619_4801# a_4367_3213# 2.05e-21
C2686 a_4074_4775# a_3899_3605# 1.33e-23
C2687 a_3900_5167# a_4073_3213# 3.52e-21
C2688 check[5] D[0] 0.417f
C2689 x20.Q_N a_3899_3605# 2.96e-20
C2690 a_2060_2640# x54.Q_N 1.48e-19
C2691 a_6010_3239# a_4970_3239# 7.73e-20
C2692 a_6465_3213# a_6375_3605# 6.69e-20
C2693 a_8858_4775# a_8998_4801# 0.07f
C2694 a_7363_4801# a_6759_3213# 1.05e-20
C2695 a_6759_3213# a_7072_3239# 0.124f
C2696 a_6291_3605# a_6198_3239# 0.0367f
C2697 check[4] a_9172_2366# 2.2e-20
C2698 a_8403_4801# a_8792_4801# 0.0019f
C2699 a_8237_4801# a_9370_4801# 2.56e-19
C2700 a_9152_4775# a_9323_5083# 0.00652f
C2701 x36.Q_N a_10794_3239# 3.85e-19
C2702 x48.Q a_2788_5674# 1.65e-19
C2703 a_6305_4112# a_6411_4112# 0.051f
C2704 a_6845_4386# a_6781_4478# 2.13e-19
C2705 a_6547_4086# a_6983_4478# 0.00412f
C2706 VDD a_4368_4775# 0.453f
C2707 a_6846_4086# a_6505_4394# 1.25e-19
C2708 a_9238_4086# x7.X 3.21e-20
C2709 a_2289_4801# a_1511_4112# 0.00374f
C2710 x4.X a_8696_2366# 0.112f
C2711 VDD a_11544_4775# 0.449f
C2712 x7.X a_11833_2340# 0.00593f
C2713 a_6011_4801# check[5] 1.26e-20
C2714 a_9639_4775# a_10345_3239# 4.94e-20
C2715 D[0] a_8402_3239# 0.00637f
C2716 x5.A a_2853_5648# 1.67e-20
C2717 a_7246_3213# a_6844_2640# 3.43e-19
C2718 check[1] a_4658_4086# 4.01e-21
C2719 a_6759_3213# a_6845_2340# 2.19e-19
C2720 check[4] a_10795_4801# 0.164f
C2721 x72.Q_N a_7953_3239# 0.178f
C2722 a_1061_4801# a_2289_4801# 0.0334f
C2723 x4.X a_1508_5167# 0.138f
C2724 a_1682_4775# a_1976_4775# 0.198f
C2725 a_1227_4801# a_2463_4775# 0.0267f
C2726 a_3600_4086# a_4155_4086# 0.197f
C2727 a_3505_4086# a_4453_4386# 8.38e-21
C2728 a_1511_4112# a_4454_4086# 7.27e-20
C2729 x4.X a_11194_2366# 3.78e-20
C2730 check[2] a_11630_4086# 1.95e-19
C2731 x4.X x75.Q_N 0.00464f
C2732 a_3900_5167# x27.Q_N 8.65e-20
C2733 a_4368_4775# a_5089_5083# 0.00185f
C2734 check[2] a_9638_3213# 0.0022f
C2735 x5.X x33.Q_N 0.00113f
C2736 check[6] a_5896_2340# 0.00282f
C2737 a_11630_4086# a_10628_3239# 6.54e-20
C2738 a_11629_4386# a_10794_3239# 4.11e-20
C2739 a_10776_4086# a_11543_3213# 8.83e-19
C2740 a_11331_4086# a_11249_3213# 1.02e-19
C2741 a_11089_4112# a_11075_3605# 1.61e-19
C2742 x30.Q_N a_5844_3239# 2.88e-19
C2743 a_6606_4801# a_6759_3213# 1.61e-20
C2744 a_6546_2340# a_6845_2340# 0.0334f
C2745 a_9151_3213# a_10794_3239# 1.89e-19
C2746 a_6304_2366# a_7049_2340# 0.199f
C2747 a_9638_3213# a_10628_3239# 0.00116f
C2748 check[0] x30.Q_N 0.00106f
C2749 a_5991_2340# a_7317_2550# 4.7e-22
C2750 a_3452_3239# a_6198_3239# 3.65e-21
C2751 a_4367_3213# a_6291_3605# 4.38e-20
C2752 a_4680_3239# a_6010_3239# 5.35e-20
C2753 a_9151_3213# a_9872_3521# 0.00185f
C2754 x4.X a_3913_4112# 0.112f
C2755 a_11076_5167# x36.Q_N 1.74e-20
C2756 a_11544_4775# a_12265_5083# 0.00185f
C2757 VDD a_8897_4394# 0.00506f
C2758 x4.X a_11195_4112# 0.00334f
C2759 a_4453_4386# x45.Q_N 2.05e-19
C2760 a_9710_4296# a_10156_4112# 0.0367f
C2761 a_9237_4386# a_9377_4112# 0.00126f
C2762 a_8939_4086# a_9578_4112# 0.00316f
C2763 VDD a_7363_4801# 0.0101f
C2764 VDD a_7072_3239# 0.18f
C2765 check[2] a_9236_2640# 8.03e-20
C2766 check[6] a_7073_4801# 4.06e-20
C2767 a_8384_4086# a_8857_3213# 2.45e-19
C2768 a_8697_4112# a_8402_3239# 4.9e-19
C2769 x33.Q_N a_9237_4386# 0.0344f
C2770 a_11331_4086# a_10775_2340# 1.3e-22
C2771 a_11089_4112# a_11088_2366# 1.8e-19
C2772 a_8998_4801# x42.Q_N 2.35e-19
C2773 x20.Q_N x51.Q_N 4.6e-19
C2774 D[4] a_8696_2366# 8.79e-19
C2775 a_9465_4801# check[4] 1.08e-19
C2776 eob a_1822_4801# 0.00828f
C2777 x33.Q_N a_11629_2340# 7.03e-21
C2778 a_2853_5648# x27.D 3.86e-19
C2779 check[0] a_3373_5674# 0.0228f
C2780 check[2] a_2463_4775# 7.62e-20
C2781 a_2389_5648# a_2289_4801# 0.0019f
C2782 x7.X a_4112_2648# 1.53e-19
C2783 a_1822_4801# x4.A 2.88e-19
C2784 VDD a_6845_2340# 0.784f
C2785 a_5992_4086# a_5844_3239# 8.29e-19
C2786 a_4454_4086# a_4154_2340# 3.47e-21
C2787 a_4453_4386# a_4452_2640# 1.32e-20
C2788 a_4658_4086# a_3912_2366# 7.14e-22
C2789 check[0] a_5992_4086# 0.0142f
C2790 a_8384_4086# a_8383_2340# 5.27e-19
C2791 a_11544_4775# a_11331_4086# 3.72e-19
C2792 a_10795_4801# a_11834_4086# 0.00221f
C2793 a_11250_4775# a_11630_4086# 0.00336f
C2794 a_12031_4775# a_11089_4112# 0.00161f
C2795 a_11249_3213# a_11194_2366# 5.71e-21
C2796 a_8938_2340# a_9577_2366# 0.00316f
C2797 check[1] x5.X 0.767f
C2798 a_9236_2640# a_9376_2366# 0.00126f
C2799 a_8696_2366# a_10775_2340# 6.25e-21
C2800 a_3618_3239# a_3899_3605# 0.152f
C2801 a_3452_3239# a_4367_3213# 0.125f
C2802 check[1] a_6292_5167# 1.94e-19
C2803 check[2] a_4453_4386# 1.41e-20
C2804 a_1062_5674# a_1338_5674# 0.00202f
C2805 eob a_621_4112# 9.72e-19
C2806 VDD a_10155_2366# 0.109f
C2807 x4.X a_4657_2340# 0.0013f
C2808 VDD a_6606_4801# 0.0332f
C2809 VDD a_3899_3605# 0.182f
C2810 a_4318_5083# check[6] 1.19e-21
C2811 x45.Q_N D[0] 0.00168f
C2812 VDD a_12264_3521# 0.00506f
C2813 a_621_4112# x4.A 6.66e-19
C2814 reset a_1511_4112# 1.58e-19
C2815 x3.A a_897_4112# 0.3f
C2816 a_11195_4112# a_11249_3213# 3.34e-20
C2817 x27.Q_N a_6844_2640# 1.07e-20
C2818 a_10775_2340# a_11194_2366# 0.0397f
C2819 a_11088_2366# a_11766_2732# 0.00652f
C2820 a_11330_2340# a_11564_2732# 0.00976f
C2821 check[4] a_8802_2366# 1.3e-19
C2822 check[5] a_9102_5083# 8.63e-22
C2823 check[1] a_9237_4386# 1.6e-19
C2824 a_11494_5083# check[3] 2.79e-19
C2825 x4.X x7.A 5.72e-19
C2826 x5.X a_7050_4086# 9.61e-19
C2827 x4.X D[4] 5.2e-19
C2828 x4.X a_11249_3213# 0.00509f
C2829 a_6760_4775# a_6846_4086# 4.63e-19
C2830 a_2289_4801# a_3619_4801# 5.38e-20
C2831 a_7247_4775# a_6845_4386# 6.17e-19
C2832 a_9237_4386# a_9954_4112# 0.0019f
C2833 a_6011_4801# x45.Q_N 7.77e-20
C2834 VDD a_10346_4801# 0.192f
C2835 x4.X x69.Q_N 0.00454f
C2836 a_2463_4775# x20.Q_N 0.129f
C2837 check[5] a_7317_2550# 0.00103f
C2838 x27.Q_N a_4073_3213# 4.88e-19
C2839 a_7246_3213# a_9151_3213# 3.71e-20
C2840 a_4452_2640# x54.Q_N 5.46e-21
C2841 a_4453_2340# a_4925_2550# 0.15f
C2842 VDD a_2784_5996# 0.00533f
C2843 x36.Q_N a_12146_3239# 0.00341f
C2844 VDD a_5897_4086# 0.189f
C2845 x4.X a_7186_4112# 0.00311f
C2846 x36.Q_N a_11761_3239# 4.03e-19
C2847 a_6305_4112# x42.Q_N 5.52e-21
C2848 a_4368_4775# a_3913_4112# 5.67e-20
C2849 a_3619_4801# a_4454_4086# 1.18e-19
C2850 a_4074_4775# a_4453_4386# 3.92e-19
C2851 a_3453_4801# a_4658_4086# 6.96e-19
C2852 a_3900_5167# a_4155_4086# 2.46e-20
C2853 a_6846_4086# a_9238_4086# 1.37e-19
C2854 x4.X a_10775_2340# 0.11f
C2855 x20.Q_N a_4453_4386# 1.28e-19
C2856 x45.Q_N a_5561_3239# 1.19e-20
C2857 a_6978_4801# check[5] 1.84e-20
C2858 a_8402_3239# a_10345_3239# 7.94e-21
C2859 D[5] a_7049_2340# 7e-20
C2860 a_8236_3239# D[1] 7.04e-20
C2861 D[7] a_2060_2640# 1.7e-19
C2862 a_1112_2340# a_2061_2340# 1.03e-19
C2863 D[0] a_9369_3239# 5.51e-20
C2864 check[4] a_11762_4801# 5.42e-20
C2865 x77.Y a_4538_3521# 2.52e-20
C2866 a_6305_4112# x7.X 2.29e-20
C2867 a_1061_4801# a_3807_4801# 3.65e-21
C2868 x4.X a_4368_4775# 0.101f
C2869 a_1338_5674# x5.X 0.225f
C2870 check[2] a_6011_4801# 1.18e-19
C2871 x27.Q_N a_5372_4112# 0.0147f
C2872 x4.X a_11544_4775# 0.105f
C2873 VDD x51.Q_N 0.085f
C2874 check[2] a_11543_3213# 1.77e-20
C2875 x39.Q_N a_11714_3521# 0.00203f
C2876 a_10628_3239# a_11543_3213# 0.126f
C2877 a_10794_3239# a_11075_3605# 0.155f
C2878 a_7317_2550# a_7185_2366# 0.0258f
C2879 a_6844_2640# a_8938_2340# 3.87e-20
C2880 a_4854_3213# a_5371_2366# 2.38e-19
C2881 a_6845_2340# a_8696_2366# 3.1e-19
C2882 check[1] a_9656_4394# 1.56e-20
C2883 x30.Q_N a_6399_3239# 6.75e-20
C2884 x30.Q_N x33.Q_N 2.51e-20
C2885 a_4213_3239# a_4789_3239# 2.46e-21
C2886 x5.X a_7764_4112# 9.62e-19
C2887 VDD a_11630_4086# 0.809f
C2888 check[2] a_8697_4112# 0.00313f
C2889 VDD a_9638_3213# 0.569f
C2890 a_3170_4801# a_3453_4801# 8.18e-19
C2891 check[2] a_11330_2340# 0.00111f
C2892 x20.Q_N x54.Q_N 1.47e-19
C2893 a_9441_2340# a_9374_2732# 9.46e-19
C2894 a_8696_2366# a_10155_2366# 4.94e-21
C2895 x60.Q_N a_8896_2648# 2.02e-20
C2896 x30.Q_N a_6780_2366# 9.42e-19
C2897 a_9236_2640# a_9655_2648# 2.46e-19
C2898 a_10794_3239# a_11088_2366# 5.94e-19
C2899 a_11249_3213# a_10775_2340# 2.5e-19
C2900 x4.X a_8897_4394# 1.75e-19
C2901 x5.X a_3453_4801# 0.255f
C2902 check[2] a_4681_4801# 4.32e-20
C2903 x4.X a_7363_4801# 0.00557f
C2904 x4.X a_7072_3239# 0.00457f
C2905 VDD a_9236_2640# 0.269f
C2906 x45.Q_N a_6375_3605# 8.49e-19
C2907 x5.X a_10629_4801# 0.27f
C2908 a_8403_4801# a_8858_4775# 0.153f
C2909 a_8237_4801# a_8684_5167# 0.15f
C2910 a_1520_2366# a_3504_2340# 9.77e-21
C2911 a_1207_2340# a_1996_2366# 4.2e-20
C2912 a_10680_2340# a_11629_2340# 1.03e-19
C2913 check[4] a_8383_2340# 2.57e-20
C2914 x36.Q_N a_11629_4386# 0.0351f
C2915 a_11390_4801# x39.Q_N 2.02e-19
C2916 a_11250_4775# a_11543_3213# 7.57e-21
C2917 a_10629_4801# a_11856_3239# 4.76e-21
C2918 eob a_1520_2366# 1.28e-19
C2919 a_4367_3213# a_5088_3521# 0.00185f
C2920 check[1] x30.Q_N 0.0373f
C2921 VDD a_2463_4775# 0.704f
C2922 a_1227_4801# a_897_4112# 4.21e-19
C2923 x48.Q a_4113_4394# 5.88e-19
C2924 x48.Q x7.X 3.3e-20
C2925 VDD a_12345_2732# 0.0042f
C2926 x4.X a_6845_2340# 0.00277f
C2927 a_4971_4801# a_4926_4296# 1.9e-20
C2928 x48.Q a_4539_5083# 6.59e-19
C2929 x4.A a_1520_2366# 6.86e-19
C2930 a_4453_4386# a_3618_3239# 4.11e-20
C2931 a_3913_4112# a_3899_3605# 1.61e-19
C2932 a_3600_4086# a_4367_3213# 8.83e-19
C2933 a_4454_4086# a_3452_3239# 6.54e-20
C2934 a_4155_4086# a_4073_3213# 1.02e-19
C2935 x45.Q_N a_7317_2550# 0.00196f
C2936 a_3599_2340# a_4112_2648# 0.00945f
C2937 a_7246_3213# a_7953_3239# 0.0968f
C2938 a_6759_3213# D[0] 4.66e-19
C2939 VDD a_4453_4386# 0.593f
C2940 check[2] a_9375_4478# 1.05e-20
C2941 VDD a_12346_4478# 0.0042f
C2942 x4.X a_10155_2366# 7.73e-20
C2943 x4.X a_6606_4801# 7.25e-19
C2944 x4.X a_11965_3239# 1.05e-19
C2945 a_3453_4801# a_3984_5167# 0.0018f
C2946 a_4074_4775# a_4681_4801# 0.00187f
C2947 a_3900_5167# a_4855_4775# 4.7e-22
C2948 a_3619_4801# a_3807_4801# 0.162f
C2949 x4.X a_3899_3605# 0.018f
C2950 x4.X a_12264_3521# 0.00103f
C2951 a_10776_4086# a_12102_4296# 4.7e-22
C2952 a_9578_4112# x39.Q_N 5.6e-20
C2953 a_1822_4801# a_2398_4801# 2.46e-21
C2954 check[2] a_9102_5083# 1.52e-19
C2955 a_11331_4086# a_11630_4086# 0.0334f
C2956 a_11089_4112# a_11834_4086# 0.199f
C2957 x5.X a_9639_4775# 0.00985f
C2958 x20.Q_N a_4681_4801# 2.69e-20
C2959 check[1] a_3373_5674# 0.027f
C2960 a_2853_5648# a_3876_6040# 0.00747f
C2961 x45.Q_N a_4854_3213# 1.37e-20
C2962 a_6011_4801# a_6759_3213# 2.05e-21
C2963 a_6292_5167# a_6465_3213# 3.52e-21
C2964 a_7247_4775# a_8684_5167# 7.98e-21
C2965 a_6466_4775# a_6291_3605# 1.33e-23
C2966 check[1] a_5992_4086# 5.87e-20
C2967 a_8402_3239# a_8590_3239# 0.163f
C2968 a_8857_3213# a_9464_3239# 0.00187f
C2969 a_8683_3605# a_9638_3213# 4.7e-22
C2970 a_8236_3239# a_8767_3605# 0.0018f
C2971 a_3258_5648# a_1511_4112# 3.06e-19
C2972 a_10629_4801# a_11160_5167# 0.0018f
C2973 a_10795_4801# a_10983_4801# 0.162f
C2974 a_11250_4775# a_11857_4801# 0.00187f
C2975 a_6605_3239# a_7181_3239# 2.46e-21
C2976 a_11076_5167# a_12031_4775# 4.7e-22
C2977 sel_bit[1] a_1511_4112# 3.24e-20
C2978 a_3600_4086# a_4389_4112# 4.2e-20
C2979 a_4453_4386# a_5170_4478# 4.45e-20
C2980 a_4454_4086# a_4872_4394# 0.00276f
C2981 x4.X a_10346_4801# 0.0067f
C2982 x27.Q_N a_4155_4086# 1.3e-22
C2983 clk_sar a_897_4112# 1.96e-20
C2984 check[2] a_10345_3239# 0.00302f
C2985 a_8403_4801# x42.Q_N 7.79e-20
C2986 a_9639_4775# a_9237_4386# 6.17e-19
C2987 a_9152_4775# a_9238_4086# 4.63e-19
C2988 a_9578_4112# a_9709_2550# 1.72e-22
C2989 a_3373_5674# a_3877_5674# 5.33e-19
C2990 sel_bit[1] a_1061_4801# 7.04e-20
C2991 a_7049_2340# a_7763_2366# 6.99e-20
C2992 a_6845_2340# D[4] 0.336f
C2993 a_7317_2550# a_7561_2732# 0.00972f
C2994 a_10345_3239# a_10628_3239# 8.18e-19
C2995 a_9638_3213# a_8696_2366# 8.4e-19
C2996 a_8402_3239# a_9441_2340# 0.00154f
C2997 a_9151_3213# a_8938_2340# 2.17e-19
C2998 a_5561_3239# a_6759_3213# 5.62e-20
C2999 a_8857_3213# a_9237_2340# 0.00199f
C3000 a_4854_3213# a_4452_2640# 3.43e-19
C3001 a_4367_3213# a_4453_2340# 2.19e-19
C3002 x33.Q_N x60.Q_N 4.08e-19
C3003 x4.X a_5897_4086# 0.00454f
C3004 a_4593_4112# x45.Q_N 3.1e-20
C3005 a_6547_4086# a_6845_4386# 0.137f
C3006 a_6305_4112# a_6846_4086# 0.125f
C3007 VDD D[0] 0.301f
C3008 check[1] eob 0.00405f
C3009 a_8403_4801# x7.X 2.9e-21
C3010 VDD x54.Q_N 0.0807f
C3011 a_6466_4775# a_6710_5083# 0.0104f
C3012 a_6011_4801# a_6931_5083# 1.09e-19
C3013 x30.Q_N a_6410_2366# 0.0102f
C3014 a_8383_2340# a_9237_2340# 0.0492f
C3015 a_8696_2366# a_9236_2640# 0.139f
C3016 a_9152_4775# a_9755_4801# 0.0552f
C3017 a_9754_3239# a_9573_3239# 4.11e-20
C3018 sel_bit[0] a_621_4112# 8.01e-21
C3019 a_10794_3239# x66.Q_N 3.85e-21
C3020 a_11856_3239# a_11942_3605# 0.00976f
C3021 VDD a_6011_4801# 0.593f
C3022 x4.X x51.Q_N 0.0098f
C3023 VDD a_11543_3213# 0.352f
C3024 x7.X a_5896_2340# 7.85e-19
C3025 a_4454_4086# D[5] 1.26e-20
C3026 a_11834_4086# a_11767_4478# 9.46e-19
C3027 a_10776_4086# a_11565_4112# 4.2e-20
C3028 VDD a_11966_4801# 7.87e-19
C3029 x30.Q_N a_7764_4112# 0.0147f
C3030 x39.Q_N a_11289_4394# 2.02e-20
C3031 a_11629_4386# a_12048_4394# 2.46e-19
C3032 x42.Q_N a_9754_3239# 0.00969f
C3033 a_1762_2340# a_1996_2732# 0.00976f
C3034 a_1207_2340# a_1626_2366# 0.0397f
C3035 a_1520_2366# a_2198_2732# 0.00652f
C3036 x27.Q_N a_4925_2550# 0.181f
C3037 a_9236_2640# a_11194_2366# 2.19e-20
C3038 a_10155_2366# a_10775_2340# 8.26e-21
C3039 check[4] a_10794_3239# 1.18e-19
C3040 a_2389_5648# a_3258_5648# 0.0296f
C3041 sel_bit[0] check[0] 0.163f
C3042 a_2853_5648# x48.Q 0.016f
C3043 x77.Y a_5844_3239# 2.13e-19
C3044 a_3618_3239# a_5561_3239# 3.23e-21
C3045 a_3452_3239# x75.Q 6.31e-20
C3046 check[0] x77.Y 2.24e-20
C3047 a_2389_5648# sel_bit[1] 0.0628f
C3048 VDD a_8697_4112# 0.448f
C3049 check[1] x60.Q_N 0.0122f
C3050 x4.X a_11630_4086# 0.0441f
C3051 x4.X a_9638_3213# 0.116f
C3052 VDD a_5561_3239# 0.19f
C3053 VDD a_11330_2340# 0.177f
C3054 a_9710_4296# x42.Q_N 0.00244f
C3055 x45.Q_N a_8590_3239# 1.34e-20
C3056 a_7050_4086# a_7362_3239# 5.48e-21
C3057 x27.Q_N a_5845_4801# 4.37e-19
C3058 D[6] a_2777_2366# 1.54e-19
C3059 a_4681_4801# a_3618_3239# 6.75e-21
C3060 x5.X a_11184_4801# 2.88e-19
C3061 a_2200_2366# a_2401_2366# 3.34e-19
C3062 a_3504_2340# a_3912_2366# 6.04e-19
C3063 x20.Q_N D[7] 5.48e-19
C3064 a_8858_4775# a_9370_4801# 9.75e-19
C3065 a_8684_5167# a_8792_4801# 0.00812f
C3066 a_8237_4801# x33.Q_N 1.26e-19
C3067 a_6010_3239# a_6709_3521# 2.46e-19
C3068 a_9465_4801# a_9323_5083# 0.00412f
C3069 check[4] a_9577_2366# 4.82e-19
C3070 a_9639_4775# a_9551_5167# 7.71e-20
C3071 a_9152_4775# a_8998_4801# 0.00943f
C3072 a_5844_3239# a_6930_3521# 0.00907f
C3073 x36.Q_N a_11075_3605# 0.00192f
C3074 x48.Q a_3671_5674# 0.0017f
C3075 x36.Q_N a_12147_4801# 3.8e-19
C3076 VDD a_4681_4801# 0.346f
C3077 a_6846_4086# a_6983_4478# 0.00907f
C3078 x45.Q_N a_5170_4112# 3.4e-20
C3079 x4.X a_9236_2640# 0.00898f
C3080 x5.X check[5] 0.17f
C3081 VDD a_11857_4801# 0.343f
C3082 x7.X x63.Q_N 2.11e-19
C3083 check[6] a_5844_3239# 0.00782f
C3084 a_6292_5167# check[5] 7.62e-21
C3085 check[0] check[6] 0.45f
C3086 a_6760_4775# a_7954_4801# 6.04e-19
C3087 a_1338_5674# eob 9.5e-19
C3088 a_7953_3239# a_9151_3213# 5.62e-20
C3089 D[0] a_8683_3605# 2.17e-19
C3090 a_7246_3213# a_7049_2340# 2.52e-19
C3091 a_6759_3213# a_7317_2550# 1.62e-19
C3092 check[4] a_11076_5167# 0.0011f
C3093 a_3373_5674# a_3453_4801# 1.45e-21
C3094 x36.Q_N a_11088_2366# 0.0928f
C3095 a_1061_4801# a_1592_5167# 0.0018f
C3096 a_1227_4801# a_1415_4801# 0.163f
C3097 x4.X a_2463_4775# 0.148f
C3098 a_1682_4775# a_2289_4801# 0.00187f
C3099 a_2969_6040# x20.Q_N 1.2e-20
C3100 a_3600_4086# a_4454_4086# 0.0492f
C3101 a_1338_5674# x4.A 7.27e-19
C3102 a_3913_4112# a_4453_4386# 0.139f
C3103 a_4855_4775# a_5372_4112# 4.23e-19
C3104 x4.X a_12345_2732# 1.17e-19
C3105 x5.X a_10776_4086# 0.0184f
C3106 check[2] a_12102_4296# 4.54e-20
C3107 a_4855_4775# x27.Q_N 0.128f
C3108 check[6] a_4592_2366# 8.47e-20
C3109 a_11834_4086# a_10794_3239# 2.9e-19
C3110 a_11089_4112# a_12030_3213# 9.49e-19
C3111 a_11331_4086# a_11543_3213# 2.12e-19
C3112 a_11630_4086# a_11249_3213# 5.04e-19
C3113 a_12147_4801# a_11629_4386# 8.84e-21
C3114 D[0] a_8696_2366# 3.91e-20
C3115 x30.Q_N a_6465_3213# 5.84e-19
C3116 a_8236_3239# a_10982_3239# 3.65e-21
C3117 a_6844_2640# a_7049_2340# 0.153f
C3118 a_9151_3213# a_11075_3605# 4.38e-20
C3119 a_6304_2366# x57.Q_N 0.00553f
C3120 a_9464_3239# a_10794_3239# 3.48e-20
C3121 a_4854_3213# a_6759_3213# 3.71e-20
C3122 a_9638_3213# x69.Q_N 0.124f
C3123 x4.X a_4453_4386# 0.0483f
C3124 check[1] a_8237_4801# 0.00245f
C3125 a_12031_4775# x36.Q_N 0.126f
C3126 VDD a_9375_4478# 0.0163f
C3127 x4.X a_12346_4478# 9.15e-19
C3128 a_4658_4086# x45.Q_N 3.93e-20
C3129 VDD a_9102_5083# 0.00984f
C3130 a_9237_4386# a_10776_4086# 1.52e-19
C3131 a_9238_4086# a_9578_4112# 6.04e-20
C3132 VDD a_6375_3605# 0.0042f
C3133 x42.Q_N a_10681_4086# 1.37e-20
C3134 a_9442_4086# a_9377_4112# 9.75e-19
C3135 a_9237_4386# a_8402_3239# 4.11e-20
C3136 a_8697_4112# a_8683_3605# 1.61e-19
C3137 a_8939_4086# a_8857_3213# 1.02e-19
C3138 a_8384_4086# a_9151_3213# 8.83e-19
C3139 a_9238_4086# a_8236_3239# 6.54e-20
C3140 a_11629_4386# a_11088_2366# 1.93e-22
C3141 x30.Q_N a_5991_2340# 0.142f
C3142 a_7763_2366# a_9237_2340# 3.65e-21
C3143 eob a_3453_4801# 5.9e-20
C3144 x75.Q D[5] 9.96e-19
C3145 D[4] a_9236_2640# 3.87e-20
C3146 eob a_2194_4801# 0.00151f
C3147 D[1] a_11389_3239# 1.6e-19
C3148 VDD a_897_4112# 0.418f
C3149 a_10681_4086# x7.X 2.05e-21
C3150 VDD a_10345_3239# 0.19f
C3151 x7.X a_4590_2732# 9.45e-19
C3152 VDD a_7317_2550# 0.172f
C3153 a_6305_4112# a_6010_3239# 4.9e-19
C3154 check[2] a_11564_2366# 1.34e-19
C3155 a_5992_4086# a_6465_3213# 2.45e-19
C3156 a_4454_4086# a_4453_2340# 1.55e-19
C3157 a_4453_4386# a_4657_2340# 1.26e-21
C3158 check[0] a_6547_4086# 3.86e-19
C3159 a_8939_4086# a_8383_2340# 1.3e-22
C3160 a_8697_4112# a_8696_2366# 1.8e-19
C3161 a_12031_4775# a_11629_4386# 6.17e-19
C3162 a_10795_4801# x39.Q_N 7.79e-20
C3163 a_11544_4775# a_11630_4086# 4.63e-19
C3164 a_9236_2640# a_10775_2340# 3.6e-19
C3165 a_9237_2340# a_9577_2366# 6.04e-20
C3166 a_9441_2340# a_9376_2366# 9.75e-19
C3167 a_3452_3239# a_4680_3239# 0.0334f
C3168 a_3618_3239# a_4854_3213# 0.0264f
C3169 a_4073_3213# a_4367_3213# 0.198f
C3170 check[1] a_7247_4775# 0.0127f
C3171 x33.Q_N a_9574_4801# 7.27e-21
C3172 a_1227_4801# a_3170_4801# 1.76e-19
C3173 a_1061_4801# x27.D 5.94e-20
C3174 a_1062_5674# check[2] 7.36e-19
C3175 check[2] a_4658_4086# 4.4e-21
C3176 x5.X a_3505_4086# 0.00259f
C3177 x5.A a_2389_5648# 4.35e-20
C3178 clk_sar a_1062_5674# 0.185f
C3179 VDD a_6978_4801# 0.00445f
C3180 x4.X D[0] 0.0011f
C3181 x5.X a_11565_4478# 1.76e-19
C3182 x4.X x54.Q_N 0.00996f
C3183 VDD D[7] 0.225f
C3184 a_5992_4086# a_5991_2340# 5.27e-19
C3185 VDD a_4854_3213# 0.572f
C3186 D[6] a_3504_2340# 0.103f
C3187 a_2060_2640# a_2777_2366# 0.0019f
C3188 x27.Q_N a_7049_2340# 8.08e-21
C3189 a_11628_2640# a_11766_2732# 1.09e-19
C3190 a_11088_2366# a_12047_2648# 1.21e-20
C3191 a_11330_2340# a_11194_2366# 0.0282f
C3192 check[1] a_9442_4086# 1.18e-19
C3193 x5.X a_1227_4801# 0.0165f
C3194 eob D[6] 8.49e-20
C3195 x75.Q_N a_5561_3239# 0.178f
C3196 a_11943_5167# check[3] 4.39e-19
C3197 x4.X a_6011_4801# 0.00494f
C3198 x5.X x45.Q_N 0.00731f
C3199 x4.X a_11543_3213# 0.111f
C3200 a_6760_4775# a_7318_4296# 2.85e-19
C3201 a_7247_4775# a_7050_4086# 4.44e-19
C3202 a_6292_5167# x45.Q_N 9.97e-20
C3203 x4.X a_11966_4801# 2.39e-19
C3204 a_1415_4801# x20.Q_N 5.43e-21
C3205 a_8803_4112# a_8857_3213# 3.34e-20
C3206 x27.Q_N a_6400_4801# 2.58e-20
C3207 x33.Q_N a_10156_4112# 0.0147f
C3208 VDD a_3648_5972# 0.0123f
C3209 x27.Q_N a_4367_3213# 0.00484f
C3210 a_7246_3213# a_9464_3239# 1.86e-21
C3211 a_6759_3213# a_8590_3239# 3.42e-20
C3212 VDD a_2969_6040# 0.00654f
C3213 x36.Q_N D[3] 0.00274f
C3214 VDD a_4593_4112# 0.00494f
C3215 x4.X a_8697_4112# 0.109f
C3216 x36.Q_N x66.Q_N 0.02f
C3217 a_4368_4775# a_4453_4386# 7.46e-19
C3218 a_3807_4801# a_3600_4086# 3.44e-19
C3219 a_2579_4801# a_1511_4112# 3.99e-19
C3220 a_4681_4801# a_3913_4112# 3.76e-19
C3221 check[2] a_3170_4801# 1.57e-20
C3222 a_6845_4386# x42.Q_N 1.95e-19
C3223 x20.Q_N a_4658_4086# 2.19e-20
C3224 x4.X a_11330_2340# 0.0071f
C3225 x4.X a_5561_3239# 0.00286f
C3226 check[0] a_6411_4112# 4.09e-19
C3227 x30.Q_N check[5] 0.902f
C3228 D[0] D[4] 0.338f
C3229 a_8857_3213# D[1] 1.23e-20
C3230 D[5] x57.Q_N 0.00107f
C3231 D[7] a_2265_2340# 2.67e-19
C3232 check[4] x36.Q_N 8.5e-21
C3233 x77.Y a_4213_3239# 0.0313f
C3234 x4.X a_4681_4801# 0.00584f
C3235 sel_bit[0] check[1] 0.583f
C3236 a_6845_4386# x7.X 2.52e-20
C3237 check[2] x5.X 0.832f
C3238 clk_sar x5.X 0.00873f
C3239 check[2] a_6292_5167# 5.02e-20
C3240 x4.X a_11857_4801# 0.00316f
C3241 x5.X a_10628_3239# 9.1e-20
C3242 x20.Q_N a_1720_2648# 2.75e-19
C3243 a_11834_4086# a_12146_3239# 5.48e-21
C3244 x30.Q_N a_5371_2366# 1.34e-20
C3245 a_8237_4801# a_10629_4801# 0.00176f
C3246 a_9638_3213# a_10155_2366# 2.38e-19
C3247 x30.Q_N a_8402_3239# 3.97e-20
C3248 x39.Q_N a_11389_3239# 0.0314f
C3249 a_621_4112# comparator_out 2.33e-19
C3250 a_6844_2640# a_9237_2340# 2.9e-21
C3251 a_10628_3239# a_11856_3239# 0.0334f
C3252 a_6845_2340# a_9236_2640# 4e-20
C3253 a_10794_3239# a_12030_3213# 0.0264f
C3254 a_7317_2550# a_8696_2366# 6.06e-21
C3255 a_11249_3213# a_11543_3213# 0.199f
C3256 x69.Q_N a_11543_3213# 2.97e-20
C3257 check[2] a_9237_4386# 0.163f
C3258 VDD a_12102_4296# 0.317f
C3259 sel_bit[0] a_3877_5674# 2.93e-19
C3260 x27.D a_3619_4801# 0.159f
C3261 VDD a_8590_3239# 0.109f
C3262 a_10156_4112# a_9954_4112# 3.67e-19
C3263 a_7247_4775# a_7764_4112# 4.23e-19
C3264 x48.Q a_4971_4801# 4.12e-19
C3265 x20.Q_N a_3170_4801# 0.187f
C3266 a_2697_5083# x27.D 7.73e-21
C3267 check[2] a_11629_2340# 1.99e-19
C3268 x42.Q_N a_9322_3521# 0.00203f
C3269 a_9441_2340# a_9655_2648# 0.0104f
C3270 a_9237_2340# a_9953_2732# 0.0018f
C3271 x30.Q_N a_7185_2366# 0.0403f
C3272 a_9236_2640# a_10155_2366# 0.159f
C3273 a_11249_3213# a_11330_2340# 4.18e-20
C3274 a_11075_3605# a_11088_2366# 1.71e-19
C3275 a_11543_3213# a_10775_2340# 9.06e-19
C3276 check[4] a_9151_3213# 1.06e-19
C3277 a_10794_3239# a_11628_2640# 4.04e-20
C3278 a_10346_4801# a_9638_3213# 3.19e-20
C3279 a_10628_3239# a_11629_2340# 6.52e-20
C3280 check[1] check[6] 6.18e-20
C3281 eob x3.A 0.00121f
C3282 VDD a_5170_4112# 1.14e-19
C3283 x4.X a_9375_4478# 0.00114f
C3284 x5.X a_4074_4775# 3.66e-19
C3285 a_2389_5648# a_2579_4801# 2.13e-20
C3286 a_8289_4086# a_9238_4086# 7e-20
C3287 x7.X a_6780_2732# 1.8e-19
C3288 x4.X a_6375_3605# 9.07e-19
C3289 x5.X x20.Q_N 0.00434f
C3290 a_4368_4775# a_6011_4801# 1.1e-19
C3291 a_4855_4775# a_5845_4801# 0.00116f
C3292 VDD a_9441_2340# 0.304f
C3293 x3.A x4.A 4.66e-19
C3294 x5.X a_11250_4775# 0.00324f
C3295 a_8237_4801# a_9639_4775# 0.0492f
C3296 a_8403_4801# a_9152_4775# 0.139f
C3297 a_8858_4775# a_8684_5167# 0.205f
C3298 a_1520_2366# a_2200_2366# 3.73e-19
C3299 a_1762_2340# a_1996_2366# 0.00707f
C3300 a_2060_2640# a_3504_2340# 6.83e-19
C3301 check[4] a_8938_2340# 1.33e-19
C3302 a_10775_2340# a_11330_2340# 0.197f
C3303 a_11544_4775# a_11543_3213# 0.00121f
C3304 x77.Y a_3912_2366# 7.49e-20
C3305 a_11544_4775# a_11966_4801# 2.87e-21
C3306 a_12031_4775# a_12147_4801# 0.0397f
C3307 eob a_2060_2640# 1.44e-19
C3308 a_4854_3213# x75.Q_N 0.124f
C3309 x4.X a_897_4112# 1.27e-19
C3310 VDD a_1415_4801# 0.12f
C3311 x48.Q a_4591_4478# 6.11e-19
C3312 x4.X a_10345_3239# 0.00275f
C3313 x4.X a_7317_2550# 0.00147f
C3314 x48.Q a_4214_4801# 0.00132f
C3315 a_1338_5674# sel_bit[0] 0.0571f
C3316 a_4155_4086# a_4367_3213# 2.12e-19
C3317 a_4658_4086# a_3618_3239# 2.9e-19
C3318 a_4454_4086# a_4073_3213# 5.04e-19
C3319 a_3913_4112# a_4854_3213# 9.49e-19
C3320 a_3912_2366# a_4388_2732# 0.00133f
C3321 a_7072_3239# D[0] 5.18e-20
C3322 VDD a_4658_4086# 0.489f
C3323 VDD a_1062_5674# 0.234f
C3324 x36.Q_N a_9237_2340# 1.55e-19
C3325 VDD a_11565_4112# 3.47e-19
C3326 check[2] a_9656_4394# 7.77e-21
C3327 x4.X a_6978_4801# 5.55e-19
C3328 a_3619_4801# a_2579_4801# 7.73e-20
C3329 x4.X a_4854_3213# 0.117f
C3330 a_4074_4775# a_3984_5167# 6.69e-20
C3331 x4.X D[7] 0.00353f
C3332 a_3900_5167# a_3807_4801# 0.0367f
C3333 a_4368_4775# a_4681_4801# 0.124f
C3334 x5.X a_8591_4801# 0.00545f
C3335 x30.Q_N x45.Q_N 0.0041f
C3336 check[2] a_9551_5167# 1.87e-19
C3337 a_11089_4112# x39.Q_N 0.0933f
C3338 a_11629_4386# a_11834_4086# 0.153f
C3339 a_2853_5648# a_2993_5674# 1.56e-19
C3340 check[6] a_3912_2366# 1.31e-20
C3341 a_7073_4801# a_6010_3239# 6.75e-21
C3342 check[1] a_6547_4086# 7.52e-20
C3343 check[0] a_7561_2366# 1.87e-20
C3344 D[0] a_6845_2340# 0.0271f
C3345 a_8402_3239# a_7362_3239# 1.22e-20
C3346 a_9151_3213# a_9464_3239# 0.124f
C3347 a_8857_3213# a_8767_3605# 6.69e-20
C3348 a_8683_3605# a_8590_3239# 0.0367f
C3349 a_4453_2340# x57.Q_N 2.94e-19
C3350 a_11250_4775# a_11160_5167# 6.69e-20
C3351 a_11544_4775# a_11857_4801# 0.124f
C3352 a_11076_5167# a_10983_4801# 0.0367f
C3353 a_10795_4801# a_9755_4801# 4.87e-21
C3354 x36.Q_N a_12547_2366# 0.0317f
C3355 eob a_653_3238# 0.0383f
C3356 a_4453_4386# a_5897_4086# 3.56e-19
C3357 a_4658_4086# a_5170_4478# 6.69e-20
C3358 a_4155_4086# a_4389_4112# 0.00707f
C3359 a_4454_4086# a_5372_4112# 0.0664f
C3360 a_3913_4112# a_4593_4112# 3.73e-19
C3361 VDD a_1720_2648# 0.00736f
C3362 a_8384_4086# a_9173_4478# 7.71e-20
C3363 a_8697_4112# a_8897_4394# 0.00185f
C3364 x27.Q_N a_4454_4086# 0.0256f
C3365 a_9152_4775# a_9710_4296# 2.85e-19
C3366 a_897_4112# x7.A 1.11e-19
C3367 a_8684_5167# x42.Q_N 9.99e-20
C3368 a_9639_4775# a_9442_4086# 4.44e-19
C3369 x3.A a_929_3238# 2.98e-19
C3370 sel_bit[0] a_3453_4801# 4.34e-20
C3371 a_3453_4801# x77.Y 9.38e-22
C3372 x30.Q_N a_4452_2640# 0.00116f
C3373 sel_bit[1] a_1682_4775# 6.18e-20
C3374 D[1] a_10794_3239# 0.00642f
C3375 a_9151_3213# a_9237_2340# 2.19e-19
C3376 x36.Q_N a_12548_4112# 0.0133f
C3377 a_9638_3213# a_9236_2640# 3.43e-19
C3378 a_4367_3213# a_4925_2550# 1.62e-19
C3379 x69.Q_N a_10345_3239# 0.178f
C3380 x4.X a_4593_4112# 0.0012f
C3381 a_4854_3213# a_4657_2340# 2.52e-19
C3382 VDD a_3170_4801# 0.212f
C3383 a_6547_4086# a_7050_4086# 0.00187f
C3384 a_5992_4086# x45.Q_N 0.154f
C3385 a_6845_4386# a_6846_4086# 0.75f
C3386 a_6305_4112# a_7318_4296# 0.0633f
C3387 x7.X a_2777_2732# 8.11e-19
C3388 x5.X a_6931_5083# 5.11e-19
C3389 x7.X a_5844_3239# 0.147f
C3390 check[2] x30.Q_N 6.73e-21
C3391 a_3505_4086# a_3504_2340# 1.07e-20
C3392 check[0] x7.X 0.121f
C3393 a_6199_4801# a_6376_5167# 8.94e-19
C3394 a_6760_4775# a_6710_5083# 1.21e-20
C3395 a_7186_4112# a_7317_2550# 1.72e-22
C3396 a_6011_4801# a_6606_4801# 0.00118f
C3397 check[0] a_4539_5083# 4.79e-19
C3398 a_8938_2340# a_9237_2340# 0.0334f
C3399 a_12030_3213# a_12146_3239# 0.0397f
C3400 a_8383_2340# a_9709_2550# 4.7e-22
C3401 a_9465_4801# a_9755_4801# 0.0282f
C3402 a_9639_4775# a_9574_4801# 4.2e-20
C3403 a_11543_3213# a_11965_3239# 2.87e-21
C3404 a_8696_2366# a_9441_2340# 0.199f
C3405 a_11543_3213# a_12264_3521# 0.00185f
C3406 VDD x5.X 2.88f
C3407 VDD a_6292_5167# 0.317f
C3408 a_3453_4801# check[6] 8.06e-20
C3409 a_3619_4801# a_5562_4801# 1.64e-20
C3410 VDD a_11856_3239# 0.18f
C3411 a_11331_4086# a_11565_4112# 0.00707f
C3412 a_11630_4086# a_12346_4478# 0.0018f
C3413 a_11834_4086# a_12048_4394# 0.0104f
C3414 eob a_1227_4801# 0.413f
C3415 a_11629_4386# a_12548_4112# 0.163f
C3416 a_11089_4112# a_11769_4112# 3.73e-19
C3417 a_7954_4801# a_8403_4801# 5.4e-19
C3418 check[5] a_8237_4801# 0.414f
C3419 a_2060_2640# a_2198_2732# 1.09e-19
C3420 a_1762_2340# a_1626_2366# 0.0282f
C3421 a_1520_2366# a_2479_2648# 1.21e-20
C3422 check[1] a_6411_4112# 1.13e-20
C3423 x30.Q_N a_9376_2366# 2.98e-20
C3424 D[3] a_11088_2366# 8.67e-19
C3425 a_12146_3239# a_11628_2640# 5.05e-21
C3426 check[2] a_3373_5674# 0.0404f
C3427 x77.Y D[6] 4.91e-19
C3428 check[4] a_12147_4801# 1.37e-20
C3429 a_10629_4801# check[3] 0.00126f
C3430 a_10795_4801# a_12738_4801# 8.38e-21
C3431 a_1227_4801# x4.A 0.00377f
C3432 check[2] a_5992_4086# 3.43e-20
C3433 VDD a_9237_4386# 0.59f
C3434 x5.X a_5170_4478# 1.85e-19
C3435 x4.X a_12102_4296# 0.021f
C3436 x48.Q a_1511_4112# 0.00368f
C3437 x4.X a_8590_3239# 0.0062f
C3438 x7.X a_8896_2648# 1.53e-19
C3439 a_1976_4775# a_2289_4801# 0.124f
C3440 a_1508_5167# a_1415_4801# 0.0367f
C3441 VDD a_11629_2340# 0.784f
C3442 x27.Q_N a_6466_4775# 1.88e-20
C3443 a_9639_4775# a_10156_4112# 4.23e-19
C3444 a_653_3238# a_929_3238# 0.00202f
C3445 x45.Q_N a_7362_3239# 0.00968f
C3446 x5.X a_12265_5083# 1.33e-19
C3447 a_4368_4775# a_4854_3213# 1.06e-20
C3448 a_4855_4775# a_4367_3213# 1.08e-22
C3449 a_8237_4801# a_8402_3239# 8.16e-19
C3450 a_8403_4801# a_8236_3239# 9.04e-19
C3451 a_11194_2366# a_11564_2366# 4.11e-20
C3452 a_3504_2340# a_4452_2640# 9.65e-21
C3453 x20.Q_N a_3806_3239# 0.00103f
C3454 a_9152_4775# a_9370_4801# 3.73e-19
C3455 a_9465_4801# a_8998_4801# 0.00316f
C3456 a_8858_4775# x33.Q_N 2.07e-20
C3457 a_6010_3239# a_7158_3605# 2.13e-19
C3458 check[4] a_11088_2366# 2.47e-20
C3459 a_6465_3213# a_6930_3521# 9.46e-19
C3460 a_5844_3239# a_6605_3239# 6.04e-20
C3461 x4.X a_5170_4112# 7.21e-19
C3462 x36.Q_N a_12030_3213# 0.0126f
C3463 a_12031_4775# x66.Q_N 4.45e-20
C3464 x48.Q a_1061_4801# 4.14e-21
C3465 a_6846_4086# a_7264_4394# 0.00276f
C3466 a_6845_4386# a_7562_4478# 4.45e-20
C3467 a_5992_4086# a_6781_4112# 4.2e-20
C3468 VDD a_3984_5167# 0.0046f
C3469 x4.X a_9441_2340# 0.00148f
C3470 VDD a_11160_5167# 0.0042f
C3471 a_7247_4775# check[5] 0.0104f
C3472 check[2] eob 0.0123f
C3473 D[0] a_9638_3213# 1.68e-20
C3474 clk_sar eob 4.74e-20
C3475 check[4] a_12031_4775# 1.91e-20
C3476 a_7072_3239# a_7317_2550# 1.85e-20
C3477 x36.Q_N a_11628_2640# 0.572f
C3478 a_1061_4801# a_2147_5083# 0.00907f
C3479 x4.X a_1415_4801# 9.23e-21
C3480 a_1682_4775# a_1592_5167# 6.69e-20
C3481 a_3600_4086# a_4926_4296# 4.7e-22
C3482 a_3913_4112# a_4658_4086# 0.199f
C3483 a_3505_4086# x48.Q_N 0.178f
C3484 a_4155_4086# a_4454_4086# 0.0334f
C3485 x5.X a_11331_4086# 8.88e-19
C3486 a_3807_4801# x27.Q_N 5.03e-21
C3487 a_11195_4112# a_11565_4112# 4.11e-20
C3488 check[6] a_5991_2340# 1.42e-21
C3489 a_11630_4086# a_11543_3213# 1.61e-19
C3490 a_11629_4386# a_12030_3213# 3.78e-19
C3491 x39.Q_N a_10794_3239# 0.348f
C3492 a_12147_4801# a_11834_4086# 7.76e-20
C3493 x30.Q_N a_6759_3213# 0.00506f
C3494 a_6844_2640# x57.Q_N 4.82e-21
C3495 a_6845_2340# a_7317_2550# 0.15f
C3496 a_9638_3213# a_11543_3213# 3.71e-20
C3497 a_4854_3213# a_7072_3239# 1.86e-21
C3498 a_4367_3213# a_6198_3239# 3.42e-20
C3499 x33.Q_N a_9573_3239# 1.68e-19
C3500 x4.X a_4658_4086# 0.0102f
C3501 a_10983_4801# x36.Q_N 5.41e-22
C3502 a_1227_4801# a_929_3238# 1.49e-22
C3503 a_2853_5648# check[0] 0.164f
C3504 VDD a_9656_4394# 0.00984f
C3505 x4.X a_11565_4112# 8.15e-20
C3506 VDD a_2777_2366# 8.32e-19
C3507 a_2389_5648# x48.Q 0.00138f
C3508 VDD a_9551_5167# 0.00371f
C3509 VDD a_4789_3239# 1.15e-19
C3510 a_9238_4086# a_11089_4112# 5.07e-21
C3511 x42.Q_N a_9377_4112# 0.00167f
C3512 a_9710_4296# a_9578_4112# 0.0258f
C3513 a_9237_4386# a_11331_4086# 2.53e-20
C3514 x7.X a_1520_2366# 0.00311f
C3515 a_4019_4112# x77.Y 1.79e-19
C3516 x20.Q_N a_3504_2340# 6.66e-19
C3517 a_9442_4086# a_8402_3239# 2.9e-19
C3518 a_8697_4112# a_9638_3213# 9.49e-19
C3519 a_9238_4086# a_8857_3213# 5.04e-19
C3520 a_8939_4086# a_9151_3213# 2.12e-19
C3521 x33.Q_N x42.Q_N 0.00395f
C3522 a_11834_4086# a_11088_2366# 7.14e-22
C3523 a_11629_4386# a_11628_2640# 1.32e-20
C3524 a_11630_4086# a_11330_2340# 3.47e-21
C3525 sel_bit[0] x3.A 6.99e-21
C3526 check[5] a_9574_4801# 1.69e-20
C3527 a_10628_3239# D[2] 6.24e-20
C3528 D[4] a_9441_2340# 6.5e-20
C3529 D[1] a_12146_3239# 1.57e-20
C3530 x30.Q_N a_6546_2340# 0.16f
C3531 a_10794_3239# a_12737_3239# 6.86e-21
C3532 D[1] a_11761_3239# 5.48e-20
C3533 eob x20.Q_N 0.367f
C3534 x4.X a_1720_2648# 0.00102f
C3535 x27.D a_3600_4086# 0.00292f
C3536 check[0] a_3671_5674# 3.04e-19
C3537 x5.X a_1508_5167# 0.00288f
C3538 x20.Q_N x4.A 5.76e-19
C3539 x7.X a_4871_2648# 6.94e-19
C3540 check[2] a_11969_2366# 4.38e-19
C3541 a_6305_4112# a_6291_3605# 1.61e-19
C3542 a_6846_4086# a_5844_3239# 6.54e-20
C3543 a_6547_4086# a_6465_3213# 1.02e-19
C3544 a_5992_4086# a_6759_3213# 8.83e-19
C3545 a_6845_4386# a_6010_3239# 4.11e-20
C3546 x33.Q_N x7.X 0.263f
C3547 check[0] a_6846_4086# 2.15e-19
C3548 a_4926_4296# a_4453_2340# 6.08e-21
C3549 a_9237_4386# a_8696_2366# 1.93e-22
C3550 a_12031_4775# a_11834_4086# 4.44e-19
C3551 a_6606_4801# a_6978_4801# 3.34e-19
C3552 x27.Q_N a_4970_3239# 0.00341f
C3553 a_11544_4775# a_12102_4296# 2.85e-19
C3554 a_11076_5167# x39.Q_N 1e-19
C3555 a_1207_2340# a_1520_2366# 0.273f
C3556 a_10346_4801# a_10345_3239# 9.85e-20
C3557 a_9237_2340# a_11088_2366# 3.08e-19
C3558 a_9709_2550# a_9577_2366# 0.0258f
C3559 a_9236_2640# a_11330_2340# 4.16e-20
C3560 a_3452_3239# a_3983_3605# 0.0018f
C3561 a_3618_3239# a_3806_3239# 0.159f
C3562 a_4073_3213# a_4680_3239# 0.00187f
C3563 a_3899_3605# a_4854_3213# 4.7e-22
C3564 a_1682_4775# x27.D 2.67e-21
C3565 x4.X a_3170_4801# 9.94e-19
C3566 x5.X a_3913_4112# 1.32e-19
C3567 check[2] a_11970_4112# 3.49e-20
C3568 x48.Q a_3619_4801# 0.0352f
C3569 VDD x30.Q_N 0.444f
C3570 VDD a_3806_3239# 0.117f
C3571 a_6547_4086# a_5991_2340# 1.3e-22
C3572 a_6305_4112# a_6304_2366# 1.8e-19
C3573 x27.Q_N x57.Q_N 7.46e-20
C3574 D[6] a_2200_2366# 1.47e-19
C3575 a_2061_2340# a_4112_2648# 4.06e-20
C3576 check[5] a_8792_4801# 1.67e-19
C3577 a_11088_2366# a_12547_2366# 4.94e-21
C3578 x63.Q_N a_11288_2648# 2.02e-20
C3579 check[4] D[3] 0.00432f
C3580 a_11833_2340# a_11766_2732# 9.46e-19
C3581 a_11628_2640# a_12047_2648# 2.46e-19
C3582 a_10775_2340# a_11564_2366# 4.2e-20
C3583 check[1] x42.Q_N 0.0239f
C3584 x36.Q_N D[1] 1.36e-20
C3585 x5.X x4.X 0.0429f
C3586 x4.X a_6292_5167# 0.00132f
C3587 x4.X a_11856_3239# 0.00481f
C3588 a_7073_4801# a_7318_4296# 3.59e-20
C3589 x42.Q_N a_9954_4112# 2.4e-19
C3590 a_10156_4112# a_10776_4086# 8.26e-21
C3591 a_9237_4386# a_11195_4112# 1.71e-20
C3592 a_1976_4775# a_3807_4801# 2.23e-21
C3593 a_2463_4775# a_4681_4801# 1.86e-21
C3594 check[2] a_8237_4801# 5.48e-19
C3595 check[1] x7.X 0.134f
C3596 VDD a_3373_5674# 0.353f
C3597 a_3912_2366# a_4388_2366# 2.87e-21
C3598 x27.Q_N a_4680_3239# 0.0029f
C3599 a_6759_3213# a_7362_3239# 0.0552f
C3600 a_9873_5083# x33.Q_N 2.02e-20
C3601 VDD a_5992_4086# 0.716f
C3602 x4.X a_9237_4386# 0.048f
C3603 a_4855_4775# a_4454_4086# 0.00169f
C3604 a_4368_4775# a_4658_4086# 0.00268f
C3605 a_4681_4801# a_4453_4386# 1.96e-20
C3606 a_7050_4086# x42.Q_N 1.92e-20
C3607 x4.X a_11629_2340# 0.00254f
C3608 x20.Q_N x48.Q_N 0.00138f
C3609 x20.Q_N a_929_3238# 7.56e-20
C3610 a_6411_4112# a_6465_3213# 3.34e-20
C3611 check[6] a_5371_2366# 0.00326f
C3612 check[3] a_10776_4086# 1.93e-20
C3613 a_12031_4775# a_12548_4112# 4.23e-19
C3614 a_5991_2340# a_6504_2648# 0.00945f
C3615 a_9638_3213# a_10345_3239# 0.0968f
C3616 x33.Q_N a_8288_2340# 3.7e-19
C3617 a_9151_3213# D[1] 4.66e-19
C3618 D[7] x51.Q_N 0.00276f
C3619 x77.Y a_4585_3239# 0.00397f
C3620 a_7050_4086# x7.X 4.39e-21
C3621 VDD a_3504_2340# 0.205f
C3622 check[2] a_7247_4775# 2.07e-19
C3623 x5.X D[4] 3.43e-19
C3624 a_5845_4801# a_6466_4775# 0.117f
C3625 x20.Q_N a_2198_2732# 0.00203f
C3626 a_3505_4086# x77.Y 7.15e-21
C3627 VDD eob 2.6f
C3628 x39.Q_N a_12146_3239# 0.00968f
C3629 x39.Q_N a_11761_3239# 0.00399f
C3630 a_10794_3239# a_10982_3239# 0.163f
C3631 a_11075_3605# a_12030_3213# 4.7e-22
C3632 a_10628_3239# a_11159_3605# 0.0018f
C3633 a_11249_3213# a_11856_3239# 0.00187f
C3634 check[1] a_9173_4112# 1.03e-21
C3635 a_8997_3239# a_9573_3239# 2.46e-21
C3636 VDD x4.A 0.788f
C3637 check[2] a_9442_4086# 7.66e-19
C3638 sel_bit[0] a_1227_4801# 1.91e-20
C3639 VDD a_7362_3239# 4.88e-19
C3640 x27.D a_3900_5167# 8.53e-19
C3641 x7.X a_3912_2366# 0.00684f
C3642 check[2] a_12101_2550# 2.02e-19
C3643 x48.Q a_3452_3239# 8.21e-19
C3644 x45.Q_N x77.Y 1.27e-22
C3645 x42.Q_N a_8997_3239# 0.0309f
C3646 a_5845_4801# x75.Q 1.99e-20
C3647 x30.Q_N a_8696_2366# 8.85e-20
C3648 a_9237_2340# D[3] 0.336f
C3649 a_9709_2550# a_9953_2732# 0.00972f
C3650 a_9441_2340# a_10155_2366# 6.99e-20
C3651 a_10794_3239# a_11833_2340# 0.00154f
C3652 a_11543_3213# a_11330_2340# 2.17e-19
C3653 a_11249_3213# a_11629_2340# 0.00199f
C3654 a_12030_3213# a_11088_2366# 8.4e-19
C3655 VDD a_6781_4478# 0.00371f
C3656 check[1] a_8288_2340# 0.027f
C3657 x4.X a_9656_4394# 8.47e-19
C3658 a_8384_4086# a_8939_4086# 0.197f
C3659 a_7764_4112# x42.Q_N 5.48e-20
C3660 x5.X a_4368_4775# 4.59e-19
C3661 x4.X a_4789_3239# 1.05e-19
C3662 VDD D[2] 0.29f
C3663 VDD x60.Q_N 0.0716f
C3664 a_3453_4801# a_6199_4801# 3.65e-21
C3665 a_4681_4801# a_6011_4801# 3.02e-20
C3666 x5.X a_11544_4775# 0.00155f
C3667 x45.Q_N a_6930_3521# 0.00203f
C3668 a_2777_2732# a_2979_2366# 8.94e-19
C3669 a_8684_5167# a_9152_4775# 0.0633f
C3670 a_8237_4801# a_8591_4801# 0.0664f
C3671 a_8403_4801# a_9465_4801# 0.137f
C3672 a_5844_3239# a_6010_3239# 0.782f
C3673 check[0] a_6010_3239# 0.0252f
C3674 a_1520_2366# a_3599_2340# 8.34e-21
C3675 a_2060_2640# a_2200_2366# 0.00126f
C3676 a_1762_2340# a_2401_2366# 0.00316f
C3677 x36.Q_N x39.Q_N 0.00386f
C3678 check[4] a_9237_2340# 0.0399f
C3679 a_11088_2366# a_11628_2640# 0.139f
C3680 a_12031_4775# a_12030_3213# 0.00237f
C3681 a_10775_2340# a_11629_2340# 0.0492f
C3682 x77.Y a_4452_2640# 4.61e-20
C3683 a_11857_4801# a_11966_4801# 0.00707f
C3684 eob a_2265_2340# 9.03e-20
C3685 a_7764_4112# x7.X 4.77e-20
C3686 VDD a_1926_5083# 0.0117f
C3687 x48.Q a_4872_4394# 1.99e-19
C3688 check[6] x45.Q_N 6.19e-19
C3689 a_2853_5648# check[1] 0.0514f
C3690 x48.Q a_4586_4801# 3.31e-19
C3691 x7.X a_10680_2340# 7.8e-19
C3692 check[2] sel_bit[0] 0.0781f
C3693 a_4454_4086# a_4367_3213# 1.61e-19
C3694 a_4453_4386# a_4854_3213# 3.78e-19
C3695 clk_sar sel_bit[0] 0.343f
C3696 a_4453_2340# a_4112_2648# 1.25e-19
C3697 D[6] a_4388_2366# 1.34e-19
C3698 a_3912_2366# a_4018_2366# 0.0552f
C3699 a_4452_2640# a_4388_2732# 2.13e-19
C3700 a_4154_2340# a_4590_2732# 0.00412f
C3701 a_4970_3239# a_4925_2550# 1.01e-20
C3702 x36.Q_N a_12737_3239# 0.0107f
C3703 VDD x48.Q_N 0.0812f
C3704 sel_bit[1] a_1976_4775# 8.83e-20
C3705 VDD a_929_3238# 0.426f
C3706 VDD a_11970_4112# 0.0326f
C3707 check[2] a_10156_4112# 0.165f
C3708 x5.X a_8897_4394# 5.64e-19
C3709 x4.X x30.Q_N 0.426f
C3710 a_3619_4801# a_4318_5083# 2.46e-19
C3711 a_3453_4801# a_4539_5083# 0.00907f
C3712 x4.X a_3806_3239# 0.00861f
C3713 x20.Q_N a_2398_4801# 9.16e-20
C3714 x5.X a_7363_4801# 2.04e-19
C3715 a_11630_4086# a_12102_4296# 0.15f
C3716 a_11629_4386# x39.Q_N 0.00118f
C3717 a_2853_5648# a_3877_5674# 8.24e-20
C3718 check[1] a_3671_5674# 5.38e-19
C3719 check[6] a_4452_2640# 0.0327f
C3720 a_6760_4775# a_7246_3213# 1.06e-20
C3721 a_7247_4775# a_8591_4801# 8.26e-21
C3722 a_7247_4775# a_6759_3213# 1.08e-22
C3723 x39.Q_N a_9151_3213# 3.3e-20
C3724 check[1] a_6846_4086# 0.441f
C3725 a_5896_2340# a_6304_2366# 6.04e-19
C3726 a_4592_2366# a_4793_2366# 3.34e-19
C3727 a_8402_3239# a_9101_3521# 2.46e-19
C3728 a_8236_3239# a_9322_3521# 0.00907f
C3729 x36.Q_N a_11768_2366# 0.00473f
C3730 a_10629_4801# a_11715_5083# 0.00907f
C3731 a_10795_4801# a_11494_5083# 2.46e-19
C3732 a_4926_4296# a_5372_4112# 0.0367f
C3733 a_4453_4386# a_4593_4112# 0.00126f
C3734 a_4155_4086# a_4794_4112# 0.00316f
C3735 VDD a_2198_2732# 0.0198f
C3736 a_8939_4086# a_9173_4478# 0.00976f
C3737 a_8384_4086# a_8803_4112# 0.0397f
C3738 check[2] check[6] 7.32e-20
C3739 a_8697_4112# a_9375_4478# 0.00652f
C3740 VDD a_8237_4801# 0.81f
C3741 x27.Q_N a_4926_4296# 5.7e-19
C3742 x5.X a_6845_2340# 2.59e-20
C3743 a_9465_4801# a_9710_4296# 3.59e-20
C3744 sel_bit[0] a_4074_4775# 0.00112f
C3745 a_4074_4775# x77.Y 5.16e-21
C3746 a_3373_5674# x4.X 5.96e-20
C3747 sel_bit[0] x20.Q_N 2.7e-20
C3748 x20.Q_N x77.Y 0.0156f
C3749 D[1] a_11075_3605# 2.08e-19
C3750 a_10345_3239# a_11543_3213# 5.62e-20
C3751 eob a_1508_5167# 0.0514f
C3752 a_9151_3213# a_9709_2550# 1.62e-19
C3753 a_4213_3239# a_3599_2340# 4.6e-20
C3754 check[3] a_10628_3239# 1.99e-20
C3755 a_4680_3239# a_4925_2550# 1.85e-20
C3756 a_9638_3213# a_9441_2340# 2.52e-19
C3757 x4.X a_5992_4086# 0.1f
C3758 a_6845_4386# a_7318_4296# 0.155f
C3759 a_6547_4086# x45.Q_N 0.0285f
C3760 a_6846_4086# a_7050_4086# 0.117f
C3761 a_1508_5167# x4.A 0.00373f
C3762 x7.X D[6] 0.00566f
C3763 check[0] a_4591_4478# 1.2e-20
C3764 x7.X a_6465_3213# 4.84e-19
C3765 x5.X a_6606_4801# 9.34e-19
C3766 a_6760_4775# a_7159_5167# 0.00133f
C3767 a_5845_4801# a_7481_5083# 1.25e-19
C3768 a_6011_4801# a_6978_4801# 0.00126f
C3769 a_6292_5167# a_6606_4801# 0.0258f
C3770 x30.Q_N D[4] 0.005f
C3771 a_1338_5674# a_2853_5648# 1e-19
C3772 D[1] a_11088_2366# 3.91e-20
C3773 a_11856_3239# a_11965_3239# 0.00707f
C3774 a_9873_5083# a_10629_4801# 4.06e-20
C3775 a_9236_2640# a_9441_2340# 0.153f
C3776 a_8696_2366# x60.Q_N 0.00553f
C3777 a_12030_3213# x66.Q_N 0.124f
C3778 x4.X a_3504_2340# 0.0105f
C3779 VDD a_7247_4775# 0.72f
C3780 VDD a_11159_3605# 0.0042f
C3781 a_4074_4775# check[6] 4.81e-21
C3782 x7.X a_5991_2340# 0.00445f
C3783 a_4794_4112# a_4925_2550# 1.72e-22
C3784 a_11629_4386# a_11769_4112# 0.00126f
C3785 x5.X a_10346_4801# 0.0293f
C3786 a_11331_4086# a_11970_4112# 0.00316f
C3787 a_11834_4086# a_12548_4112# 6.99e-20
C3788 a_12102_4296# a_12346_4478# 0.00972f
C3789 eob x4.X 0.224f
C3790 check[5] a_8858_4775# 6.94e-19
C3791 a_2265_2340# a_2198_2732# 9.46e-19
C3792 a_2060_2640# a_2479_2648# 2.46e-19
C3793 x51.Q_N a_1720_2648# 2.02e-20
C3794 a_1207_2340# D[6] 3.57e-20
C3795 a_1520_2366# a_2979_2366# 6.59e-21
C3796 a_10155_2366# a_11629_2340# 3.65e-21
C3797 D[3] a_11628_2640# 4.01e-20
C3798 check[2] a_2788_5674# 0.00675f
C3799 a_12146_3239# a_11833_2340# 3.49e-20
C3800 a_4367_3213# x75.Q 3.3e-19
C3801 a_4854_3213# a_5561_3239# 0.0968f
C3802 a_11250_4775# check[3] 0.00109f
C3803 x4.X x4.A 0.00766f
C3804 a_4453_4386# a_5170_4112# 0.0019f
C3805 x5.X a_5897_4086# 0.0764f
C3806 VDD a_9442_4086# 0.487f
C3807 x48.Q a_3600_4086# 0.00969f
C3808 x4.X a_7362_3239# 5.65e-19
C3809 x7.X a_9374_2732# 9.52e-19
C3810 VDD a_12101_2550# 0.172f
C3811 x27.Q_N a_6760_4775# 6.16e-21
C3812 comparator_out a_653_3238# 0.196f
C3813 a_4681_4801# a_4854_3213# 4.82e-21
C3814 D[6] a_4018_2366# 0.0021f
C3815 a_4855_4775# a_4680_3239# 1.33e-23
C3816 a_8684_5167# a_8236_3239# 8.3e-21
C3817 a_5844_3239# a_8236_3239# 0.00176f
C3818 a_8403_4801# a_8857_3213# 3.18e-21
C3819 a_3599_2340# a_3912_2366# 0.273f
C3820 a_8591_4801# a_8792_4801# 3.67e-19
C3821 a_9465_4801# a_9370_4801# 0.00276f
C3822 a_5844_3239# a_6977_3239# 2.56e-19
C3823 a_6759_3213# a_6930_3521# 0.00652f
C3824 a_9152_4775# x33.Q_N 0.0059f
C3825 a_9639_4775# a_9873_5083# 0.00945f
C3826 a_6010_3239# a_6399_3239# 0.0019f
C3827 a_2853_5648# a_3453_4801# 7.76e-20
C3828 a_6465_3213# a_6605_3239# 0.07f
C3829 x4.X a_6781_4478# 2.12e-19
C3830 x48.Q a_1682_4775# 4.88e-21
C3831 a_6547_4086# a_6781_4112# 0.00707f
C3832 a_6845_4386# a_8289_4086# 4.36e-19
C3833 a_7050_4086# a_7562_4478# 6.69e-20
C3834 a_6305_4112# a_6985_4112# 3.73e-19
C3835 x45.Q_N a_6411_4112# 0.0455f
C3836 VDD a_2398_4801# 6.04e-19
C3837 a_6846_4086# a_7764_4112# 0.0664f
C3838 a_1822_4801# a_1511_4112# 1.33e-19
C3839 x4.X D[2] 4e-19
C3840 x4.X x60.Q_N 0.00784f
C3841 VDD a_9574_4801# 7.87e-19
C3842 check[5] a_7561_2366# 5.2e-20
C3843 check[6] a_6759_3213# 8.24e-21
C3844 D[5] a_5896_2340# 0.0999f
C3845 check[0] a_6984_2366# 3.17e-19
C3846 D[0] a_8590_3239# 5.04e-19
C3847 a_6605_3239# a_5991_2340# 4.6e-20
C3848 check[4] a_10983_4801# 0.164f
C3849 eob x7.A 0.0353f
C3850 x77.Y a_3618_3239# 0.528f
C3851 x36.Q_N a_11833_2340# 0.179f
C3852 a_1682_4775# a_2147_5083# 9.46e-19
C3853 a_1227_4801# a_2375_5167# 2.13e-19
C3854 a_1061_4801# a_1822_4801# 6.04e-20
C3855 a_3913_4112# x48.Q_N 0.00553f
C3856 a_4453_4386# a_4658_4086# 0.153f
C3857 a_4855_4775# a_4794_4112# 1.79e-20
C3858 x5.X a_11630_4086# 0.26f
C3859 VDD sel_bit[0] 1.26f
C3860 VDD x77.Y 0.423f
C3861 a_621_4112# a_1511_4112# 2.76e-19
C3862 check[5] x42.Q_N 6.88e-19
C3863 a_11834_4086# a_12030_3213# 2.47e-19
C3864 x39.Q_N a_11075_3605# 0.152f
C3865 a_12102_4296# a_11543_3213# 1.71e-19
C3866 x30.Q_N a_7072_3239# 0.00298f
C3867 x30.Q_N a_7363_4801# 0.00129f
C3868 a_9151_3213# a_10982_3239# 3.42e-20
C3869 a_9638_3213# a_11856_3239# 1.86e-21
C3870 a_4367_3213# a_4970_3239# 0.0552f
C3871 x4.X x48.Q_N 0.00819f
C3872 x4.X a_929_3238# 0.00384f
C3873 VDD a_10156_4112# 0.109f
C3874 x4.X a_11970_4112# 0.00309f
C3875 VDD a_4388_2732# 0.00402f
C3876 check[5] x7.X 0.0221f
C3877 x7.X a_2060_2640# 0.113f
C3878 a_9237_4386# a_11630_4086# 2.9e-21
C3879 VDD a_6930_3521# 0.0163f
C3880 a_2463_4775# a_3170_4801# 0.0968f
C3881 x42.Q_N a_10776_4086# 7.84e-21
C3882 a_1976_4775# x27.D 0.00388f
C3883 a_9238_4086# a_9151_3213# 1.61e-19
C3884 check[6] a_6931_5083# 1.5e-21
C3885 x42.Q_N a_8402_3239# 0.345f
C3886 a_9237_4386# a_9638_3213# 3.78e-19
C3887 x20.Q_N a_2200_2366# 0.00397f
C3888 x39.Q_N a_11088_2366# 6.35e-20
C3889 a_11629_4386# a_11833_2340# 1.26e-21
C3890 a_897_4112# D[7] 1.81e-20
C3891 a_11630_4086# a_11629_2340# 1.55e-19
C3892 check[6] a_3618_3239# 7.95e-22
C3893 D[1] D[3] 0.345f
C3894 x30.Q_N a_6845_2340# 0.0463f
C3895 a_11249_3213# D[2] 1.23e-20
C3896 D[4] x60.Q_N 0.00109f
C3897 a_7562_4478# a_7764_4112# 8.94e-19
C3898 x4.X a_2198_2732# 9.81e-19
C3899 VDD check[6] 0.503f
C3900 a_6411_4112# a_6781_4112# 4.11e-20
C3901 a_10776_4086# x7.X 0.00196f
C3902 x4.X a_8237_4801# 0.0043f
C3903 x5.X a_2463_4775# 0.016f
C3904 x7.X a_5371_2366# 0.155f
C3905 x7.X a_8402_3239# 0.147f
C3906 VDD check[3] 0.745f
C3907 a_6305_4112# a_7246_3213# 9.49e-19
C3908 a_6547_4086# a_6759_3213# 2.12e-19
C3909 a_6846_4086# a_6465_3213# 5.04e-19
C3910 a_7050_4086# a_6010_3239# 2.9e-19
C3911 check[0] a_7318_4296# 4.24e-20
C3912 a_9237_4386# a_9236_2640# 1.32e-20
C3913 a_9238_4086# a_8938_2340# 3.47e-21
C3914 a_9442_4086# a_8696_2366# 7.14e-22
C3915 a_1207_2340# a_2060_2640# 0.0264f
C3916 a_1520_2366# a_1762_2340# 0.124f
C3917 a_11857_4801# a_12102_4296# 3.59e-20
C3918 a_6606_4801# x30.Q_N 1.33e-19
C3919 a_12030_3213# a_12547_2366# 2.38e-19
C3920 check[4] D[1] 0.435f
C3921 a_9237_2340# a_11628_2640# 4e-20
C3922 a_9236_2640# a_11629_2340# 2.9e-21
C3923 a_9709_2550# a_11088_2366# 5.19e-21
C3924 a_9755_4801# a_9151_3213# 1.05e-20
C3925 a_4367_3213# a_4680_3239# 0.124f
C3926 a_4073_3213# a_3983_3605# 6.69e-20
C3927 a_3618_3239# a_4317_3521# 2.46e-19
C3928 a_3899_3605# a_3806_3239# 0.0367f
C3929 a_3452_3239# a_4538_3521# 0.00907f
C3930 x33.Q_N a_11390_4801# 6.84e-20
C3931 x5.X a_4453_4386# 0.009f
C3932 x48.Q a_3900_5167# 0.00702f
C3933 x7.A a_929_3238# 0.3f
C3934 a_653_3238# x7.X 0.00275f
C3935 a_6845_4386# a_6304_2366# 1.93e-22
C3936 VDD a_4317_3521# 0.0107f
C3937 a_5089_5083# check[6] 5.84e-21
C3938 x27.Q_N a_5562_4801# 0.182f
C3939 a_2060_2640# a_4018_2366# 2.19e-20
C3940 a_12548_4112# a_12030_3213# 2.07e-19
C3941 D[6] a_3599_2340# 0.0144f
C3942 a_2979_2366# a_3912_2366# 3.42e-20
C3943 a_11330_2340# a_11564_2366# 0.00707f
C3944 a_12031_4775# a_12737_3239# 4.94e-20
C3945 a_11629_2340# a_12345_2732# 0.0018f
C3946 a_11628_2640# a_12547_2366# 0.159f
C3947 a_11088_2366# a_11768_2366# 3.73e-19
C3948 a_11833_2340# a_12047_2648# 0.0104f
C3949 x36.Q_N a_12738_4801# 0.184f
C3950 a_12265_5083# check[3] 0.0011f
C3951 x4.X a_7247_4775# 0.103f
C3952 x4.X a_11159_3605# 9.07e-19
C3953 x7.X a_11564_2732# 1.8e-19
C3954 a_9377_4112# a_9578_4112# 3.34e-19
C3955 a_6606_4801# a_5992_4086# 1.08e-19
C3956 check[2] a_8858_4775# 5.69e-19
C3957 a_1976_4775# a_2579_4801# 0.0551f
C3958 a_10681_4086# a_11089_4112# 4.37e-19
C3959 a_3912_2366# a_4793_2366# 0.00943f
C3960 a_4154_2340# a_4592_2366# 0.00276f
C3961 a_4453_2340# a_5896_2340# 8.18e-19
C3962 VDD a_2788_5674# 6.52e-19
C3963 a_7072_3239# a_7362_3239# 0.0282f
C3964 x33.Q_N a_8236_3239# 2.78e-19
C3965 a_7246_3213# a_7181_3239# 4.2e-20
C3966 a_8998_4801# a_9151_3213# 1.61e-20
C3967 VDD a_6547_4086# 0.34f
C3968 a_3505_4086# x7.X 2.05e-21
C3969 x4.X a_9442_4086# 0.00986f
C3970 a_4681_4801# a_4658_4086# 2.59e-19
C3971 a_4855_4775# a_4926_4296# 2.97e-21
C3972 x4.X a_12101_2550# 0.00146f
C3973 x5.X D[0] 0.00133f
C3974 sel_bit[0] a_1508_5167# 3.52e-20
C3975 a_6304_2366# a_6780_2732# 0.00133f
C3976 check[3] a_11331_4086# 4.58e-20
C3977 a_2883_5674# a_3258_5648# 0.014f
C3978 a_9464_3239# D[1] 5.18e-20
C3979 a_2883_5674# sel_bit[1] 0.0353f
C3980 a_1227_4801# x7.X 2.05e-22
C3981 check[1] a_7954_4801# 0.0169f
C3982 a_5897_4086# a_5992_4086# 0.0968f
C3983 x77.Y x75.Q_N 3.94e-19
C3984 a_4389_4112# a_4794_4112# 2.46e-21
C3985 x45.Q_N x7.X 0.00129f
C3986 x4.X a_2398_4801# 0.00124f
C3987 VDD a_2200_2366# 0.00214f
C3988 x5.X a_6011_4801# 0.0199f
C3989 x4.X a_9574_4801# 2.39e-19
C3990 a_1511_4112# a_1520_2366# 7.01e-19
C3991 a_6011_4801# a_6292_5167# 0.155f
C3992 a_5845_4801# a_6760_4775# 0.125f
C3993 sel_bit[0] a_3913_4112# 5.05e-19
C3994 x20.Q_N a_2479_2648# 0.00136f
C3995 a_3913_4112# x77.Y 3.94e-20
C3996 check[0] a_3619_4801# 0.00149f
C3997 x5.X a_11966_4801# 5.38e-20
C3998 x39.Q_N x66.Q_N 3.91e-19
C3999 D[1] a_9237_2340# 0.0263f
C4000 a_9152_4775# a_10629_4801# 1.67e-19
C4001 a_11075_3605# a_10982_3239# 0.0367f
C4002 a_6845_2340# x60.Q_N 2.94e-19
C4003 a_11543_3213# a_11856_3239# 0.124f
C4004 a_11249_3213# a_11159_3605# 6.69e-20
C4005 a_10794_3239# a_9754_3239# 9.75e-21
C4006 check[1] a_9578_4112# 3.76e-20
C4007 check[1] a_8236_3239# 0.0444f
C4008 check[2] x42.Q_N 8.18e-19
C4009 VDD a_6504_2648# 0.00506f
C4010 x5.X a_8697_4112# 0.00599f
C4011 sel_bit[0] x4.X 4e-20
C4012 check[5] a_6846_4086# 0.0346f
C4013 VDD a_9101_3521# 0.00984f
C4014 x4.X x77.Y 0.07f
C4015 a_7247_4775# a_7186_4112# 1.79e-20
C4016 x7.X a_4452_2640# 0.109f
C4017 x27.D a_4855_4775# 4.69e-21
C4018 x5.X a_5561_3239# 0.00125f
C4019 x42.Q_N a_10628_3239# 1.47e-19
C4020 check[4] x39.Q_N 6.54e-19
C4021 x42.Q_N a_9369_3239# 0.00401f
C4022 x30.Q_N a_9236_2640# 1.21e-20
C4023 check[6] x75.Q_N 0.00302f
C4024 D[2] a_11965_3239# 9.32e-21
C4025 a_12030_3213# a_11628_2640# 3.43e-19
C4026 check[3] a_11194_2366# 1.29e-19
C4027 a_11543_3213# a_11629_2340# 2.19e-19
C4028 x66.Q_N a_12737_3239# 0.178f
C4029 VDD a_6411_4112# 0.00996f
C4030 x4.X a_10156_4112# 0.00621f
C4031 check[2] x7.X 0.125f
C4032 x4.X a_4388_2732# 4.32e-19
C4033 x5.X a_4681_4801# 1.74e-19
C4034 a_8384_4086# a_9238_4086# 0.0492f
C4035 check[6] a_3913_4112# 7.75e-22
C4036 a_8697_4112# a_9237_4386# 0.139f
C4037 x4.X a_6930_3521# 9.99e-19
C4038 x4.X a_8792_4801# 8.46e-20
C4039 a_1062_5674# a_897_4112# 9.53e-20
C4040 x7.X a_7561_2732# 8.23e-19
C4041 x7.X a_10628_3239# 0.148f
C4042 x45.Q_N a_6605_3239# 0.031f
C4043 x27.Q_N a_5169_2366# 0.00224f
C4044 x5.X a_11857_4801# 0.00141f
C4045 a_2979_2366# D[6] 6.09e-19
C4046 a_6010_3239# a_6465_3213# 0.153f
C4047 a_2060_2640# a_3599_2340# 3.6e-19
C4048 a_2061_2340# a_2401_2366# 6.04e-20
C4049 D[3] a_11768_2366# 7.83e-20
C4050 a_8858_4775# a_8591_4801# 6.99e-20
C4051 a_8403_4801# a_8768_5167# 4.45e-20
C4052 a_9152_4775# a_9639_4775# 0.273f
C4053 a_5844_3239# a_6291_3605# 0.15f
C4054 a_2265_2340# a_2200_2366# 9.75e-19
C4055 check[0] a_6291_3605# 7.4e-20
C4056 check[4] a_9709_2550# 0.00101f
C4057 a_11330_2340# a_11629_2340# 0.0334f
C4058 a_11088_2366# a_11833_2340# 0.199f
C4059 a_10775_2340# a_12101_2550# 4.7e-22
C4060 x77.Y a_4657_2340# 1.11e-19
C4061 x4.X check[6] 0.0328f
C4062 VDD a_2375_5167# 0.00488f
C4063 x4.X check[3] 0.316f
C4064 a_4926_4296# a_4367_3213# 1.71e-19
C4065 a_4658_4086# a_4854_3213# 2.47e-19
C4066 a_4453_2340# a_4590_2732# 0.00907f
C4067 D[6] a_4793_2366# 4.25e-19
C4068 check[1] a_1511_4112# 5.91e-22
C4069 a_5844_3239# a_6304_2366# 1.89e-19
C4070 a_6010_3239# a_5991_2340# 3.73e-19
C4071 check[0] a_6304_2366# 0.00297f
C4072 sel_bit[1] a_2289_4801# 1.47e-20
C4073 x20.Q_N a_4113_4394# 6.16e-20
C4074 VDD comparator_out 0.186f
C4075 x5.X a_9375_4478# 7.3e-19
C4076 check[2] a_9173_4112# 1.17e-20
C4077 x20.Q_N x7.X 0.0882f
C4078 a_3619_4801# a_4767_5167# 2.13e-19
C4079 a_3453_4801# a_4214_4801# 6.04e-20
C4080 x4.X a_4317_3521# 0.00111f
C4081 a_4074_4775# a_4539_5083# 9.46e-19
C4082 x5.X a_9102_5083# 3.46e-19
C4083 check[2] a_9873_5083# 4.31e-19
C4084 a_11834_4086# x39.Q_N 0.00118f
C4085 check[6] a_4657_2340# 6.83e-20
C4086 a_7247_4775# a_7072_3239# 1.33e-23
C4087 a_7247_4775# a_7363_4801# 0.0397f
C4088 a_7073_4801# a_7246_3213# 4.82e-21
C4089 a_6760_4775# a_7182_4801# 2.87e-21
C4090 a_5896_2340# a_6844_2640# 8.38e-21
C4091 a_3452_3239# a_5844_3239# 0.00176f
C4092 check[1] a_7318_4296# 0.0013f
C4093 a_8236_3239# a_8997_3239# 6.04e-20
C4094 a_8857_3213# a_9322_3521# 9.46e-19
C4095 a_8402_3239# a_9550_3605# 2.13e-19
C4096 check[0] a_3452_3239# 2.98e-21
C4097 a_11250_4775# a_11715_5083# 9.46e-19
C4098 a_10795_4801# a_11943_5167# 2.13e-19
C4099 x36.Q_N a_12345_2366# 0.00224f
C4100 a_10629_4801# a_11390_4801# 6.04e-20
C4101 x33.Q_N a_8791_3239# 6.75e-20
C4102 a_4454_4086# a_4794_4112# 6.04e-20
C4103 a_4453_4386# a_5992_4086# 1.24e-19
C4104 a_4658_4086# a_4593_4112# 9.75e-19
C4105 VDD a_2479_2648# 0.0122f
C4106 VDD a_8858_4775# 0.488f
C4107 a_8939_4086# a_8803_4112# 0.0282f
C4108 a_9237_4386# a_9375_4478# 1.09e-19
C4109 a_8697_4112# a_9656_4394# 1.21e-20
C4110 x5.X a_897_4112# 0.00452f
C4111 a_5562_4801# a_5845_4801# 8.18e-19
C4112 x5.X a_10345_3239# 0.00125f
C4113 a_8998_4801# a_8384_4086# 1.08e-19
C4114 x42.Q_N a_6759_3213# 3.3e-20
C4115 a_11630_4086# D[2] 3.53e-19
C4116 x20.Q_N a_1207_2340# 0.144f
C4117 a_8237_4801# a_10346_4801# 1.03e-19
C4118 x30.Q_N D[0] 3.29e-19
C4119 D[1] a_12030_3213# 1.69e-20
C4120 x33.Q_N a_9172_2366# 9.42e-19
C4121 a_9464_3239# a_9709_2550# 1.85e-20
C4122 eob a_2463_4775# 0.00567f
C4123 x4.X a_6547_4086# 0.00727f
C4124 a_7050_4086# a_7318_4296# 0.205f
C4125 a_6846_4086# x45.Q_N 0.00113f
C4126 VDD a_4388_2366# 1.64e-19
C4127 x7.X a_6759_3213# 7.49e-19
C4128 a_8591_4801# x7.X 1.94e-20
C4129 a_3505_4086# a_3599_2340# 1.57e-20
C4130 check[0] a_4872_4394# 8.58e-21
C4131 x5.X a_6978_4801# 2.58e-19
C4132 a_929_3238# x51.Q_N 1.42e-19
C4133 x20.Q_N a_4018_2366# 1.31e-20
C4134 a_7073_4801# a_7159_5167# 0.00976f
C4135 a_4971_4801# a_4790_4801# 4.11e-20
C4136 a_6011_4801# x30.Q_N 1.04e-19
C4137 a_2389_5648# check[1] 0.0168f
C4138 check[2] a_2853_5648# 0.112f
C4139 a_9236_2640# x60.Q_N 5.14e-21
C4140 a_9237_2340# a_9709_2550# 0.15f
C4141 check[3] a_10775_2340# 2.56e-20
C4142 x33.Q_N a_10795_4801# 2.19e-19
C4143 a_1338_5674# a_1511_4112# 4.25e-21
C4144 VDD a_6199_4801# 0.109f
C4145 x48.Q a_1976_4775# 4.67e-19
C4146 a_4855_4775# a_5562_4801# 0.0968f
C4147 x7.X a_6546_2340# 0.00104f
C4148 a_4368_4775# check[6] 0.00421f
C4149 x39.Q_N a_12548_4112# 8.27e-20
C4150 a_11629_4386# a_12346_4112# 0.0019f
C4151 a_9238_4086# D[3] 1.26e-20
C4152 a_11630_4086# a_11970_4112# 6.04e-20
C4153 a_11834_4086# a_11769_4112# 9.75e-19
C4154 x27.Q_N a_5896_2340# 1.79e-19
C4155 a_2265_2340# a_2479_2648# 0.0104f
C4156 check[5] a_9152_4775# 0.00306f
C4157 a_1762_2340# D[6] 2.05e-19
C4158 check[5] a_6010_3239# 2.24e-21
C4159 a_2060_2640# a_2979_2366# 0.163f
C4160 a_2061_2340# a_2777_2732# 0.0018f
C4161 check[1] a_8289_4086# 0.125f
C4162 D[3] a_11833_2340# 6.82e-20
C4163 check[2] a_3671_5674# 0.00323f
C4164 a_1338_5674# a_1061_4801# 0.0022f
C4165 a_11544_4775# check[3] 0.00913f
C4166 a_12031_4775# a_12738_4801# 0.0968f
C4167 check[1] a_9172_2366# 1.35e-19
C4168 VDD x42.Q_N 0.457f
C4169 check[2] a_6846_4086# 2.36e-20
C4170 x4.X a_6504_2648# 0.00102f
C4171 x48.Q a_4155_4086# 0.00101f
C4172 a_5845_4801# a_6305_4112# 3.05e-19
C4173 a_6011_4801# a_5992_4086# 6.63e-19
C4174 x7.X a_9655_2648# 7e-19
C4175 x4.X a_9101_3521# 2.91e-19
C4176 a_1976_4775# a_2147_5083# 0.00652f
C4177 sel_bit[1] reset 1.45e-20
C4178 x7.X a_3618_3239# 4.91e-19
C4179 a_9639_4775# a_9578_4112# 1.79e-20
C4180 a_4214_4801# a_4790_4801# 2.46e-21
C4181 x27.Q_N a_7073_4801# 7.65e-21
C4182 check[4] a_9238_4086# 0.0367f
C4183 a_5844_3239# D[5] 5.19e-19
C4184 a_3504_2340# x54.Q_N 0.178f
C4185 a_8684_5167# a_8857_3213# 3.52e-21
C4186 a_3599_2340# a_4452_2640# 0.0264f
C4187 check[0] D[5] 0.228f
C4188 a_8858_4775# a_8683_3605# 1.33e-23
C4189 a_8403_4801# a_9151_3213# 2.05e-21
C4190 a_3912_2366# a_4154_2340# 0.124f
C4191 a_7072_3239# a_6930_3521# 0.00412f
C4192 check[1] a_3619_4801# 7.46e-20
C4193 a_6465_3213# a_6977_3239# 9.75e-19
C4194 a_6291_3605# a_6399_3239# 0.00812f
C4195 a_5844_3239# x72.Q_N 1.07e-19
C4196 a_2853_5648# a_4074_4775# 1.12e-19
C4197 a_6759_3213# a_6605_3239# 0.00943f
C4198 a_9465_4801# x33.Q_N 8.55e-20
C4199 a_7246_3213# a_7158_3605# 7.71e-20
C4200 VDD a_4113_4394# 0.00555f
C4201 x4.X a_6411_4112# 0.00336f
C4202 a_2853_5648# x20.Q_N 2.38e-20
C4203 VDD x7.X 1.93f
C4204 VDD a_4539_5083# 0.0172f
C4205 a_7318_4296# a_7764_4112# 0.0367f
C4206 a_6547_4086# a_7186_4112# 0.00316f
C4207 a_6845_4386# a_6985_4112# 0.00126f
C4208 VDD a_11715_5083# 0.0163f
C4209 check[6] a_7363_4801# 1.16e-20
C4210 a_4925_2550# a_5169_2366# 0.00812f
C4211 D[0] a_7362_3239# 8.51e-20
C4212 check[4] a_9755_4801# 2.75e-19
C4213 x77.Y a_3899_3605# 0.181f
C4214 x36.Q_N x63.Q_N 4.08e-19
C4215 a_1061_4801# a_3453_4801# 0.00176f
C4216 a_1338_5674# a_2389_5648# 0.00448f
C4217 a_1682_4775# a_1822_4801# 0.07f
C4218 a_1061_4801# a_2194_4801# 2.56e-19
C4219 a_1227_4801# a_1616_4801# 0.0019f
C4220 a_4453_4386# x48.Q_N 4.82e-21
C4221 a_4454_4086# a_4926_4296# 0.15f
C4222 VDD a_1207_2340# 0.607f
C4223 x5.X a_12102_4296# 1.62e-19
C4224 check[6] a_6845_2340# 3.11e-22
C4225 x39.Q_N a_12030_3213# 0.144f
C4226 a_12102_4296# a_11856_3239# 2.37e-20
C4227 a_6304_2366# a_6780_2366# 2.87e-21
C4228 x33.Q_N a_8802_2366# 0.0102f
C4229 a_9151_3213# a_9754_3239# 0.0552f
C4230 a_5088_3521# a_5844_3239# 4.06e-20
C4231 a_4680_3239# a_4970_3239# 0.0282f
C4232 a_4854_3213# a_4789_3239# 4.2e-20
C4233 VDD a_9173_4112# 3.55e-19
C4234 x4.X comparator_out 1.47e-19
C4235 VDD a_4018_2366# 0.0028f
C4236 sel_bit[0] a_2784_5996# 0.00164f
C4237 x7.X a_2265_2340# 0.00311f
C4238 VDD a_9873_5083# 0.00506f
C4239 a_8939_4086# x39.Q_N 1.36e-20
C4240 a_2289_4801# x27.D 1.17e-20
C4241 VDD a_6605_3239# 5.47e-21
C4242 check[0] a_3600_4086# 9e-20
C4243 a_9710_4296# a_9151_3213# 1.71e-19
C4244 a_9442_4086# a_9638_3213# 2.47e-19
C4245 x42.Q_N a_8683_3605# 0.152f
C4246 check[6] a_6606_4801# 1.78e-19
C4247 x20.Q_N a_3599_2340# 3.36e-19
C4248 x39.Q_N a_11628_2640# 4.61e-20
C4249 a_8383_2340# a_8896_2648# 0.00945f
C4250 a_12102_4296# a_11629_2340# 6.08e-21
C4251 a_11543_3213# D[2] 3.13e-19
C4252 a_12030_3213# a_12737_3239# 0.0968f
C4253 x30.Q_N a_7317_2550# 0.181f
C4254 a_8998_4801# check[4] 1.23e-20
C4255 check[1] a_6304_2366# 1.25e-21
C4256 a_6845_4386# a_7562_4112# 0.0019f
C4257 x4.X a_2479_2648# 2.86e-19
C4258 x4.X a_8858_4775# 9.41e-19
C4259 x5.X a_1415_4801# 0.00367f
C4260 VDD a_8288_2340# 0.189f
C4261 x7.X a_8683_3605# 0.0011f
C4262 a_6845_4386# a_7246_3213# 3.78e-19
C4263 x45.Q_N a_6010_3239# 0.346f
C4264 a_6846_4086# a_6759_3213# 1.61e-19
C4265 a_9237_4386# a_9441_2340# 1.26e-21
C4266 x42.Q_N a_8696_2366# 6.41e-20
C4267 a_9238_4086# a_9237_2340# 1.55e-19
C4268 a_7954_4801# check[5] 0.129f
C4269 a_1762_2340# a_2060_2640# 0.137f
C4270 a_6978_4801# x30.Q_N 1.41e-19
C4271 a_11390_4801# a_10776_4086# 1.08e-19
C4272 a_1520_2366# a_2061_2340# 0.125f
C4273 D[2] a_11330_2340# 2.3e-20
C4274 a_4073_3213# a_4538_3521# 9.46e-19
C4275 a_3618_3239# a_4766_3605# 2.13e-19
C4276 a_3452_3239# a_4213_3239# 6.04e-20
C4277 x33.Q_N a_11762_4801# 3.57e-20
C4278 check[1] a_6710_5083# 1.55e-19
C4279 check[1] a_8802_2366# 0.00244f
C4280 a_1062_5674# x5.X 0.00571f
C4281 x5.X a_4658_4086# 4.53e-19
C4282 check[6] a_5897_4086# 0.00265f
C4283 x48.Q a_4855_4775# 0.00105f
C4284 x7.X a_8696_2366# 0.00714f
C4285 VDD a_4766_3605# 0.00394f
C4286 a_6846_4086# a_6546_2340# 3.47e-21
C4287 a_7050_4086# a_6304_2366# 7.14e-22
C4288 a_6845_4386# a_6844_2640# 1.32e-20
C4289 comparator_out x7.A 0.0101f
C4290 VDD a_2853_5648# 0.413f
C4291 check[5] a_8236_3239# 0.00639f
C4292 D[6] a_4154_2340# 8.45e-19
C4293 a_8237_4801# D[0] 1.99e-20
C4294 check[0] a_4453_2340# 0.00712f
C4295 a_12101_2550# a_12345_2732# 0.00972f
C4296 a_11833_2340# a_12547_2366# 6.99e-20
C4297 a_11330_2340# a_11969_2366# 0.00316f
C4298 a_11628_2640# a_11768_2366# 0.00126f
C4299 x4.X a_6199_4801# 2.3e-19
C4300 a_3453_4801# a_3619_4801# 0.75f
C4301 x4.X a_9573_3239# 1.05e-19
C4302 a_10156_4112# a_11630_4086# 3.65e-21
C4303 check[2] a_9152_4775# 0.00242f
C4304 a_10681_4086# a_11629_4386# 7.74e-21
C4305 a_2697_5083# a_3453_4801# 4.06e-20
C4306 a_2463_4775# a_2398_4801# 4.2e-20
C4307 a_2289_4801# a_2579_4801# 0.0282f
C4308 a_1616_4801# x20.Q_N 4.31e-20
C4309 x7.X x75.Q_N 1.48e-19
C4310 a_6011_4801# a_8237_4801# 4e-20
C4311 a_5845_4801# a_8403_4801# 2.9e-21
C4312 a_10156_4112# a_9638_3213# 2.07e-19
C4313 a_5169_2732# a_5371_2366# 8.94e-19
C4314 check[5] a_6984_2366# 9.43e-20
C4315 VDD a_3671_5674# 7.34e-19
C4316 a_4453_2340# a_4592_2366# 2.56e-19
C4317 a_3912_2366# a_6304_2366# 8.41e-21
C4318 a_8236_3239# a_8402_3239# 0.782f
C4319 a_4452_2640# a_4793_2366# 0.00118f
C4320 a_4154_2340# a_5991_2340# 1.86e-21
C4321 x33.Q_N a_8857_3213# 5.46e-19
C4322 a_10629_4801# a_10795_4801# 0.751f
C4323 a_7480_3521# a_8236_3239# 4.06e-20
C4324 eob a_897_4112# 0.0036f
C4325 a_3913_4112# a_4113_4394# 0.00185f
C4326 a_3600_4086# a_4389_4478# 7.71e-20
C4327 VDD a_6846_4086# 0.805f
C4328 x4.X x42.Q_N 0.252f
C4329 a_3913_4112# x7.X 2.29e-20
C4330 x5.X a_3170_4801# 0.0367f
C4331 a_897_4112# x4.A 0.238f
C4332 a_8403_4801# a_8384_4086# 6.63e-19
C4333 a_8237_4801# a_8697_4112# 3.05e-19
C4334 check[0] a_6985_4112# 3.21e-20
C4335 a_3648_5972# a_3373_5674# 0.0156f
C4336 sel_bit[0] a_2463_4775# 5.11e-20
C4337 x39.Q_N D[1] 3.4e-19
C4338 D[5] a_6780_2366# 3.51e-20
C4339 sel_bit[1] a_3258_5648# 0.259f
C4340 a_6546_2340# a_6982_2732# 0.00412f
C4341 a_6304_2366# a_6410_2366# 0.0552f
C4342 a_6844_2640# a_6780_2732# 2.13e-19
C4343 a_6845_2340# a_6504_2648# 1.25e-19
C4344 check[3] a_11630_4086# 0.223f
C4345 a_3452_3239# a_3912_2366# 1.89e-19
C4346 a_3618_3239# a_3599_2340# 3.73e-19
C4347 a_7362_3239# a_7317_2550# 1.01e-20
C4348 x4.X a_4113_4394# 1.78e-19
C4349 x33.Q_N a_8383_2340# 0.142f
C4350 x4.X x7.X 0.88f
C4351 eob D[7] 2.2e-20
C4352 VDD a_3599_2340# 0.58f
C4353 x5.X a_6292_5167# 0.00462f
C4354 a_1511_4112# a_2060_2640# 0.00164f
C4355 a_5845_4801# a_7073_4801# 0.0334f
C4356 check[0] a_3900_5167# 8.76e-19
C4357 a_6466_4775# a_6760_4775# 0.199f
C4358 a_6011_4801# a_7247_4775# 0.0264f
C4359 a_4453_4386# x77.Y 1.11e-20
C4360 x20.Q_N a_2979_2366# 0.00156f
C4361 a_6984_2366# a_7185_2366# 3.34e-19
C4362 a_8288_2340# a_8696_2366# 6.04e-19
C4363 a_9639_4775# a_10795_4801# 1.25e-19
C4364 a_9465_4801# a_10629_4801# 6.38e-20
C4365 a_10628_3239# a_11714_3521# 0.00907f
C4366 a_10794_3239# a_11493_3521# 2.46e-19
C4367 check[1] x72.Q_N 4.68e-20
C4368 x5.X a_9237_4386# 0.00958f
C4369 x4.X a_1207_2340# 0.117f
C4370 VDD a_6982_2732# 0.0163f
C4371 x27.D a_3807_4801# 0.164f
C4372 x7.X a_4657_2340# 0.00586f
C4373 VDD a_9550_3605# 0.00371f
C4374 a_10776_4086# a_11289_4394# 0.00945f
C4375 x5.X a_11629_2340# 4.23e-20
C4376 x42.Q_N x69.Q_N 3.92e-19
C4377 x30.Q_N a_9441_2340# 9.31e-21
C4378 a_12030_3213# a_11833_2340# 2.52e-19
C4379 a_11543_3213# a_12101_2550# 1.62e-19
C4380 VDD a_7562_4478# 0.0042f
C4381 x4.X a_9173_4112# 8.4e-20
C4382 check[1] a_8383_2340# 0.0126f
C4383 x4.X a_4018_2366# 3.78e-20
C4384 x7.A x7.X 0.00565f
C4385 a_7186_4112# x42.Q_N 4.05e-20
C4386 a_5562_4801# a_4454_4086# 6.67e-19
C4387 check[6] a_4453_4386# 0.0318f
C4388 a_8939_4086# a_9238_4086# 0.0334f
C4389 a_8697_4112# a_9442_4086# 0.199f
C4390 a_8384_4086# a_9710_4296# 4.7e-22
C4391 x7.X D[4] 0.00125f
C4392 x4.X a_6605_3239# 0.00267f
C4393 a_897_4112# a_929_3238# 0.00635f
C4394 x7.X a_11249_3213# 4.81e-19
C4395 a_4368_4775# a_6199_4801# 1.49e-21
C4396 x45.Q_N a_8236_3239# 1.49e-19
C4397 a_4855_4775# a_7073_4801# 1.86e-21
C4398 x7.X x69.Q_N 1.46e-19
C4399 check[0] a_7562_4112# 5.56e-22
C4400 a_3453_4801# a_3452_3239# 6.9e-19
C4401 x5.X a_11160_5167# 4.21e-19
C4402 x45.Q_N a_6977_3239# 0.00399f
C4403 a_2533_2550# a_2401_2366# 0.0258f
C4404 a_9152_4775# a_8591_4801# 2.47e-21
C4405 a_8684_5167# a_8768_5167# 0.00972f
C4406 a_6465_3213# a_6291_3605# 0.205f
C4407 a_2060_2640# a_4154_2340# 4.16e-20
C4408 a_6010_3239# a_6759_3213# 0.139f
C4409 a_9639_4775# a_9465_4801# 0.197f
C4410 a_5844_3239# a_7246_3213# 0.0492f
C4411 a_2061_2340# a_3912_2366# 3.12e-19
C4412 a_8237_4801# a_9102_5083# 0.00276f
C4413 a_11088_2366# x63.Q_N 0.00553f
C4414 a_11628_2640# a_11833_2340# 0.153f
C4415 a_2883_5674# x48.Q 0.00144f
C4416 VDD a_1616_4801# 6e-19
C4417 x4.X a_8288_2340# 0.00317f
C4418 check[2] a_7954_4801# 4.53e-20
C4419 x7.X a_10775_2340# 0.00442f
C4420 a_3600_4086# a_4213_3239# 1.16e-20
C4421 a_4926_4296# a_4680_3239# 2.37e-20
C4422 a_929_3238# D[7] 0.00104f
C4423 a_4453_2340# a_4871_2648# 0.00276f
C4424 a_3912_2366# D[5] 2.89e-20
C4425 a_4452_2640# a_5169_2732# 4.45e-20
C4426 check[1] a_3600_4086# 1.19e-20
C4427 a_2853_5648# a_3913_4112# 4.72e-21
C4428 a_6291_3605# a_5991_2340# 3.9e-20
C4429 a_5844_3239# a_6844_2640# 6.01e-20
C4430 a_6465_3213# a_6304_2366# 0.0014f
C4431 check[0] a_6844_2640# 2.7e-19
C4432 a_1511_4112# a_3505_4086# 0.0121f
C4433 check[2] a_9578_4112# 1.87e-19
C4434 x5.X a_9656_4394# 2.97e-19
C4435 x20.Q_N a_4591_4478# 6.94e-20
C4436 a_4074_4775# a_4214_4801# 0.07f
C4437 a_3619_4801# a_4008_4801# 0.0019f
C4438 a_3453_4801# a_4586_4801# 2.56e-19
C4439 a_4368_4775# a_4539_5083# 0.00652f
C4440 check[2] a_8236_3239# 6.24e-22
C4441 x4.X a_4766_3605# 6.48e-19
C4442 check[5] a_8289_4086# 0.00275f
C4443 x5.X a_9551_5167# 1.06e-19
C4444 x20.Q_N a_4214_4801# 1.27e-19
C4445 a_2853_5648# x4.X 5.73e-20
C4446 D[5] a_6410_2366# 5.42e-19
C4447 a_7073_4801# a_7182_4801# 0.00707f
C4448 a_5991_2340# a_6304_2366# 0.273f
C4449 a_8236_3239# a_10628_3239# 0.00176f
C4450 a_3452_3239# D[6] 2.82e-19
C4451 x33.Q_N a_7763_2366# 1.34e-20
C4452 x33.Q_N a_10794_3239# 3.79e-20
C4453 a_8236_3239# a_9369_3239# 2.56e-19
C4454 a_8402_3239# a_8791_3239# 0.0019f
C4455 a_8857_3213# a_8997_3239# 0.07f
C4456 a_9151_3213# a_9322_3521# 0.00652f
C4457 x77.Y a_5561_3239# 3.29e-19
C4458 a_1227_4801# a_1511_4112# 0.00301f
C4459 x5.A sel_bit[1] 0.0352f
C4460 a_10795_4801# a_11184_4801# 0.0019f
C4461 a_11544_4775# a_11715_5083# 0.00652f
C4462 a_10629_4801# a_11762_4801# 2.56e-19
C4463 a_11250_4775# a_11390_4801# 0.07f
C4464 a_4454_4086# a_6305_4112# 5.07e-21
C4465 a_4453_4386# a_6547_4086# 2.47e-20
C4466 a_4926_4296# a_4794_4112# 0.0258f
C4467 VDD a_2979_2366# 0.117f
C4468 VDD a_9152_4775# 0.449f
C4469 VDD a_6010_3239# 0.274f
C4470 a_8697_4112# a_10156_4112# 8.23e-22
C4471 a_9442_4086# a_9375_4478# 9.46e-19
C4472 x42.Q_N a_8897_4394# 2.02e-20
C4473 a_9237_4386# a_9656_4394# 2.46e-19
C4474 check[6] a_6011_4801# 0.162f
C4475 x20.Q_N a_1762_2340# 0.162f
C4476 x39.Q_N a_12737_3239# 3.23e-19
C4477 D[4] a_8288_2340# 0.1f
C4478 a_1061_4801# a_1227_4801# 0.619f
C4479 a_8403_4801# check[4] 1.14e-20
C4480 eob a_1415_4801# 0.151f
C4481 D[1] a_10982_3239# 4.96e-19
C4482 a_8997_3239# a_8383_2340# 4.6e-20
C4483 x33.Q_N a_9577_2366# 0.0403f
C4484 a_12738_4801# a_12030_3213# 3.19e-20
C4485 check[3] a_11543_3213# 1.04e-19
C4486 x4.X a_6846_4086# 0.0467f
C4487 a_7318_4296# x45.Q_N 0.00243f
C4488 VDD a_4793_2366# 9.91e-19
C4489 check[0] a_5372_4112# 0.165f
C4490 a_3913_4112# a_3599_2340# 5.05e-21
C4491 x7.X a_7072_3239# 1.93e-19
C4492 x5.X x30.Q_N 8.83e-19
C4493 a_9238_4086# D[1] 3.36e-19
C4494 a_6760_4775# a_7481_5083# 0.00185f
C4495 a_6292_5167# x30.Q_N 7.29e-20
C4496 a_10629_4801# a_11089_4112# 3.05e-19
C4497 check[0] x27.Q_N 0.0367f
C4498 a_10795_4801# a_10776_4086# 6.63e-19
C4499 check[6] a_5561_3239# 0.027f
C4500 x27.Q_N a_5844_3239# 8.96e-20
C4501 a_1062_5674# eob 4.55e-20
C4502 x33.Q_N a_11076_5167# 1.6e-19
C4503 check[3] a_11330_2340# 1.32e-19
C4504 check[2] a_1511_4112# 5.19e-20
C4505 sel_bit[1] x27.D 4.45e-19
C4506 a_1062_5674# x4.A 8.16e-22
C4507 VDD a_4971_4801# 0.0111f
C4508 check[2] a_11289_4394# 9.25e-20
C4509 VDD a_9172_2732# 0.00371f
C4510 x4.X a_3599_2340# 0.117f
C4511 x48.Q a_2289_4801# 8.99e-20
C4512 a_4681_4801# check[6] 4.98e-20
C4513 VDD a_11714_3521# 0.0163f
C4514 x7.X a_6845_2340# 0.182f
C4515 a_12102_4296# a_11970_4112# 0.0258f
C4516 x39.Q_N a_11769_4112# 0.00167f
C4517 x27.Q_N a_4592_2366# 0.00474f
C4518 check[5] a_9465_4801# 6.82e-20
C4519 a_2265_2340# a_2979_2366# 6.99e-20
C4520 a_2061_2340# D[6] 0.338f
C4521 a_2533_2550# a_2777_2732# 0.00972f
C4522 check[1] a_6985_4112# 7.78e-20
C4523 D[3] x63.Q_N 0.00107f
C4524 x5.X a_3373_5674# 1.23e-19
C4525 a_1338_5674# a_1682_4775# 0.00186f
C4526 a_2389_5648# a_1227_4801# 3.08e-19
C4527 a_11857_4801# check[3] 0.00257f
C4528 clk_sar a_1061_4801# 1.18e-19
C4529 x5.X a_5992_4086# 0.0202f
C4530 check[1] a_9577_2366# 4.4e-19
C4531 check[2] a_7318_4296# 2.18e-22
C4532 a_4453_4386# a_6411_4112# 9.75e-21
C4533 x4.X a_6982_2732# 9.81e-19
C4534 x48.Q a_4454_4086# 2.06e-19
C4535 a_5845_4801# a_6845_4386# 9.86e-20
C4536 a_6466_4775# a_6305_4112# 0.0025f
C4537 a_6292_5167# a_5992_4086# 4.9e-20
C4538 a_1508_5167# a_1616_4801# 0.00812f
C4539 a_2463_4775# a_2375_5167# 7.71e-20
C4540 a_2289_4801# a_2147_5083# 0.00412f
C4541 x7.X a_10155_2366# 0.155f
C4542 x4.X a_9550_3605# 4.4e-19
C4543 a_1976_4775# a_1822_4801# 0.00943f
C4544 a_6846_4086# D[4] 1.26e-20
C4545 x7.X a_3899_3605# 1.95e-19
C4546 sel_bit[0] a_897_4112# 8.65e-21
C4547 check[5] a_6304_2366# 1.15e-20
C4548 a_12547_2366# a_12345_2366# 3.67e-19
C4549 a_11564_2366# a_11969_2366# 2.46e-21
C4550 a_9465_4801# a_8402_3239# 6.75e-21
C4551 a_6759_3213# a_8236_3239# 3.41e-19
C4552 a_3912_2366# a_4453_2340# 0.125f
C4553 a_4154_2340# a_4452_2640# 0.137f
C4554 eob a_3170_4801# 0.00132f
C4555 check[1] a_3900_5167# 4.17e-20
C4556 a_6759_3213# a_6977_3239# 3.73e-19
C4557 a_7072_3239# a_6605_3239# 0.00316f
C4558 VDD a_4591_4478# 0.0172f
C4559 x4.X a_7562_4478# 9.15e-19
C4560 a_3453_4801# a_3600_4086# 0.00159f
C4561 VDD a_4214_4801# 0.035f
C4562 a_6845_4386# a_8384_4086# 2.16e-19
C4563 a_6846_4086# a_7186_4112# 6.04e-20
C4564 a_7050_4086# a_6985_4112# 9.75e-19
C4565 x45.Q_N a_8289_4086# 8.9e-21
C4566 x20.Q_N a_1511_4112# 0.0407f
C4567 a_1415_4801# a_929_3238# 4.09e-20
C4568 VDD a_11390_4801# 0.0332f
C4569 a_6710_5083# check[5] 3.95e-22
C4570 a_5371_2366# a_6304_2366# 3.42e-20
C4571 x5.X eob 0.155f
C4572 D[5] a_5991_2340# 0.0123f
C4573 x33.Q_N a_6844_2640# 0.00104f
C4574 a_1227_4801# a_3619_4801# 7.69e-21
C4575 x77.Y a_4854_3213# 0.142f
C4576 a_2389_5648# check[2] 0.138f
C4577 a_5897_4086# x7.X 2.05e-21
C4578 a_1061_4801# x20.Q_N 2.14e-19
C4579 a_1682_4775# a_2194_4801# 9.75e-19
C4580 x5.X x4.A 5.96e-19
C4581 VDD a_7954_4801# 0.193f
C4582 VDD a_1762_2340# 0.201f
C4583 a_11565_4112# a_11970_4112# 2.46e-21
C4584 a_12548_4112# a_12346_4112# 3.67e-19
C4585 x39.Q_N a_10982_3239# 7.52e-20
C4586 a_10776_4086# a_11389_3239# 1.16e-20
C4587 a_6845_2340# a_8288_2340# 8.18e-19
C4588 check[1] a_7562_4112# 1.69e-19
C4589 a_6546_2340# a_6984_2366# 0.00276f
C4590 a_6304_2366# a_7185_2366# 0.00943f
C4591 a_9638_3213# a_9573_3239# 4.2e-20
C4592 a_9464_3239# a_9754_3239# 0.0282f
C4593 x75.Q_N a_6010_3239# 2.12e-19
C4594 check[1] a_7246_3213# 0.00245f
C4595 x5.X a_6781_4478# 3.2e-19
C4596 VDD a_9578_4112# 0.0326f
C4597 check[2] a_8289_4086# 1.35e-21
C4598 sel_bit[0] a_3648_5972# 2.6e-19
C4599 VDD a_5169_2732# 0.00436f
C4600 VDD a_8236_3239# 0.791f
C4601 VDD a_6977_3239# 6.2e-19
C4602 check[0] a_4155_4086# 4.34e-20
C4603 a_9238_4086# x39.Q_N 3.57e-19
C4604 x5.X D[2] 0.0046f
C4605 check[6] a_6978_4801# 6.18e-20
C4606 check[4] a_10681_4086# 0.00276f
C4607 a_9710_4296# a_9464_3239# 2.37e-20
C4608 x42.Q_N a_9638_3213# 0.144f
C4609 x20.Q_N a_4154_2340# 2.93e-20
C4610 x39.Q_N a_11833_2340# 1.11e-19
C4611 check[6] a_4854_3213# 0.00397f
C4612 a_8696_2366# a_9172_2732# 0.00133f
C4613 a_9370_4801# check[4] 9.79e-21
C4614 a_11856_3239# D[2] 5.2e-20
C4615 check[1] a_6844_2640# 7.55e-20
C4616 check[2] a_3619_4801# 6.48e-20
C4617 x4.X a_2979_2366# 4.09e-19
C4618 x4.X a_6010_3239# 0.0446f
C4619 x4.X a_9152_4775# 0.104f
C4620 x5.X a_1926_5083# 3.49e-19
C4621 a_11630_4086# x7.X 3e-20
C4622 a_2389_5648# x20.Q_N 2.12e-20
C4623 VDD a_6984_2366# 6.2e-19
C4624 x7.X a_9638_3213# 0.00374f
C4625 check[2] a_10795_4801# 0.00106f
C4626 a_7318_4296# a_6759_3213# 1.71e-19
C4627 a_7050_4086# a_7246_3213# 2.47e-19
C4628 x45.Q_N a_6291_3605# 0.152f
C4629 a_9710_4296# a_9237_2340# 6.08e-21
C4630 x42.Q_N a_9236_2640# 4.61e-20
C4631 a_1207_2340# x51.Q_N 0.124f
C4632 a_1762_2340# a_2265_2340# 0.00187f
C4633 a_1520_2366# a_2533_2550# 0.0633f
C4634 a_2060_2640# a_2061_2340# 0.783f
C4635 a_10795_4801# a_10628_3239# 9.04e-19
C4636 a_10629_4801# a_10794_3239# 8.16e-19
C4637 D[2] a_11629_2340# 0.271f
C4638 a_9237_2340# x63.Q_N 2.94e-19
C4639 check[1] a_7159_5167# 1.92e-19
C4640 a_3618_3239# a_4007_3239# 0.0019f
C4641 x33.Q_N x36.Q_N 2.37e-20
C4642 a_3452_3239# a_4585_3239# 2.56e-19
C4643 a_4367_3213# a_4538_3521# 0.00652f
C4644 a_4073_3213# a_4213_3239# 0.07f
C4645 x5.X a_929_3238# 2.33e-20
C4646 VDD a_11288_2648# 0.00506f
C4647 x48.Q a_3807_4801# 0.00791f
C4648 VDD a_4007_3239# 2.82e-19
C4649 x7.X a_9236_2640# 0.108f
C4650 a_6845_4386# a_7049_2340# 1.26e-21
C4651 a_6846_4086# a_6845_2340# 1.55e-19
C4652 x45.Q_N a_6304_2366# 6.37e-20
C4653 a_3505_4086# a_3452_3239# 5.06e-19
C4654 x27.Q_N a_6780_2366# 9.28e-21
C4655 D[6] a_4453_2340# 2.08e-19
C4656 a_5844_3239# a_7953_3239# 1.03e-19
C4657 a_11629_2340# a_11969_2366# 6.04e-20
C4658 a_11833_2340# a_11768_2366# 9.75e-19
C4659 check[5] x72.Q_N 0.00322f
C4660 a_11628_2640# a_12345_2366# 0.00105f
C4661 VDD a_1511_4112# 1.55f
C4662 VDD a_11289_4394# 0.00506f
C4663 x4.X a_4971_4801# 0.00557f
C4664 x4.X a_9172_2732# 4.32e-19
C4665 a_3619_4801# a_4074_4775# 0.153f
C4666 a_3453_4801# a_3900_5167# 0.15f
C4667 check[2] a_9465_4801# 0.00105f
C4668 x7.X a_12345_2732# 8.26e-19
C4669 x4.X a_11714_3521# 9.99e-19
C4670 x20.Q_N a_3619_4801# 4.85e-19
C4671 x5.X a_8237_4801# 0.27f
C4672 a_10776_4086# a_11089_4112# 0.272f
C4673 a_2697_5083# x20.Q_N 2.02e-20
C4674 a_5845_4801# a_5844_3239# 6.9e-19
C4675 a_2853_5648# a_2784_5996# 0.00105f
C4676 check[0] a_5845_4801# 0.00285f
C4677 check[5] a_8383_2340# 3.32e-21
C4678 a_4452_2640# a_6304_2366# 1.95e-19
C4679 a_8236_3239# a_8683_3605# 0.15f
C4680 x27.Q_N a_4213_3239# 6.11e-19
C4681 VDD a_1061_4801# 0.901f
C4682 a_4657_2340# a_4793_2366# 0.07f
C4683 a_4453_2340# a_5991_2340# 0.00116f
C4684 a_8402_3239# a_8857_3213# 0.153f
C4685 a_10629_4801# a_11076_5167# 0.15f
C4686 a_10795_4801# a_11250_4775# 0.153f
C4687 x72.Q_N a_8402_3239# 9.24e-20
C4688 x33.Q_N a_9151_3213# 0.00498f
C4689 check[1] x27.Q_N 3.1e-20
C4690 a_3600_4086# a_4019_4112# 0.0397f
C4691 a_7480_3521# x72.Q_N 2.02e-20
C4692 VDD a_7318_4296# 0.317f
C4693 a_4155_4086# a_4389_4478# 0.00976f
C4694 a_3913_4112# a_4591_4478# 0.00652f
C4695 a_4453_4386# x7.X 2.5e-20
C4696 a_7764_4112# a_7562_4112# 3.67e-19
C4697 a_8858_4775# a_8697_4112# 0.0025f
C4698 a_8237_4801# a_9237_4386# 9.86e-20
C4699 a_8684_5167# a_8384_4086# 4.9e-20
C4700 a_7764_4112# a_7246_3213# 2.07e-19
C4701 a_9578_4112# a_8696_2366# 1.26e-20
C4702 D[5] a_7185_2366# 7.82e-20
C4703 a_6845_2340# a_6982_2732# 0.00907f
C4704 a_2883_5674# a_2993_5674# 0.00857f
C4705 D[7] a_2200_2366# 3.49e-19
C4706 check[3] a_12102_4296# 0.00213f
C4707 a_8402_3239# a_8383_2340# 3.73e-19
C4708 a_8236_3239# a_8696_2366# 1.89e-19
C4709 D[0] a_9573_3239# 1.29e-20
C4710 x4.X a_4591_4478# 0.00114f
C4711 a_3452_3239# a_4452_2640# 6.01e-20
C4712 a_3899_3605# a_3599_2340# 3.9e-20
C4713 a_4073_3213# a_3912_2366# 0.0014f
C4714 x33.Q_N a_8938_2340# 0.16f
C4715 a_5897_4086# a_6846_4086# 7e-20
C4716 x4.X a_4214_4801# 7.25e-19
C4717 VDD a_4154_2340# 0.182f
C4718 x5.X a_7247_4775# 0.00983f
C4719 x4.X a_11390_4801# 7.25e-19
C4720 a_1511_4112# a_2265_2340# 0.00119f
C4721 a_6011_4801# a_6199_4801# 0.162f
C4722 a_1062_5674# sel_bit[0] 0.0421f
C4723 a_6466_4775# a_7073_4801# 0.00187f
C4724 a_6292_5167# a_7247_4775# 4.7e-22
C4725 a_5845_4801# a_6376_5167# 0.0018f
C4726 check[0] a_4855_4775# 0.0127f
C4727 x42.Q_N D[0] 3.91e-19
C4728 a_4658_4086# x77.Y 1.87e-21
C4729 a_8288_2340# a_9236_2640# 9.02e-21
C4730 a_9639_4775# a_11076_5167# 7.98e-21
C4731 x75.Q a_5896_2340# 0.00129f
C4732 x30.Q_N a_7362_3239# 0.00342f
C4733 a_10628_3239# a_11389_3239# 6.04e-20
C4734 a_11249_3213# a_11714_3521# 9.46e-19
C4735 a_12738_4801# a_12737_3239# 9.85e-20
C4736 a_10794_3239# a_11942_3605# 2.13e-19
C4737 VDD a_2389_5648# 0.695f
C4738 check[1] a_9151_3213# 1.78e-20
C4739 x4.X a_7954_4801# 0.00672f
C4740 VDD a_7263_2648# 0.00984f
C4741 x4.X a_1762_2340# 0.00671f
C4742 x5.X a_9442_4086# 9.38e-19
C4743 x7.X D[0] 0.0253f
C4744 x7.X x54.Q_N 0.00122f
C4745 eob a_3373_5674# 1.33e-19
C4746 a_11089_4112# a_11565_4478# 0.00133f
C4747 x27.Q_N a_3912_2366# 0.0928f
C4748 x30.Q_N x60.Q_N 8.43e-20
C4749 check[3] a_11564_2366# 2.19e-20
C4750 a_11856_3239# a_12101_2550# 1.85e-20
C4751 VDD a_8289_4086# 0.189f
C4752 x4.X a_9578_4112# 0.0031f
C4753 check[1] a_8938_2340# 0.00112f
C4754 x4.X a_5169_2732# 1.17e-19
C4755 a_6011_4801# x7.X 2.9e-21
C4756 x4.X a_8236_3239# 0.0456f
C4757 a_8697_4112# x42.Q_N 0.0927f
C4758 a_9237_4386# a_9442_4086# 0.153f
C4759 x4.X a_6977_3239# 4.96e-19
C4760 a_4368_4775# a_4971_4801# 0.0552f
C4761 x7.X a_11543_3213# 6.77e-19
C4762 a_3619_4801# a_3618_3239# 1.39e-19
C4763 x5.X a_9574_4801# 5.36e-20
C4764 x45.Q_N x72.Q_N 3.9e-19
C4765 x27.Q_N a_6410_2366# 8.39e-20
C4766 x20.Q_N a_3452_3239# 0.00411f
C4767 a_3170_4801# x77.Y 5.69e-20
C4768 a_8858_4775# a_9102_5083# 0.0104f
C4769 a_8403_4801# a_9323_5083# 1.09e-19
C4770 a_6291_3605# a_6759_3213# 0.0633f
C4771 a_2060_2640# a_4453_2340# 2.9e-21
C4772 a_2533_2550# a_3912_2366# 6.92e-21
C4773 a_2061_2340# a_4452_2640# 4e-20
C4774 a_5844_3239# a_6198_3239# 0.0708f
C4775 a_6010_3239# a_7072_3239# 0.137f
C4776 check[0] a_6198_3239# 0.00621f
C4777 a_2853_5648# a_2463_4775# 9.54e-20
C4778 a_11629_2340# a_12101_2550# 0.15f
C4779 a_11628_2640# x63.Q_N 5.46e-21
C4780 x48.Q a_3258_5648# 0.00631f
C4781 a_5992_4086# a_6781_4478# 7.71e-20
C4782 a_6305_4112# a_6505_4394# 0.00185f
C4783 VDD a_3619_4801# 0.617f
C4784 sel_bit[1] x48.Q 0.173f
C4785 VDD a_2697_5083# 0.00615f
C4786 a_1508_5167# a_1511_4112# 3.47e-19
C4787 a_8697_4112# x7.X 2.29e-20
C4788 VDD a_10795_4801# 0.593f
C4789 x7.X a_5561_3239# 0.00108f
C4790 x7.X a_11330_2340# 0.00103f
C4791 sel_bit[0] x5.X 0.0929f
C4792 check[5] a_7763_2366# 0.0034f
C4793 a_4657_2340# a_5169_2732# 6.69e-20
C4794 eob x4.A 0.0197f
C4795 a_4452_2640# D[5] 0.00524f
C4796 a_4453_2340# a_5371_2366# 0.0708f
C4797 a_5844_3239# a_7049_2340# 4.77e-19
C4798 a_6465_3213# a_6844_2640# 2.68e-19
C4799 a_6291_3605# a_6546_2340# 2.41e-20
C4800 a_6759_3213# a_6304_2366# 3.36e-20
C4801 check[0] a_7049_2340# 4.27e-19
C4802 a_6010_3239# a_6845_2340# 6.38e-20
C4803 a_6605_3239# D[0] 1.08e-20
C4804 x36.Q_N a_10680_2340# 3.7e-19
C4805 a_1061_4801# a_1508_5167# 0.138f
C4806 a_1511_4112# a_3913_4112# 1e-19
C4807 a_3505_4086# a_3600_4086# 0.0968f
C4808 x5.X a_10156_4112# 9.37e-19
C4809 check[2] a_11089_4112# 0.00131f
C4810 x4.X a_11288_2648# 0.00102f
C4811 x4.X a_4007_3239# 6.32e-19
C4812 a_4368_4775# a_4214_4801# 0.00943f
C4813 a_3900_5167# a_4008_4801# 0.00812f
C4814 a_3453_4801# x27.Q_N 2.36e-19
C4815 a_4681_4801# a_4539_5083# 0.00412f
C4816 a_4855_4775# a_4767_5167# 7.71e-20
C4817 a_4074_4775# a_4586_4801# 9.75e-19
C4818 x5.X a_8792_4801# 2.86e-19
C4819 x20.Q_N a_4586_4801# 5.69e-20
C4820 a_10776_4086# a_10794_3239# 3.48e-19
C4821 a_11089_4112# a_10628_3239# 2.21e-19
C4822 x30.Q_N a_8237_4801# 3.15e-19
C4823 a_8236_3239# D[4] 5.41e-19
C4824 D[0] a_8288_2340# 0.00665f
C4825 a_5896_2340# x57.Q_N 0.178f
C4826 a_6304_2366# a_6546_2340# 0.124f
C4827 a_5991_2340# a_6844_2640# 0.0264f
C4828 a_4367_3213# a_5844_3239# 3.41e-19
C4829 check[0] a_4367_3213# 2.58e-20
C4830 a_8857_3213# a_9369_3239# 9.75e-19
C4831 a_9638_3213# a_9550_3605# 7.71e-20
C4832 a_9151_3213# a_8997_3239# 0.00943f
C4833 a_8236_3239# x69.Q_N 1.07e-19
C4834 x4.X a_1511_4112# 1.74f
C4835 a_8683_3605# a_8791_3239# 0.00812f
C4836 a_9464_3239# a_9322_3521# 0.00412f
C4837 a_11250_4775# a_11762_4801# 9.75e-19
C4838 a_10629_4801# x36.Q_N 1.22e-19
C4839 a_11544_4775# a_11390_4801# 0.00943f
C4840 a_11076_5167# a_11184_4801# 0.00812f
C4841 a_11857_4801# a_11715_5083# 0.00412f
C4842 a_12031_4775# a_11943_5167# 7.71e-20
C4843 x4.X a_11289_4394# 1.75e-19
C4844 a_4453_4386# a_6846_4086# 2.9e-21
C4845 a_9237_4386# a_10156_4112# 0.162f
C4846 VDD a_6291_3605# 0.176f
C4847 VDD a_9465_4801# 0.343f
C4848 a_8697_4112# a_9173_4112# 2.87e-21
C4849 a_9442_4086# a_9656_4394# 0.0104f
C4850 a_9238_4086# a_9954_4478# 0.0018f
C4851 x5.X check[6] 0.168f
C4852 check[6] a_6292_5167# 0.00105f
C4853 x5.X check[3] 0.285f
C4854 x20.Q_N a_2061_2340# 0.0469f
C4855 a_1227_4801# a_1682_4775# 0.145f
C4856 a_8684_5167# check[4] 4.29e-21
C4857 a_9152_4775# a_10346_4801# 6.04e-19
C4858 a_7317_2550# a_7561_2366# 0.00812f
C4859 a_1061_4801# x4.X 0.0131f
C4860 D[1] a_9754_3239# 8.74e-20
C4861 eob a_1926_5083# 0.00171f
C4862 x33.Q_N a_11088_2366# 8.24e-20
C4863 x4.X a_7318_4296# 0.0211f
C4864 check[1] a_7953_3239# 0.00311f
C4865 VDD a_6304_2366# 0.348f
C4866 check[0] a_4389_4112# 8.48e-21
C4867 x27.Q_N D[6] 0.00313f
C4868 x42.Q_N a_10345_3239# 3.23e-19
C4869 a_7247_4775# x30.Q_N 0.126f
C4870 a_11076_5167# a_10776_4086# 4.9e-20
C4871 a_11250_4775# a_11089_4112# 0.0025f
C4872 a_10629_4801# a_11629_4386# 9.86e-20
C4873 eob a_929_3238# 0.0549f
C4874 a_8696_2366# a_9172_2366# 2.87e-21
C4875 a_3452_3239# a_3618_3239# 0.638f
C4876 check[1] a_5845_4801# 5.4e-19
C4877 check[3] a_11629_2340# 0.0405f
C4878 check[2] a_3600_4086# 1.65e-20
C4879 VDD a_8802_2366# 4.84e-19
C4880 a_897_4112# x7.X 4.72e-19
C4881 check[2] a_11767_4478# 5.02e-20
C4882 VDD a_6710_5083# 0.00984f
C4883 x4.A a_929_3238# 3.84e-19
C4884 x4.X a_4154_2340# 0.00377f
C4885 VDD a_3452_3239# 0.821f
C4886 x7.X a_10345_3239# 0.00106f
C4887 a_6846_4086# D[0] 3.2e-19
C4888 VDD a_11389_3239# 5.47e-21
C4889 x7.X a_7317_2550# 0.00825f
C4890 x39.Q_N a_12346_4112# 2.43e-19
C4891 x27.Q_N a_5991_2340# 1.43e-19
C4892 check[5] a_7246_3213# 0.00432f
C4893 a_2533_2550# D[6] 0.00108f
C4894 a_10775_2340# a_11288_2648# 0.00945f
C4895 check[1] a_8384_4086# 0.0126f
C4896 a_2389_5648# x4.X 0.00219f
C4897 x77.Y a_4789_3239# 7.87e-19
C4898 a_11160_5167# check[3] 1.13e-19
C4899 x5.X a_6547_4086# 0.00115f
C4900 x4.X a_7263_2648# 2.86e-19
C4901 x48.Q a_4926_4296# 1.36e-19
C4902 a_5845_4801# a_7050_4086# 6.96e-19
C4903 a_6760_4775# a_6305_4112# 5.67e-20
C4904 a_6292_5167# a_6547_4086# 2.46e-20
C4905 a_6466_4775# a_6845_4386# 3.92e-19
C4906 a_6011_4801# a_6846_4086# 1.18e-19
C4907 a_1976_4775# a_3453_4801# 1.75e-19
C4908 x4.X a_8791_3239# 6.32e-19
C4909 a_2289_4801# a_1822_4801# 0.00316f
C4910 a_4019_4112# a_4073_3213# 3.34e-20
C4911 a_1976_4775# a_2194_4801# 3.73e-19
C4912 x7.X a_4854_3213# 0.00379f
C4913 x7.X D[7] 9.14e-20
C4914 x27.Q_N a_4790_4801# 8.36e-20
C4915 check[5] a_6844_2640# 0.0314f
C4916 a_9152_4775# a_9638_3213# 1.06e-20
C4917 a_9639_4775# a_9151_3213# 1.08e-22
C4918 a_6759_3213# a_8857_3213# 4.53e-20
C4919 a_7246_3213# a_8402_3239# 1.84e-19
C4920 a_7072_3239# a_8236_3239# 6.38e-20
C4921 a_4154_2340# a_4657_2340# 0.00187f
C4922 a_3912_2366# a_4925_2550# 0.0633f
C4923 a_3599_2340# x54.Q_N 0.124f
C4924 a_4452_2640# a_4453_2340# 0.781f
C4925 check[1] a_4855_4775# 1.73e-19
C4926 a_6198_3239# a_6399_3239# 3.67e-19
C4927 a_7072_3239# a_6977_3239# 0.00276f
C4928 a_7246_3213# a_7480_3521# 0.00945f
C4929 a_6759_3213# x72.Q_N 0.00553f
C4930 VDD a_4872_4394# 0.0102f
C4931 x4.X a_8289_4086# 0.00368f
C4932 a_4074_4775# a_3600_4086# 4.54e-19
C4933 a_6845_4386# a_8939_4086# 3.16e-20
C4934 VDD a_4586_4801# 0.00495f
C4935 a_3619_4801# a_3913_4112# 9.06e-19
C4936 a_7318_4296# a_7186_4112# 0.0258f
C4937 x45.Q_N a_6985_4112# 0.00166f
C4938 a_6846_4086# a_8697_4112# 5.07e-21
C4939 x20.Q_N a_3600_4086# 0.00304f
C4940 VDD a_11762_4801# 0.00445f
C4941 a_10681_4086# D[1] 0.00123f
C4942 D[5] a_6546_2340# 2.03e-19
C4943 D[7] a_1207_2340# 0.00629f
C4944 a_1112_2340# a_1520_2366# 6.04e-19
C4945 a_7246_3213# a_7185_2366# 1.2e-20
C4946 x77.Y a_3806_3239# 0.0112f
C4947 x4.X a_3619_4801# 0.00737f
C4948 a_1682_4775# x20.Q_N 1.32e-19
C4949 x27.Q_N a_4019_4112# 2.89e-22
C4950 x4.X a_10795_4801# 0.00496f
C4951 VDD a_2061_2340# 0.853f
C4952 x48.Q x27.D 0.0333f
C4953 check[2] a_10794_3239# 0.0351f
C4954 a_4008_4801# x27.Q_N 4.32e-20
C4955 a_7561_2732# a_7763_2366# 8.94e-19
C4956 a_10628_3239# a_10794_3239# 0.782f
C4957 a_6546_2340# a_8383_2340# 1.86e-21
C4958 x33.Q_N D[3] 0.00525f
C4959 a_6304_2366# a_8696_2366# 5.35e-21
C4960 a_6844_2640# a_7185_2366# 0.00118f
C4961 a_6845_2340# a_6984_2366# 2.56e-19
C4962 a_9872_3521# a_10628_3239# 4.06e-20
C4963 VDD a_11089_4112# 0.448f
C4964 sel_bit[0] a_3373_5674# 0.0563f
C4965 VDD D[5] 0.221f
C4966 VDD a_8857_3213# 0.308f
C4967 a_9710_4296# x39.Q_N 1.29e-19
C4968 a_2147_5083# x27.D 2.85e-21
C4969 VDD x72.Q_N 0.0716f
C4970 check[0] a_4454_4086# 0.44f
C4971 check[6] x30.Q_N 1.48e-21
C4972 a_8384_4086# a_8997_3239# 1.16e-20
C4973 x42.Q_N a_8590_3239# 8.76e-20
C4974 x27.Q_N a_2060_2640# 0.00112f
C4975 a_8696_2366# a_8802_2366# 0.0552f
C4976 a_8938_2340# a_9374_2732# 0.00412f
C4977 D[4] a_9172_2366# 3.13e-20
C4978 a_9237_2340# a_8896_2648# 1.25e-19
C4979 a_9236_2640# a_9172_2732# 2.13e-19
C4980 x33.Q_N check[4] 0.842f
C4981 eob a_2398_4801# 2.92e-19
C4982 a_9754_3239# a_9709_2550# 1.01e-20
C4983 a_7764_4112# a_8384_4086# 8.26e-21
C4984 check[2] a_3900_5167# 5.02e-20
C4985 a_6845_4386# a_8803_4112# 3.66e-20
C4986 x45.Q_N a_7562_4112# 2.38e-19
C4987 x4.X a_6291_3605# 0.0177f
C4988 x4.X a_9465_4801# 0.00321f
C4989 x5.X a_2375_5167# 1.58e-19
C4990 VDD a_8383_2340# 0.561f
C4991 a_3453_4801# a_5845_4801# 0.00176f
C4992 x7.X a_8590_3239# 0.158f
C4993 x45.Q_N a_7246_3213# 0.144f
C4994 a_7363_4801# a_7318_4296# 1.9e-20
C4995 a_7318_4296# a_7072_3239# 2.37e-20
C4996 x27.Q_N a_5371_2366# 0.0318f
C4997 x42.Q_N a_9441_2340# 1.11e-19
C4998 a_1762_2340# x51.Q_N 9.58e-21
C4999 x77.Y a_3504_2340# 3.35e-21
C5000 a_10795_4801# a_11249_3213# 3.18e-21
C5001 a_2061_2340# a_2265_2340# 0.117f
C5002 a_10680_2340# a_11088_2366# 6.04e-19
C5003 a_9376_2366# a_9577_2366# 3.34e-19
C5004 a_2060_2640# a_2533_2550# 0.155f
C5005 a_11076_5167# a_10628_3239# 8.3e-21
C5006 D[2] a_12101_2550# 2.21e-19
C5007 a_3452_3239# x75.Q_N 1.07e-19
C5008 a_4680_3239# a_4538_3521# 0.00412f
C5009 a_3899_3605# a_4007_3239# 0.00812f
C5010 a_4367_3213# a_4213_3239# 0.00943f
C5011 a_4073_3213# a_4585_3239# 9.75e-19
C5012 a_4854_3213# a_4766_3605# 7.71e-20
C5013 sel_bit[0] eob 0.294f
C5014 eob x77.Y 0.05f
C5015 check[6] a_5992_4086# 0.00385f
C5016 VDD a_11766_2732# 0.0163f
C5017 x4.X a_6304_2366# 0.112f
C5018 x48.Q a_2579_4801# 1.65e-19
C5019 a_4971_4801# a_4453_4386# 8.84e-21
C5020 x45.Q_N a_6844_2640# 4.61e-20
C5021 a_7318_4296# a_6845_2340# 6.08e-21
C5022 VDD a_5088_3521# 0.00529f
C5023 a_3913_4112# a_3452_3239# 2.21e-19
C5024 x7.X a_9441_2340# 0.00598f
C5025 a_3600_4086# a_3618_3239# 3.48e-19
C5026 sel_bit[0] x4.A 5.72e-21
C5027 check[5] a_9151_3213# 8.29e-21
C5028 a_6010_3239# D[0] 5.69e-21
C5029 check[4] a_9953_2366# 5.12e-20
C5030 D[6] a_4925_2550# 6.65e-20
C5031 a_12101_2550# a_11969_2366# 0.0258f
C5032 reset a_621_4112# 0.197f
C5033 VDD a_3600_4086# 0.741f
C5034 VDD a_11767_4478# 0.0163f
C5035 x4.X a_8802_2366# 3.78e-20
C5036 a_1415_4801# x7.X 2.3e-21
C5037 a_4074_4775# a_3900_5167# 0.205f
C5038 a_3453_4801# a_4855_4775# 0.0492f
C5039 a_3619_4801# a_4368_4775# 0.139f
C5040 x4.X a_3452_3239# 0.0477f
C5041 x4.X a_11389_3239# 0.00267f
C5042 x5.X a_8858_4775# 0.00316f
C5043 a_10776_4086# a_11629_4386# 0.0264f
C5044 x20.Q_N a_3900_5167# 2.13e-19
C5045 a_10681_4086# x39.Q_N 0.181f
C5046 a_11089_4112# a_11331_4086# 0.124f
C5047 x30.Q_N a_6547_4086# 1.3e-22
C5048 a_2853_5648# a_3648_5972# 0.00271f
C5049 a_6011_4801# a_6010_3239# 1.39e-19
C5050 a_7247_4775# a_8237_4801# 0.00116f
C5051 a_2853_5648# a_2969_6040# 0.00149f
C5052 check[1] a_2883_5674# 0.195f
C5053 a_9578_4112# a_9638_3213# 4.45e-20
C5054 a_6760_4775# a_8403_4801# 1.55e-19
C5055 a_8402_3239# a_9151_3213# 0.139f
C5056 a_11970_4112# a_12101_2550# 1.72e-22
C5057 a_8236_3239# a_9638_3213# 0.0492f
C5058 a_8857_3213# a_8683_3605# 0.205f
C5059 a_4925_2550# a_5991_2340# 7.98e-21
C5060 x27.Q_N a_4585_3239# 4.03e-19
C5061 a_4453_2340# a_6546_2340# 6.38e-20
C5062 a_4657_2340# a_6304_2366# 1.32e-20
C5063 VDD a_1682_4775# 0.336f
C5064 x33.Q_N a_9464_3239# 0.00295f
C5065 a_11250_4775# a_11076_5167# 0.205f
C5066 a_10795_4801# a_11544_4775# 0.139f
C5067 a_10629_4801# a_12031_4775# 0.0492f
C5068 a_4155_4086# a_4019_4112# 0.0282f
C5069 a_4453_4386# a_4591_4478# 1.09e-19
C5070 a_3913_4112# a_4872_4394# 1.21e-20
C5071 a_4658_4086# x7.X 4.39e-21
C5072 a_8858_4775# a_9237_4386# 3.92e-19
C5073 a_8403_4801# a_9238_4086# 1.18e-19
C5074 a_8237_4801# a_9442_4086# 6.96e-19
C5075 a_9152_4775# a_8697_4112# 5.67e-20
C5076 a_8684_5167# a_8939_4086# 2.46e-20
C5077 a_6844_2640# a_7561_2732# 4.45e-20
C5078 a_6845_2340# a_7263_2648# 0.00276f
C5079 a_5561_3239# a_6010_3239# 6.84e-19
C5080 x75.Q a_5844_3239# 0.335f
C5081 a_6304_2366# D[4] 1.86e-20
C5082 sel_bit[1] a_2993_5674# 4.44e-19
C5083 a_8236_3239# a_9236_2640# 6.01e-20
C5084 a_4367_3213# a_3912_2366# 3.36e-20
C5085 a_3899_3605# a_4154_2340# 2.41e-20
C5086 a_4073_3213# a_4452_2640# 2.68e-19
C5087 check[0] x75.Q 0.0176f
C5088 a_8857_3213# a_8696_2366# 0.0014f
C5089 a_3618_3239# a_4453_2340# 6.38e-20
C5090 a_3452_3239# a_4657_2340# 4.77e-19
C5091 a_8683_3605# a_8383_2340# 3.9e-20
C5092 x33.Q_N a_9237_2340# 0.0469f
C5093 x4.X a_4872_4394# 8.47e-19
C5094 a_5992_4086# a_6547_4086# 0.197f
C5095 a_5372_4112# x45.Q_N 8.9e-20
C5096 x4.X a_4586_4801# 5.55e-19
C5097 VDD a_4453_2340# 0.788f
C5098 x5.X a_6199_4801# 0.00541f
C5099 x27.Q_N x45.Q_N 2.8e-20
C5100 x4.X a_11762_4801# 5.55e-19
C5101 a_7186_4112# a_6304_2366# 1.26e-20
C5102 a_6466_4775# a_6376_5167# 6.69e-20
C5103 a_6292_5167# a_6199_4801# 0.0367f
C5104 a_6760_4775# a_7073_4801# 0.124f
C5105 sel_bit[0] x48.Q_N 3.83e-20
C5106 a_6011_4801# a_4971_4801# 1.71e-20
C5107 D[4] a_8802_2366# 5.38e-19
C5108 a_8383_2340# a_8696_2366# 0.273f
C5109 check[3] D[2] 0.449f
C5110 a_11543_3213# a_11714_3521# 0.00652f
C5111 a_10794_3239# a_11183_3239# 0.0019f
C5112 a_11249_3213# a_11389_3239# 0.07f
C5113 a_10628_3239# a_11761_3239# 2.56e-19
C5114 x5.X x42.Q_N 0.00729f
C5115 VDD a_7763_2366# 0.109f
C5116 x4.X a_2061_2340# 0.00458f
C5117 VDD a_10794_3239# 0.274f
C5118 a_11629_4386# a_11565_4478# 2.13e-19
C5119 a_11630_4086# a_11289_4394# 1.25e-19
C5120 VDD a_9872_3521# 0.00506f
C5121 a_11089_4112# a_11195_4112# 0.051f
C5122 x30.Q_N a_6411_4112# 2.89e-22
C5123 a_11331_4086# a_11767_4478# 0.00412f
C5124 x27.D a_4318_5083# 3.45e-21
C5125 eob a_2788_5674# 1.71e-19
C5126 a_1207_2340# a_1720_2648# 0.00945f
C5127 x27.Q_N a_4452_2640# 0.569f
C5128 D[3] a_10680_2340# 0.0999f
C5129 check[3] a_11969_2366# 4.79e-19
C5130 a_11389_3239# a_10775_2340# 4.6e-20
C5131 a_2389_5648# a_2784_5996# 0.0102f
C5132 VDD a_6985_4112# 0.00445f
C5133 check[1] a_9237_2340# 1.98e-19
C5134 x4.X a_11089_4112# 0.109f
C5135 x5.X x7.X 6.95e-20
C5136 x4.X D[5] 5.17e-19
C5137 x4.X a_8857_3213# 0.00506f
C5138 a_9238_4086# a_9710_4296# 0.15f
C5139 a_9237_4386# x42.Q_N 0.00118f
C5140 check[2] x27.Q_N 3.57e-20
C5141 x4.X x72.Q_N 0.00455f
C5142 x7.X a_11856_3239# 1.89e-19
C5143 a_4681_4801# a_4971_4801# 0.0282f
C5144 a_4855_4775# a_4790_4801# 4.2e-20
C5145 a_4074_4775# a_4073_3213# 2.59e-19
C5146 a_3900_5167# a_3618_3239# 1.65e-21
C5147 x5.X a_11715_5083# 6.65e-19
C5148 a_3619_4801# a_3899_3605# 8.52e-21
C5149 a_4368_4775# a_3452_3239# 9.66e-21
C5150 check[2] x36.Q_N 0.0011f
C5151 check[5] a_7953_3239# 0.0271f
C5152 x20.Q_N a_4073_3213# 8.02e-21
C5153 a_8591_4801# a_8768_5167# 8.94e-19
C5154 a_8403_4801# a_8998_4801# 0.00118f
C5155 a_9152_4775# a_9102_5083# 1.21e-20
C5156 a_6759_3213# a_7246_3213# 0.273f
C5157 a_6465_3213# a_6198_3239# 6.99e-20
C5158 a_6010_3239# a_6375_3605# 4.45e-20
C5159 a_11390_4801# a_11543_3213# 1.61e-20
C5160 x36.Q_N a_10628_3239# 2.75e-19
C5161 a_11390_4801# a_11966_4801# 2.46e-21
C5162 VDD a_3900_5167# 0.324f
C5163 a_5088_3521# x75.Q_N 2.02e-20
C5164 a_6547_4086# a_6781_4478# 0.00976f
C5165 a_6305_4112# a_6983_4478# 0.00652f
C5166 a_5992_4086# a_6411_4112# 0.0397f
C5167 a_9237_4386# x7.X 2.49e-20
C5168 a_2463_4775# a_1511_4112# 0.0111f
C5169 x4.X a_8383_2340# 0.111f
C5170 VDD a_11076_5167# 0.317f
C5171 x7.X a_11629_2340# 0.183f
C5172 a_6011_4801# a_7954_4801# 8.38e-21
C5173 a_5845_4801# check[5] 8.72e-20
C5174 a_9755_4801# a_9710_4296# 1.9e-20
C5175 a_7953_3239# a_8402_3239# 3.93e-19
C5176 a_4925_2550# a_5371_2366# 0.0367f
C5177 D[0] a_8236_3239# 0.348f
C5178 a_6198_3239# a_5991_2340# 2.02e-19
C5179 a_7072_3239# a_6304_2366# 2.17e-19
C5180 check[1] a_4454_4086# 2.15e-20
C5181 a_6759_3213# a_6844_2640# 5.32e-19
C5182 a_6977_3239# D[0] 1.36e-20
C5183 a_10346_4801# a_10795_4801# 3.41e-19
C5184 check[4] a_10629_4801# 0.413f
C5185 check[0] x57.Q_N 0.0113f
C5186 a_1061_4801# a_2463_4775# 0.0492f
C5187 a_1682_4775# a_1508_5167# 0.205f
C5188 a_1227_4801# a_1976_4775# 0.132f
C5189 a_3600_4086# a_3913_4112# 0.273f
C5190 x4.X a_11766_2732# 9.81e-19
C5191 check[2] a_11629_4386# 1.44e-19
C5192 a_4681_4801# a_4214_4801# 0.00316f
C5193 check[2] a_9151_3213# 2.41e-20
C5194 x4.X a_5088_3521# 0.0012f
C5195 a_4368_4775# a_4586_4801# 3.73e-19
C5196 a_4074_4775# x27.Q_N 1.34e-19
C5197 check[5] a_8384_4086# 0.0042f
C5198 x20.Q_N x27.Q_N 1.21e-20
C5199 a_11089_4112# a_11249_3213# 0.00148f
C5200 a_11629_4386# a_10628_3239# 6.5e-20
C5201 a_11331_4086# a_10794_3239# 1.07e-20
C5202 a_9151_3213# a_10628_3239# 3.41e-19
C5203 a_6304_2366# a_6845_2340# 0.125f
C5204 a_6546_2340# a_6844_2640# 0.137f
C5205 a_4367_3213# a_6465_3213# 4.53e-20
C5206 a_4680_3239# a_5844_3239# 6.38e-20
C5207 a_4854_3213# a_6010_3239# 3.57e-19
C5208 a_9151_3213# a_9369_3239# 3.73e-19
C5209 a_9464_3239# a_8997_3239# 0.00316f
C5210 x4.X a_3600_4086# 0.106f
C5211 a_11250_4775# x36.Q_N 2.08e-20
C5212 a_11857_4801# a_11390_4801# 0.00316f
C5213 a_11544_4775# a_11762_4801# 3.73e-19
C5214 x4.X a_11767_4478# 0.00114f
C5215 a_4155_4086# x45.Q_N 1.43e-20
C5216 a_9238_4086# a_10681_4086# 2.08e-19
C5217 a_9710_4296# a_9954_4478# 0.00972f
C5218 a_8697_4112# a_9578_4112# 0.00943f
C5219 a_9442_4086# a_10156_4112# 6.99e-20
C5220 a_8939_4086# a_9377_4112# 0.00276f
C5221 VDD a_8768_5167# 0.0042f
C5222 VDD a_7246_3213# 0.569f
C5223 sel_bit[1] a_621_4112# 1.03e-20
C5224 check[6] a_7247_4775# 2.19e-20
C5225 a_8384_4086# a_8402_3239# 3.48e-19
C5226 a_8697_4112# a_8236_3239# 2.21e-19
C5227 x33.Q_N a_8939_4086# 1.3e-22
C5228 a_11089_4112# a_10775_2340# 5.05e-21
C5229 x20.Q_N a_2533_2550# 0.153f
C5230 a_7763_2366# a_8696_2366# 3.42e-20
C5231 a_1682_4775# x4.X 0.176f
C5232 a_9639_4775# check[4] 0.0122f
C5233 D[4] a_8383_2340# 0.0132f
C5234 a_4854_3213# a_4793_2366# 1.2e-20
C5235 eob a_2375_5167# 5.84e-19
C5236 x33.Q_N a_11628_2640# 1.12e-20
C5237 check[2] a_1976_4775# 0.00168f
C5238 a_2389_5648# a_2463_4775# 0.00225f
C5239 VDD a_6844_2640# 0.269f
C5240 check[0] a_4794_4112# 1.51e-19
C5241 a_3913_4112# a_4453_2340# 1.4e-21
C5242 a_4155_4086# a_4452_2640# 4.75e-21
C5243 a_10795_4801# a_11630_4086# 1.18e-19
C5244 x30.Q_N a_7561_2366# 0.00224f
C5245 a_11076_5167# a_11331_4086# 2.46e-20
C5246 x27.Q_N a_6759_3213# 8.29e-21
C5247 a_11250_4775# a_11629_4386# 3.92e-19
C5248 a_6199_4801# x30.Q_N 4.57e-21
C5249 a_10629_4801# a_11834_4086# 6.96e-19
C5250 a_11544_4775# a_11089_4112# 5.67e-20
C5251 a_2853_5648# x5.X 6.67e-19
C5252 a_9237_2340# a_10680_2340# 8.18e-19
C5253 a_8938_2340# a_9376_2366# 0.00276f
C5254 a_8696_2366# a_9577_2366# 0.00943f
C5255 a_3618_3239# a_4073_3213# 0.149f
C5256 a_11389_3239# a_11965_3239# 2.46e-21
C5257 a_3452_3239# a_3899_3605# 0.141f
C5258 x33.Q_N a_10983_4801# 1e-19
C5259 check[3] a_12101_2550# 9.97e-19
C5260 check[1] a_6466_4775# 5.74e-19
C5261 eob comparator_out 0.0519f
C5262 VDD a_9953_2732# 0.0042f
C5263 x4.X a_4453_2340# 0.00242f
C5264 VDD a_7159_5167# 0.00371f
C5265 check[2] a_12048_4394# 1.36e-20
C5266 VDD a_12146_3239# 4.88e-19
C5267 VDD a_4073_3213# 0.314f
C5268 x45.Q_N a_7953_3239# 3.23e-19
C5269 VDD a_11761_3239# 6.2e-19
C5270 x30.Q_N x42.Q_N 1.63e-20
C5271 a_11195_4112# a_10794_3239# 4.04e-21
C5272 a_1626_2366# a_1996_2366# 4.11e-20
C5273 x27.Q_N a_6546_2340# 5.08e-20
C5274 check[5] a_7182_4801# 1.11e-20
C5275 a_11088_2366# a_11564_2732# 0.00133f
C5276 check[1] a_8939_4086# 3.29e-19
C5277 x5.X a_6846_4086# 0.261f
C5278 x4.X a_7763_2366# 8.68e-20
C5279 a_12345_2366# VSS 8.87e-19
C5280 a_11969_2366# VSS 0.182f
C5281 a_11768_2366# VSS 0.00989f
C5282 a_11564_2366# VSS 0.00207f
C5283 a_12547_2366# VSS 0.0962f
C5284 a_12345_2732# VSS 3.33e-19
C5285 a_12047_2648# VSS 4.04e-19
C5286 a_11194_2366# VSS 0.158f
C5287 a_11766_2732# VSS 0.0011f
C5288 a_11564_2732# VSS 1.58e-19
C5289 a_11288_2648# VSS 1.45e-19
C5290 a_9953_2366# VSS 6.96e-19
C5291 x63.Q_N VSS 0.1f
C5292 a_12101_2550# VSS 0.262f
C5293 a_11833_2340# VSS 0.29f
C5294 a_11629_2340# VSS 0.606f
C5295 a_11628_2640# VSS 0.419f
C5296 a_11330_2340# VSS 0.251f
C5297 a_11088_2366# VSS 0.387f
C5298 a_10775_2340# VSS 0.458f
C5299 a_9577_2366# VSS 0.18f
C5300 a_9376_2366# VSS 0.00923f
C5301 a_9172_2366# VSS 0.00192f
C5302 a_10680_2340# VSS 0.225f
C5303 D[3] VSS 0.365f
C5304 a_10155_2366# VSS 0.0926f
C5305 a_8802_2366# VSS 0.157f
C5306 a_9374_2732# VSS 3.84e-19
C5307 a_7561_2366# VSS 6.96e-19
C5308 x60.Q_N VSS 0.1f
C5309 a_9709_2550# VSS 0.256f
C5310 a_9441_2340# VSS 0.286f
C5311 a_9237_2340# VSS 0.512f
C5312 a_9236_2640# VSS 0.4f
C5313 a_8938_2340# VSS 0.249f
C5314 a_8696_2366# VSS 0.385f
C5315 a_8383_2340# VSS 0.456f
C5316 a_7185_2366# VSS 0.18f
C5317 a_6984_2366# VSS 0.00923f
C5318 a_6780_2366# VSS 0.00192f
C5319 a_8288_2340# VSS 0.225f
C5320 D[4] VSS 0.365f
C5321 a_7763_2366# VSS 0.0926f
C5322 a_6410_2366# VSS 0.157f
C5323 a_6982_2732# VSS 3.84e-19
C5324 a_5169_2366# VSS 6.96e-19
C5325 x57.Q_N VSS 0.1f
C5326 a_7317_2550# VSS 0.256f
C5327 a_7049_2340# VSS 0.286f
C5328 a_6845_2340# VSS 0.513f
C5329 a_6844_2640# VSS 0.4f
C5330 a_6546_2340# VSS 0.249f
C5331 a_6304_2366# VSS 0.385f
C5332 a_5991_2340# VSS 0.456f
C5333 a_4793_2366# VSS 0.18f
C5334 a_4592_2366# VSS 0.00923f
C5335 a_4388_2366# VSS 0.00192f
C5336 a_5896_2340# VSS 0.225f
C5337 D[5] VSS 0.393f
C5338 a_5371_2366# VSS 0.0926f
C5339 a_4018_2366# VSS 0.157f
C5340 a_4590_2732# VSS 3.84e-19
C5341 a_2777_2366# VSS 0.00168f
C5342 x54.Q_N VSS 0.1f
C5343 a_4925_2550# VSS 0.256f
C5344 a_4657_2340# VSS 0.286f
C5345 a_4453_2340# VSS 0.513f
C5346 a_4452_2640# VSS 0.4f
C5347 a_4154_2340# VSS 0.249f
C5348 a_3912_2366# VSS 0.385f
C5349 a_3599_2340# VSS 0.458f
C5350 a_2401_2366# VSS 0.18f
C5351 a_2200_2366# VSS 0.00923f
C5352 a_1996_2366# VSS 0.00192f
C5353 a_3504_2340# VSS 0.226f
C5354 D[6] VSS 0.604f
C5355 a_2979_2366# VSS 0.0988f
C5356 a_1626_2366# VSS 0.157f
C5357 a_2198_2732# VSS 3.84e-19
C5358 x51.Q_N VSS 0.1f
C5359 a_2533_2550# VSS 0.263f
C5360 a_2265_2340# VSS 0.289f
C5361 a_2061_2340# VSS 0.517f
C5362 a_2060_2640# VSS 0.527f
C5363 a_1762_2340# VSS 0.25f
C5364 a_1520_2366# VSS 0.387f
C5365 a_1207_2340# VSS 0.466f
C5366 D[7] VSS 0.535f
C5367 a_1112_2340# VSS 0.246f
C5368 a_11965_3239# VSS 0.00208f
C5369 a_12146_3239# VSS 0.159f
C5370 D[2] VSS 1.11f
C5371 a_12737_3239# VSS 0.252f
C5372 x66.Q_N VSS 0.102f
C5373 a_12264_3521# VSS 3.9e-19
C5374 a_11761_3239# VSS 0.00967f
C5375 a_11183_3239# VSS 0.00168f
C5376 a_11389_3239# VSS 0.181f
C5377 a_11942_3605# VSS 2.25e-19
C5378 a_11714_3521# VSS 0.00103f
C5379 a_11493_3521# VSS 2.34e-19
C5380 a_9573_3239# VSS 0.00192f
C5381 a_9754_3239# VSS 0.157f
C5382 a_10982_3239# VSS 0.0988f
C5383 a_11856_3239# VSS 0.25f
C5384 a_12030_3213# VSS 0.463f
C5385 a_11543_3213# VSS 0.389f
C5386 a_11075_3605# VSS 0.259f
C5387 a_11249_3213# VSS 0.281f
C5388 a_10794_3239# VSS 0.519f
C5389 a_10628_3239# VSS 0.509f
C5390 D[1] VSS 0.467f
C5391 a_10345_3239# VSS 0.222f
C5392 x69.Q_N VSS 0.1f
C5393 a_9369_3239# VSS 0.00923f
C5394 a_8791_3239# VSS 0.00168f
C5395 a_8997_3239# VSS 0.18f
C5396 a_9322_3521# VSS 3.84e-19
C5397 a_7181_3239# VSS 0.00192f
C5398 a_7362_3239# VSS 0.157f
C5399 a_8590_3239# VSS 0.0988f
C5400 a_9464_3239# VSS 0.246f
C5401 a_9638_3213# VSS 0.446f
C5402 a_9151_3213# VSS 0.38f
C5403 a_8683_3605# VSS 0.258f
C5404 a_8857_3213# VSS 0.28f
C5405 a_8402_3239# VSS 0.519f
C5406 a_8236_3239# VSS 0.506f
C5407 D[0] VSS 0.471f
C5408 a_7953_3239# VSS 0.222f
C5409 x72.Q_N VSS 0.1f
C5410 a_6977_3239# VSS 0.00923f
C5411 a_6399_3239# VSS 0.00168f
C5412 a_6605_3239# VSS 0.18f
C5413 a_6930_3521# VSS 3.84e-19
C5414 a_4789_3239# VSS 0.00196f
C5415 a_4970_3239# VSS 0.157f
C5416 a_6198_3239# VSS 0.0988f
C5417 a_7072_3239# VSS 0.246f
C5418 a_7246_3213# VSS 0.446f
C5419 a_6759_3213# VSS 0.38f
C5420 a_6291_3605# VSS 0.258f
C5421 a_6465_3213# VSS 0.28f
C5422 a_6010_3239# VSS 0.519f
C5423 a_5844_3239# VSS 0.506f
C5424 x75.Q VSS 0.239f
C5425 a_5561_3239# VSS 0.222f
C5426 x75.Q_N VSS 0.1f
C5427 a_4585_3239# VSS 0.00943f
C5428 a_4007_3239# VSS 0.00202f
C5429 a_4213_3239# VSS 0.181f
C5430 a_4538_3521# VSS 3.84e-19
C5431 a_3806_3239# VSS 0.263f
C5432 a_4680_3239# VSS 0.246f
C5433 a_4854_3213# VSS 0.446f
C5434 a_4367_3213# VSS 0.379f
C5435 a_3899_3605# VSS 0.261f
C5436 a_4073_3213# VSS 0.28f
C5437 a_3618_3239# VSS 0.751f
C5438 a_3452_3239# VSS 0.888f
C5439 x77.Y VSS 1.02f
C5440 x7.X VSS 11.5f
C5441 a_929_3238# VSS 0.532f
C5442 x7.A VSS 0.204f
C5443 a_653_3238# VSS 0.285f
C5444 comparator_out VSS 0.577f
C5445 a_12346_4112# VSS 0.00226f
C5446 a_11970_4112# VSS 0.183f
C5447 a_11769_4112# VSS 0.00991f
C5448 a_11565_4112# VSS 0.00168f
C5449 a_12548_4112# VSS 0.102f
C5450 a_12346_4478# VSS 3.33e-19
C5451 a_12048_4394# VSS 3.91e-19
C5452 a_11195_4112# VSS 0.148f
C5453 a_11767_4478# VSS 0.00107f
C5454 a_11565_4478# VSS 1.58e-19
C5455 a_11289_4394# VSS 1.48e-19
C5456 a_9954_4112# VSS 0.00168f
C5457 x39.Q_N VSS 1.23f
C5458 a_12102_4296# VSS 0.261f
C5459 a_11834_4086# VSS 0.279f
C5460 a_11630_4086# VSS 0.588f
C5461 a_11629_4386# VSS 0.537f
C5462 a_11331_4086# VSS 0.238f
C5463 a_11089_4112# VSS 0.318f
C5464 a_10776_4086# VSS 0.425f
C5465 a_9578_4112# VSS 0.18f
C5466 a_9377_4112# VSS 0.00923f
C5467 a_9173_4112# VSS 0.00155f
C5468 a_10681_4086# VSS 0.207f
C5469 a_10156_4112# VSS 0.0984f
C5470 a_8803_4112# VSS 0.147f
C5471 a_9375_4478# VSS 3.84e-19
C5472 a_7562_4112# VSS 0.00168f
C5473 x42.Q_N VSS 1.22f
C5474 a_9710_4296# VSS 0.255f
C5475 a_9442_4086# VSS 0.275f
C5476 a_9238_4086# VSS 0.484f
C5477 a_9237_4386# VSS 0.515f
C5478 a_8939_4086# VSS 0.236f
C5479 a_8697_4112# VSS 0.316f
C5480 a_8384_4086# VSS 0.423f
C5481 a_7186_4112# VSS 0.18f
C5482 a_6985_4112# VSS 0.00923f
C5483 a_6781_4112# VSS 0.00157f
C5484 a_8289_4086# VSS 0.205f
C5485 a_7764_4112# VSS 0.0984f
C5486 a_6411_4112# VSS 0.147f
C5487 a_6983_4478# VSS 3.84e-19
C5488 a_5170_4112# VSS 0.00168f
C5489 x45.Q_N VSS 1.22f
C5490 a_7318_4296# VSS 0.255f
C5491 a_7050_4086# VSS 0.275f
C5492 a_6846_4086# VSS 0.484f
C5493 a_6845_4386# VSS 0.515f
C5494 a_6547_4086# VSS 0.236f
C5495 a_6305_4112# VSS 0.316f
C5496 a_5992_4086# VSS 0.423f
C5497 a_4794_4112# VSS 0.18f
C5498 a_4593_4112# VSS 0.00923f
C5499 a_4389_4112# VSS 0.00192f
C5500 a_5897_4086# VSS 0.211f
C5501 a_5372_4112# VSS 0.0984f
C5502 a_4019_4112# VSS 0.157f
C5503 a_4591_4478# VSS 3.84e-19
C5504 x48.Q_N VSS 0.1f
C5505 a_4926_4296# VSS 0.255f
C5506 a_4658_4086# VSS 0.275f
C5507 a_4454_4086# VSS 0.486f
C5508 a_4453_4386# VSS 0.515f
C5509 a_4155_4086# VSS 0.243f
C5510 a_3913_4112# VSS 0.373f
C5511 a_3600_4086# VSS 0.443f
C5512 a_3505_4086# VSS 0.225f
C5513 a_1511_4112# VSS 2.05f
C5514 x4.A VSS 0.931f
C5515 a_897_4112# VSS 0.511f
C5516 x3.A VSS 0.203f
C5517 a_621_4112# VSS 0.282f
C5518 reset VSS 0.244f
C5519 a_11966_4801# VSS 0.00215f
C5520 a_12147_4801# VSS 0.161f
C5521 check[3] VSS 1.3f
C5522 a_12738_4801# VSS 0.255f
C5523 x36.Q_N VSS 1.28f
C5524 a_12265_5083# VSS 5.88e-19
C5525 a_11762_4801# VSS 0.00989f
C5526 a_11184_4801# VSS 0.00168f
C5527 a_11390_4801# VSS 0.181f
C5528 a_11943_5167# VSS 2.29e-19
C5529 a_11715_5083# VSS 0.00114f
C5530 a_11494_5083# VSS 2.58e-19
C5531 a_9574_4801# VSS 0.00192f
C5532 a_9755_4801# VSS 0.157f
C5533 a_10983_4801# VSS 0.0987f
C5534 a_11857_4801# VSS 0.25f
C5535 a_12031_4775# VSS 0.46f
C5536 a_11544_4775# VSS 0.386f
C5537 a_11076_5167# VSS 0.257f
C5538 a_11250_4775# VSS 0.279f
C5539 a_10795_4801# VSS 0.517f
C5540 a_10629_4801# VSS 0.488f
C5541 check[4] VSS 0.823f
C5542 a_10346_4801# VSS 0.21f
C5543 x33.Q_N VSS 1.25f
C5544 a_9370_4801# VSS 0.00923f
C5545 a_8792_4801# VSS 0.00168f
C5546 a_8998_4801# VSS 0.18f
C5547 a_9323_5083# VSS 3.84e-19
C5548 a_7182_4801# VSS 0.00192f
C5549 a_7363_4801# VSS 0.157f
C5550 a_8591_4801# VSS 0.0987f
C5551 a_9465_4801# VSS 0.244f
C5552 a_9639_4775# VSS 0.435f
C5553 a_9152_4775# VSS 0.373f
C5554 a_8684_5167# VSS 0.257f
C5555 a_8858_4775# VSS 0.276f
C5556 a_8403_4801# VSS 0.515f
C5557 a_8237_4801# VSS 0.484f
C5558 check[5] VSS 0.83f
C5559 a_7954_4801# VSS 0.207f
C5560 x30.Q_N VSS 1.26f
C5561 a_6978_4801# VSS 0.00923f
C5562 a_6400_4801# VSS 0.00168f
C5563 a_6606_4801# VSS 0.18f
C5564 a_6931_5083# VSS 3.84e-19
C5565 a_4790_4801# VSS 0.00192f
C5566 a_4971_4801# VSS 0.157f
C5567 a_6199_4801# VSS 0.0987f
C5568 a_7073_4801# VSS 0.244f
C5569 a_7247_4775# VSS 0.435f
C5570 a_6760_4775# VSS 0.373f
C5571 a_6292_5167# VSS 0.257f
C5572 a_6466_4775# VSS 0.276f
C5573 a_6011_4801# VSS 0.515f
C5574 a_5845_4801# VSS 0.484f
C5575 check[6] VSS 0.845f
C5576 a_5562_4801# VSS 0.207f
C5577 x27.Q_N VSS 1.25f
C5578 a_4586_4801# VSS 0.00923f
C5579 a_4008_4801# VSS 0.00168f
C5580 a_4214_4801# VSS 0.18f
C5581 a_4539_5083# VSS 3.84e-19
C5582 a_2398_4801# VSS 0.00192f
C5583 a_2579_4801# VSS 0.157f
C5584 a_3807_4801# VSS 0.0987f
C5585 a_4681_4801# VSS 0.244f
C5586 a_4855_4775# VSS 0.435f
C5587 a_4368_4775# VSS 0.373f
C5588 a_3900_5167# VSS 0.257f
C5589 a_4074_4775# VSS 0.275f
C5590 a_3619_4801# VSS 0.513f
C5591 a_3453_4801# VSS 0.481f
C5592 x27.D VSS 0.243f
C5593 a_3170_4801# VSS 0.22f
C5594 x20.Q_N VSS 1.24f
C5595 a_2194_4801# VSS 0.00923f
C5596 a_1616_4801# VSS 0.00168f
C5597 a_1822_4801# VSS 0.18f
C5598 a_2147_5083# VSS 3.84e-19
C5599 a_1415_4801# VSS 0.0987f
C5600 a_2289_4801# VSS 0.242f
C5601 a_2463_4775# VSS 0.429f
C5602 a_1976_4775# VSS 0.37f
C5603 a_1508_5167# VSS 0.256f
C5604 x4.X VSS 16.5f
C5605 a_1682_4775# VSS 0.274f
C5606 a_1227_4801# VSS 0.516f
C5607 a_1061_4801# VSS 0.54f
C5608 a_3877_5674# VSS 0.00437f
C5609 a_3671_5674# VSS 0.00563f
C5610 a_2993_5674# VSS 0.00182f
C5611 a_2788_5674# VSS 0.00372f
C5612 a_3373_5674# VSS 0.115f
C5613 a_3258_5648# VSS 0.229f
C5614 check[0] VSS 2.45f
C5615 x48.Q VSS 0.615f
C5616 sel_bit[1] VSS 1.15f
C5617 a_2883_5674# VSS 0.185f
C5618 a_2784_5996# VSS 2.03e-19
C5619 eob VSS 2.51f
C5620 x5.X VSS 13f
C5621 check[1] VSS 2.75f
C5622 a_2853_5648# VSS 0.373f
C5623 sel_bit[0] VSS 0.539f
C5624 check[2] VSS 4.55f
C5625 a_2389_5648# VSS 0.479f
C5626 a_1338_5674# VSS 0.514f
C5627 x5.A VSS 0.197f
C5628 a_1062_5674# VSS 0.276f
C5629 clk_sar VSS 0.214f
C5630 VDD VSS 0.107p
C5631 check[2].t0 VSS 0.0384f
C5632 check[2].n0 VSS 0.00289f
C5633 check[2].t3 VSS 0.0197f
C5634 check[2].t2 VSS 0.0123f
C5635 check[2].n1 VSS 0.0406f
C5636 check[2].n2 VSS 0.629f
C5637 check[2].t5 VSS 0.0179f
C5638 check[2].t4 VSS 0.0125f
C5639 check[2].n3 VSS 0.0364f
C5640 check[2].n4 VSS 0.0138f
C5641 check[2].n5 VSS 0.836f
C5642 check[2].n6 VSS 0.0257f
C5643 check[2].n7 VSS 0.198f
C5644 check[2].t1 VSS 0.0144f
C5645 check[2].n8 VSS 0.0246f
C5646 x4.X.n0 VSS 0.00768f
C5647 x4.X.n1 VSS 0.00767f
C5648 x4.X.n2 VSS 0.00768f
C5649 x4.X.n3 VSS 0.00767f
C5650 x4.X.n4 VSS 0.00768f
C5651 x4.X.n5 VSS 0.00779f
C5652 x4.X.n6 VSS 0.0356f
C5653 x4.X.n7 VSS 0.00746f
C5654 x4.X.n8 VSS 0.00423f
C5655 x4.X.n9 VSS 0.00216f
C5656 x4.X.n10 VSS 0.00427f
C5657 x4.X.n11 VSS 0.0017f
C5658 x4.X.n12 VSS 0.00446f
C5659 x4.X.t4 VSS 0.00963f
C5660 x4.X.t10 VSS 0.00963f
C5661 x4.X.n13 VSS 0.0238f
C5662 x4.X.t3 VSS 0.00963f
C5663 x4.X.t14 VSS 0.00963f
C5664 x4.X.n14 VSS 0.0238f
C5665 x4.X.t11 VSS 0.00963f
C5666 x4.X.t2 VSS 0.00963f
C5667 x4.X.n15 VSS 0.0238f
C5668 x4.X.t7 VSS 0.00963f
C5669 x4.X.t0 VSS 0.00963f
C5670 x4.X.n16 VSS 0.0238f
C5671 x4.X.t6 VSS 0.00963f
C5672 x4.X.t1 VSS 0.00963f
C5673 x4.X.n17 VSS 0.0368f
C5674 x4.X.t8 VSS 0.00963f
C5675 x4.X.t12 VSS 0.00963f
C5676 x4.X.n18 VSS 0.0238f
C5677 x4.X.n19 VSS 0.0926f
C5678 x4.X.t9 VSS 0.00963f
C5679 x4.X.t13 VSS 0.00963f
C5680 x4.X.n20 VSS 0.0238f
C5681 x4.X.n21 VSS 0.0559f
C5682 x4.X.n22 VSS 0.00913f
C5683 x4.X.t5 VSS 0.00821f
C5684 x4.X.n23 VSS 0.00963f
C5685 x4.X.t66 VSS 0.0152f
C5686 x4.X.t32 VSS 0.00645f
C5687 x4.X.n24 VSS 0.0286f
C5688 x4.X.n25 VSS 0.00238f
C5689 x4.X.n26 VSS 0.0084f
C5690 x4.X.n27 VSS 0.0033f
C5691 x4.X.n28 VSS 0.0389f
C5692 x4.X.n29 VSS 0.103f
C5693 x4.X.n30 VSS 0.00153f
C5694 x4.X.t50 VSS 0.0152f
C5695 x4.X.t37 VSS 0.00644f
C5696 x4.X.n31 VSS 0.0297f
C5697 x4.X.n32 VSS 0.00977f
C5698 x4.X.n33 VSS 0.00208f
C5699 x4.X.n34 VSS 0.0273f
C5700 x4.X.n35 VSS 0.00586f
C5701 x4.X.n36 VSS 0.00803f
C5702 x4.X.n37 VSS 0.0201f
C5703 x4.X.t15 VSS 0.005f
C5704 x4.X.n38 VSS 0.00963f
C5705 x4.X.n39 VSS 0.00651f
C5706 x4.X.n40 VSS 0.00614f
C5707 x4.X.n41 VSS 0.0246f
C5708 x4.X.n42 VSS 0.0559f
C5709 x4.X.n43 VSS 0.0559f
C5710 x4.X.n44 VSS 0.0559f
C5711 x4.X.n45 VSS 0.0532f
C5712 x4.X.t18 VSS 0.00626f
C5713 x4.X.t29 VSS 0.00626f
C5714 x4.X.n46 VSS 0.0297f
C5715 x4.X.t20 VSS 0.00626f
C5716 x4.X.t24 VSS 0.00626f
C5717 x4.X.n47 VSS 0.0157f
C5718 x4.X.n48 VSS 0.0587f
C5719 x4.X.t21 VSS 0.00626f
C5720 x4.X.t25 VSS 0.00626f
C5721 x4.X.n49 VSS 0.0157f
C5722 x4.X.n50 VSS 0.0395f
C5723 x4.X.t17 VSS 0.00626f
C5724 x4.X.t27 VSS 0.00626f
C5725 x4.X.n51 VSS 0.0157f
C5726 x4.X.n52 VSS 0.0396f
C5727 x4.X.t19 VSS 0.00626f
C5728 x4.X.t28 VSS 0.00626f
C5729 x4.X.n53 VSS 0.0157f
C5730 x4.X.n54 VSS 0.0396f
C5731 x4.X.t23 VSS 0.00626f
C5732 x4.X.t30 VSS 0.00626f
C5733 x4.X.n55 VSS 0.0157f
C5734 x4.X.n56 VSS 0.0396f
C5735 x4.X.t31 VSS 0.00626f
C5736 x4.X.t26 VSS 0.00626f
C5737 x4.X.n57 VSS 0.0157f
C5738 x4.X.n58 VSS 0.0396f
C5739 x4.X.t16 VSS 0.00626f
C5740 x4.X.t22 VSS 0.00626f
C5741 x4.X.n59 VSS 0.0157f
C5742 x4.X.n60 VSS 0.0384f
C5743 x4.X.n61 VSS 0.00482f
C5744 x4.X.t58 VSS 0.009f
C5745 x4.X.t45 VSS 0.0104f
C5746 x4.X.n62 VSS 0.0242f
C5747 x4.X.n63 VSS 0.00675f
C5748 x4.X.n64 VSS 0.00238f
C5749 x4.X.n65 VSS 0.0014f
C5750 x4.X.n66 VSS 0.0083f
C5751 x4.X.n67 VSS 0.0546f
C5752 x4.X.n68 VSS 0.00482f
C5753 x4.X.t55 VSS 0.009f
C5754 x4.X.t51 VSS 0.0104f
C5755 x4.X.n69 VSS 0.0242f
C5756 x4.X.n70 VSS 0.00675f
C5757 x4.X.n71 VSS 0.00238f
C5758 x4.X.n72 VSS 0.0014f
C5759 x4.X.n73 VSS 0.00821f
C5760 x4.X.n74 VSS 0.0259f
C5761 x4.X.n75 VSS 0.113f
C5762 x4.X.n76 VSS 0.00271f
C5763 x4.X.n77 VSS 0.0014f
C5764 x4.X.t34 VSS 0.0103f
C5765 x4.X.t39 VSS 0.00868f
C5766 x4.X.n78 VSS 0.0115f
C5767 x4.X.n79 VSS 0.0128f
C5768 x4.X.n80 VSS 0.0189f
C5769 x4.X.n81 VSS 0.00271f
C5770 x4.X.n82 VSS 0.0014f
C5771 x4.X.t54 VSS 0.0103f
C5772 x4.X.t60 VSS 0.0087f
C5773 x4.X.n83 VSS 0.0117f
C5774 x4.X.n84 VSS 0.0126f
C5775 x4.X.n85 VSS 0.0588f
C5776 x4.X.n86 VSS 0.16f
C5777 x4.X.n87 VSS 0.135f
C5778 x4.X.n88 VSS 0.00482f
C5779 x4.X.t36 VSS 0.00905f
C5780 x4.X.t57 VSS 0.0103f
C5781 x4.X.n89 VSS 0.0242f
C5782 x4.X.n90 VSS 0.00661f
C5783 x4.X.n91 VSS 0.00246f
C5784 x4.X.n92 VSS 0.0014f
C5785 x4.X.n93 VSS 0.0083f
C5786 x4.X.n94 VSS 0.0547f
C5787 x4.X.n95 VSS 0.00482f
C5788 x4.X.t33 VSS 0.009f
C5789 x4.X.t63 VSS 0.0104f
C5790 x4.X.n96 VSS 0.0242f
C5791 x4.X.n97 VSS 0.00675f
C5792 x4.X.n98 VSS 0.00238f
C5793 x4.X.n99 VSS 0.0014f
C5794 x4.X.n100 VSS 0.00821f
C5795 x4.X.n101 VSS 0.0259f
C5796 x4.X.n102 VSS 0.0847f
C5797 x4.X.n103 VSS 0.125f
C5798 x4.X.n104 VSS 0.00271f
C5799 x4.X.n105 VSS 0.0014f
C5800 x4.X.t69 VSS 0.0103f
C5801 x4.X.t49 VSS 0.0087f
C5802 x4.X.n106 VSS 0.0117f
C5803 x4.X.n107 VSS 0.0126f
C5804 x4.X.n108 VSS 0.0199f
C5805 x4.X.n109 VSS 0.00271f
C5806 x4.X.n110 VSS 0.0014f
C5807 x4.X.t52 VSS 0.0103f
C5808 x4.X.t67 VSS 0.0087f
C5809 x4.X.n111 VSS 0.0117f
C5810 x4.X.n112 VSS 0.0126f
C5811 x4.X.n113 VSS 0.0589f
C5812 x4.X.n114 VSS 0.16f
C5813 x4.X.n115 VSS 0.126f
C5814 x4.X.n116 VSS 0.0047f
C5815 x4.X.t42 VSS 0.009f
C5816 x4.X.t64 VSS 0.0104f
C5817 x4.X.n117 VSS 0.0242f
C5818 x4.X.n118 VSS 0.00653f
C5819 x4.X.n119 VSS 0.00254f
C5820 x4.X.n120 VSS 0.0014f
C5821 x4.X.n121 VSS 0.0083f
C5822 x4.X.n122 VSS 0.0546f
C5823 x4.X.n123 VSS 0.00482f
C5824 x4.X.t41 VSS 0.00909f
C5825 x4.X.t38 VSS 0.0103f
C5826 x4.X.n124 VSS 0.0242f
C5827 x4.X.n125 VSS 0.00661f
C5828 x4.X.n126 VSS 0.00246f
C5829 x4.X.n127 VSS 0.0014f
C5830 x4.X.n128 VSS 0.00821f
C5831 x4.X.n129 VSS 0.0257f
C5832 x4.X.n130 VSS 0.0844f
C5833 x4.X.n131 VSS 0.125f
C5834 x4.X.n132 VSS 0.00271f
C5835 x4.X.n133 VSS 0.0014f
C5836 x4.X.t46 VSS 0.0103f
C5837 x4.X.t61 VSS 0.0087f
C5838 x4.X.n134 VSS 0.0117f
C5839 x4.X.n135 VSS 0.0126f
C5840 x4.X.n136 VSS 0.019f
C5841 x4.X.n137 VSS 0.00271f
C5842 x4.X.n138 VSS 0.0014f
C5843 x4.X.t65 VSS 0.0103f
C5844 x4.X.t43 VSS 0.00868f
C5845 x4.X.n139 VSS 0.0115f
C5846 x4.X.n140 VSS 0.0128f
C5847 x4.X.n141 VSS 0.0589f
C5848 x4.X.n142 VSS 0.161f
C5849 x4.X.n143 VSS 0.125f
C5850 x4.X.t56 VSS 0.009f
C5851 x4.X.t35 VSS 0.0104f
C5852 x4.X.n144 VSS 0.0242f
C5853 x4.X.n145 VSS 0.00631f
C5854 x4.X.n146 VSS 0.00271f
C5855 x4.X.n147 VSS 0.00141f
C5856 x4.X.n148 VSS 0.00518f
C5857 x4.X.n149 VSS 0.00686f
C5858 x4.X.n150 VSS 0.00893f
C5859 x4.X.n151 VSS 0.0541f
C5860 x4.X.t40 VSS 0.0105f
C5861 x4.X.t53 VSS 0.00892f
C5862 x4.X.n152 VSS 0.0242f
C5863 x4.X.n153 VSS 0.00639f
C5864 x4.X.n154 VSS 0.00263f
C5865 x4.X.n155 VSS 0.0014f
C5866 x4.X.n156 VSS 0.00482f
C5867 x4.X.n157 VSS 0.00769f
C5868 x4.X.n158 VSS 0.00848f
C5869 x4.X.n159 VSS 0.0259f
C5870 x4.X.n160 VSS 0.0851f
C5871 x4.X.n161 VSS 0.125f
C5872 x4.X.n162 VSS 0.00271f
C5873 x4.X.n163 VSS 0.0014f
C5874 x4.X.t48 VSS 0.0103f
C5875 x4.X.t62 VSS 0.00868f
C5876 x4.X.n164 VSS 0.0115f
C5877 x4.X.n165 VSS 0.0128f
C5878 x4.X.n166 VSS 0.0221f
C5879 x4.X.n167 VSS 0.00778f
C5880 x4.X.n168 VSS 0.0061f
C5881 x4.X.n169 VSS 0.00271f
C5882 x4.X.t47 VSS 0.009f
C5883 x4.X.t68 VSS 0.0103f
C5884 x4.X.n170 VSS 0.0128f
C5885 x4.X.n171 VSS 0.0112f
C5886 x4.X.n172 VSS 0.00148f
C5887 x4.X.n173 VSS 0.00507f
C5888 x4.X.n174 VSS 0.00813f
C5889 x4.X.n175 VSS 0.0698f
C5890 x4.X.n176 VSS 0.119f
C5891 x4.X.n177 VSS 0.103f
C5892 x4.X.t44 VSS 0.0104f
C5893 x4.X.t59 VSS 0.00899f
C5894 x4.X.n178 VSS 0.0239f
C5895 x4.X.n179 VSS 0.168f
C5896 x4.X.n180 VSS 0.304f
C5897 x4.X.n181 VSS 0.0328f
C5898 x5.X.n0 VSS 0.0705f
C5899 x5.X.n1 VSS 0.0499f
C5900 x5.X.n2 VSS 0.05f
C5901 x5.X.t24 VSS 0.0128f
C5902 x5.X.t11 VSS 0.00992f
C5903 x5.X.n3 VSS 0.0251f
C5904 x5.X.n4 VSS 0.00749f
C5905 x5.X.n5 VSS 0.00463f
C5906 x5.X.n6 VSS 0.00187f
C5907 x5.X.t15 VSS 0.0125f
C5908 x5.X.n7 VSS 0.0129f
C5909 x5.X.n8 VSS 0.00145f
C5910 x5.X.t20 VSS 0.00945f
C5911 x5.X.n9 VSS 0.0114f
C5912 x5.X.n10 VSS 0.00259f
C5913 x5.X.n11 VSS 0.00389f
C5914 x5.X.n12 VSS 0.00462f
C5915 x5.X.n13 VSS 0.00187f
C5916 x5.X.t13 VSS 0.0126f
C5917 x5.X.n14 VSS 0.013f
C5918 x5.X.n15 VSS 0.00145f
C5919 x5.X.t18 VSS 0.00933f
C5920 x5.X.n16 VSS 0.0113f
C5921 x5.X.n17 VSS 0.00287f
C5922 x5.X.n18 VSS 0.0495f
C5923 x5.X.n19 VSS 0.0664f
C5924 x5.X.n20 VSS 0.013f
C5925 x5.X.n21 VSS 0.0394f
C5926 x5.X.n22 VSS 0.322f
C5927 x5.X.n23 VSS 0.00462f
C5928 x5.X.n24 VSS 0.00187f
C5929 x5.X.t21 VSS 0.0126f
C5930 x5.X.n25 VSS 0.0129f
C5931 x5.X.n26 VSS 0.00145f
C5932 x5.X.t8 VSS 0.00941f
C5933 x5.X.n27 VSS 0.0114f
C5934 x5.X.n28 VSS 0.00272f
C5935 x5.X.n29 VSS 0.00537f
C5936 x5.X.n30 VSS 0.00462f
C5937 x5.X.n31 VSS 0.00187f
C5938 x5.X.t17 VSS 0.0126f
C5939 x5.X.n32 VSS 0.013f
C5940 x5.X.n33 VSS 0.00145f
C5941 x5.X.t25 VSS 0.00933f
C5942 x5.X.n34 VSS 0.0113f
C5943 x5.X.n35 VSS 0.00287f
C5944 x5.X.n36 VSS 0.0487f
C5945 x5.X.n37 VSS 0.0657f
C5946 x5.X.n38 VSS 0.228f
C5947 x5.X.n39 VSS 0.00462f
C5948 x5.X.n40 VSS 0.00187f
C5949 x5.X.t22 VSS 0.0126f
C5950 x5.X.n41 VSS 0.0129f
C5951 x5.X.n42 VSS 0.00145f
C5952 x5.X.t9 VSS 0.00941f
C5953 x5.X.n43 VSS 0.0114f
C5954 x5.X.n44 VSS 0.00265f
C5955 x5.X.n45 VSS 0.00551f
C5956 x5.X.n46 VSS 0.00462f
C5957 x5.X.n47 VSS 0.00187f
C5958 x5.X.t14 VSS 0.0126f
C5959 x5.X.n48 VSS 0.013f
C5960 x5.X.n49 VSS 0.00145f
C5961 x5.X.t19 VSS 0.00933f
C5962 x5.X.n50 VSS 0.0113f
C5963 x5.X.n51 VSS 0.00288f
C5964 x5.X.n52 VSS 0.0482f
C5965 x5.X.n53 VSS 0.0661f
C5966 x5.X.n54 VSS 0.228f
C5967 x5.X.n55 VSS 0.00462f
C5968 x5.X.n56 VSS 0.00187f
C5969 x5.X.t23 VSS 0.0126f
C5970 x5.X.n57 VSS 0.0129f
C5971 x5.X.n58 VSS 0.00145f
C5972 x5.X.t10 VSS 0.00941f
C5973 x5.X.n59 VSS 0.0114f
C5974 x5.X.n60 VSS 0.00273f
C5975 x5.X.n61 VSS 0.0404f
C5976 x5.X.n62 VSS 0.217f
C5977 x5.X.n63 VSS 0.00462f
C5978 x5.X.n64 VSS 0.00187f
C5979 x5.X.t12 VSS 0.0126f
C5980 x5.X.n65 VSS 0.0129f
C5981 x5.X.n66 VSS 0.00145f
C5982 x5.X.t16 VSS 0.00941f
C5983 x5.X.n67 VSS 0.0114f
C5984 x5.X.n68 VSS 0.00273f
C5985 x5.X.n69 VSS 0.00444f
C5986 x5.X.n70 VSS 0.00418f
C5987 x5.X.n71 VSS 0.186f
C5988 x5.X.t2 VSS 0.00838f
C5989 x5.X.t0 VSS 0.00838f
C5990 x5.X.n72 VSS 0.0225f
C5991 x5.X.t3 VSS 0.00838f
C5992 x5.X.t1 VSS 0.00838f
C5993 x5.X.n73 VSS 0.0191f
C5994 x5.X.n74 VSS 0.0466f
C5995 x5.X.n75 VSS 0.0293f
C5996 x5.X.t4 VSS 0.00545f
C5997 x5.X.t6 VSS 0.00545f
C5998 x5.X.n76 VSS 0.0155f
C5999 x5.X.t5 VSS 0.00545f
C6000 x5.X.t7 VSS 0.00545f
C6001 x5.X.n77 VSS 0.012f
C6002 x5.X.n78 VSS 0.0268f
C6003 eob.t8 VSS 0.0344f
C6004 eob.t9 VSS 0.0215f
C6005 eob.n0 VSS 0.0657f
C6006 eob.t4 VSS 0.0208f
C6007 eob.t2 VSS 0.0208f
C6008 eob.n1 VSS 0.0606f
C6009 eob.t7 VSS 0.0135f
C6010 eob.t5 VSS 0.0135f
C6011 eob.n2 VSS 0.0404f
C6012 eob.n3 VSS 0.184f
C6013 eob.t1 VSS 0.0208f
C6014 eob.t3 VSS 0.0208f
C6015 eob.n4 VSS 0.0421f
C6016 eob.n5 VSS 0.017f
C6017 eob.n6 VSS 0.0382f
C6018 eob.t0 VSS 0.0135f
C6019 eob.t6 VSS 0.0135f
C6020 eob.n7 VSS 0.027f
C6021 eob.n8 VSS 0.017f
C6022 eob.n9 VSS 0.0976f
C6023 eob.t11 VSS 0.0279f
C6024 eob.t10 VSS 0.0194f
C6025 eob.n10 VSS 0.0567f
C6026 eob.n11 VSS 0.0214f
C6027 eob.n12 VSS 0.574f
C6028 eob.n13 VSS 0.595f
C6029 check[1].t1 VSS 0.046f
C6030 check[1].n0 VSS 0.00347f
C6031 check[1].t3 VSS 0.0153f
C6032 check[1].t2 VSS 0.0227f
C6033 check[1].n1 VSS 0.0487f
C6034 check[1].n2 VSS 0.582f
C6035 check[1].t5 VSS 0.0215f
C6036 check[1].t4 VSS 0.0149f
C6037 check[1].n3 VSS 0.0436f
C6038 check[1].n4 VSS 0.0165f
C6039 check[1].n5 VSS 0.733f
C6040 check[1].n6 VSS 0.0312f
C6041 check[1].n7 VSS 0.227f
C6042 check[1].t0 VSS 0.0177f
C6043 check[1].n8 VSS 0.0291f
C6044 VDD.n0 VSS 0.00122f
C6045 VDD.t708 VSS 4.05e-19
C6046 VDD.t626 VSS 4.05e-19
C6047 VDD.n1 VSS 8.77e-19
C6048 VDD.t707 VSS 0.0039f
C6049 VDD.n2 VSS 0.00525f
C6050 VDD.n3 VSS 7.34e-19
C6051 VDD.n4 VSS 0.00122f
C6052 VDD.t736 VSS 4.05e-19
C6053 VDD.t684 VSS 4.05e-19
C6054 VDD.n5 VSS 8.77e-19
C6055 VDD.t735 VSS 0.0039f
C6056 VDD.n6 VSS 0.00525f
C6057 VDD.n7 VSS 7.34e-19
C6058 VDD.n8 VSS 0.00122f
C6059 VDD.t301 VSS 4.05e-19
C6060 VDD.t686 VSS 4.05e-19
C6061 VDD.n9 VSS 8.77e-19
C6062 VDD.t300 VSS 0.0039f
C6063 VDD.n10 VSS 0.00525f
C6064 VDD.n11 VSS 7.34e-19
C6065 VDD.n12 VSS 0.00207f
C6066 VDD.t212 VSS 5.37e-19
C6067 VDD.t236 VSS 5.37e-19
C6068 VDD.n13 VSS 0.0013f
C6069 VDD.n14 VSS 0.00246f
C6070 VDD.n15 VSS 0.00136f
C6071 VDD.n16 VSS 7.44e-19
C6072 VDD.n17 VSS 7.34e-19
C6073 VDD.n18 VSS 0.00207f
C6074 VDD.t601 VSS 6.33e-19
C6075 VDD.t661 VSS 6.33e-19
C6076 VDD.n19 VSS 0.00145f
C6077 VDD.n20 VSS 0.00225f
C6078 VDD.n21 VSS 7.34e-19
C6079 VDD.t602 VSS 0.00394f
C6080 VDD.n22 VSS 7.34e-19
C6081 VDD.n23 VSS 6.94e-19
C6082 VDD.t603 VSS 6.33e-19
C6083 VDD.t599 VSS 6.33e-19
C6084 VDD.n24 VSS 0.0015f
C6085 VDD.n25 VSS 0.00257f
C6086 VDD.n26 VSS 4.9e-19
C6087 VDD.n27 VSS 3.67e-19
C6088 VDD.n28 VSS 0.0012f
C6089 VDD.n29 VSS 3.27e-19
C6090 VDD.n30 VSS 4.42e-19
C6091 VDD.t577 VSS 0.00252f
C6092 VDD.n31 VSS 0.00189f
C6093 VDD.n32 VSS 1.91e-19
C6094 VDD.n33 VSS 1.16e-19
C6095 VDD.n34 VSS 9.57e-19
C6096 VDD.n35 VSS 6.78e-20
C6097 VDD.t570 VSS 0.00321f
C6098 VDD.n36 VSS 3.39e-19
C6099 VDD.t567 VSS 6.33e-19
C6100 VDD.t571 VSS 6.33e-19
C6101 VDD.n37 VSS 0.00144f
C6102 VDD.n38 VSS 1.16e-19
C6103 VDD.n39 VSS 9.23e-19
C6104 VDD.n40 VSS 4.42e-19
C6105 VDD.n41 VSS 3.27e-19
C6106 VDD.n42 VSS 5.99e-19
C6107 VDD.n43 VSS 6.78e-20
C6108 VDD.n44 VSS 1.16e-19
C6109 VDD.n45 VSS 4.42e-19
C6110 VDD.n46 VSS 1.16e-19
C6111 VDD.n47 VSS 1.91e-19
C6112 VDD.n48 VSS 1.16e-19
C6113 VDD.t569 VSS 6.33e-19
C6114 VDD.t573 VSS 6.33e-19
C6115 VDD.n49 VSS 0.00144f
C6116 VDD.n50 VSS 3.39e-19
C6117 VDD.n51 VSS 0.00343f
C6118 VDD.n52 VSS 3.27e-19
C6119 VDD.n53 VSS 4.42e-19
C6120 VDD.n54 VSS 1.91e-19
C6121 VDD.n55 VSS 1.16e-19
C6122 VDD.n56 VSS 9.57e-19
C6123 VDD.n57 VSS 6.78e-20
C6124 VDD.t354 VSS 0.00321f
C6125 VDD.n58 VSS 3.39e-19
C6126 VDD.t355 VSS 6.33e-19
C6127 VDD.t575 VSS 6.33e-19
C6128 VDD.n59 VSS 0.00144f
C6129 VDD.n60 VSS 1.16e-19
C6130 VDD.n61 VSS 9.23e-19
C6131 VDD.n62 VSS 4.42e-19
C6132 VDD.n63 VSS 3.27e-19
C6133 VDD.n64 VSS 7.28e-19
C6134 VDD.n65 VSS 6.78e-20
C6135 VDD.n66 VSS 1.16e-19
C6136 VDD.n67 VSS 4.42e-19
C6137 VDD.n68 VSS 1.16e-19
C6138 VDD.n69 VSS 1.91e-19
C6139 VDD.n70 VSS 1.16e-19
C6140 VDD.t377 VSS 6.33e-19
C6141 VDD.t365 VSS 6.33e-19
C6142 VDD.n71 VSS 0.00144f
C6143 VDD.n72 VSS 3.39e-19
C6144 VDD.n73 VSS 0.00205f
C6145 VDD.n74 VSS 3.27e-19
C6146 VDD.n75 VSS 4.42e-19
C6147 VDD.n76 VSS 1.91e-19
C6148 VDD.t379 VSS 6.33e-19
C6149 VDD.t369 VSS 6.33e-19
C6150 VDD.n77 VSS 0.00144f
C6151 VDD.n78 VSS 0.00117f
C6152 VDD.n79 VSS 0.00104f
C6153 VDD.n80 VSS 6.78e-20
C6154 VDD.t378 VSS 0.00278f
C6155 VDD.n81 VSS 2.99e-19
C6156 VDD.n82 VSS 1.84e-19
C6157 VDD.n83 VSS 0.00207f
C6158 VDD.t383 VSS 6.33e-19
C6159 VDD.t371 VSS 6.33e-19
C6160 VDD.n84 VSS 0.00144f
C6161 VDD.n85 VSS 0.00173f
C6162 VDD.n86 VSS 6.26e-19
C6163 VDD.n87 VSS 1.08e-19
C6164 VDD.t362 VSS 0.00394f
C6165 VDD.n88 VSS 7.34e-19
C6166 VDD.t353 VSS 6.33e-19
C6167 VDD.t363 VSS 6.33e-19
C6168 VDD.n89 VSS 0.00144f
C6169 VDD.n90 VSS 0.00105f
C6170 VDD.n91 VSS 0.00207f
C6171 VDD.n92 VSS 9.39e-19
C6172 VDD.n93 VSS 7.34e-19
C6173 VDD.n94 VSS 7.34e-19
C6174 VDD.t358 VSS 0.00394f
C6175 VDD.n95 VSS 7.34e-19
C6176 VDD.n96 VSS 8.3e-19
C6177 VDD.t381 VSS 6.33e-19
C6178 VDD.t375 VSS 6.33e-19
C6179 VDD.n97 VSS 0.00144f
C6180 VDD.n98 VSS 0.00173f
C6181 VDD.n99 VSS 0.00207f
C6182 VDD.n100 VSS 7.21e-19
C6183 VDD.n101 VSS 7.34e-19
C6184 VDD.n102 VSS 0.00599f
C6185 VDD.n103 VSS 7.34e-19
C6186 VDD.n104 VSS 0.00101f
C6187 VDD.t361 VSS 0.00235f
C6188 VDD.n105 VSS 0.00199f
C6189 VDD.n106 VSS 0.00207f
C6190 VDD.t555 VSS 5.71e-19
C6191 VDD.t126 VSS -1.82e-19
C6192 VDD.n107 VSS 0.00268f
C6193 VDD.n108 VSS 7.44e-19
C6194 VDD.n109 VSS 0.0012f
C6195 VDD.n110 VSS 7.34e-19
C6196 VDD.t40 VSS 0.00394f
C6197 VDD.n111 VSS 7.34e-19
C6198 VDD.t41 VSS 6.16e-19
C6199 VDD.t551 VSS -3.41e-19
C6200 VDD.n112 VSS 0.00241f
C6201 VDD.n113 VSS 0.00164f
C6202 VDD.n114 VSS 0.00207f
C6203 VDD.t240 VSS 0.00176f
C6204 VDD.n115 VSS 0.00177f
C6205 VDD.n116 VSS 0.00112f
C6206 VDD.n117 VSS 0.00428f
C6207 VDD.n118 VSS 7.34e-19
C6208 VDD.n119 VSS 0.00125f
C6209 VDD.n120 VSS 0.00207f
C6210 VDD.n121 VSS 0.00125f
C6211 VDD.n122 VSS 7.34e-19
C6212 VDD.n123 VSS 0.00415f
C6213 VDD.n124 VSS 7.34e-19
C6214 VDD.t238 VSS 6.5e-19
C6215 VDD.t513 VSS 0.00146f
C6216 VDD.n125 VSS 0.00234f
C6217 VDD.n126 VSS 0.00307f
C6218 VDD.n127 VSS 0.00207f
C6219 VDD.n128 VSS 7.89e-19
C6220 VDD.n129 VSS 7.34e-19
C6221 VDD.t510 VSS 0.00394f
C6222 VDD.n130 VSS 7.34e-19
C6223 VDD.n131 VSS 0.0012f
C6224 VDD.n132 VSS 0.00207f
C6225 VDD.n133 VSS 0.00101f
C6226 VDD.n134 VSS 7.34e-19
C6227 VDD.n135 VSS 0.00617f
C6228 VDD.n136 VSS 7.34e-19
C6229 VDD.n137 VSS 8.03e-19
C6230 VDD.t688 VSS 4.05e-19
C6231 VDD.t67 VSS 4.05e-19
C6232 VDD.n138 VSS 8.77e-19
C6233 VDD.n139 VSS 0.00101f
C6234 VDD.n140 VSS 7.34e-19
C6235 VDD.t38 VSS 0.00394f
C6236 VDD.n141 VSS 7.44e-19
C6237 VDD.n142 VSS 0.00134f
C6238 VDD.n143 VSS 0.00207f
C6239 VDD.n144 VSS 0.0012f
C6240 VDD.n145 VSS 7.34e-19
C6241 VDD.t294 VSS 0.00394f
C6242 VDD.n146 VSS 7.34e-19
C6243 VDD.t295 VSS 6.16e-19
C6244 VDD.t430 VSS -3.41e-19
C6245 VDD.n147 VSS 0.00241f
C6246 VDD.n148 VSS 0.00164f
C6247 VDD.n149 VSS 0.00207f
C6248 VDD.t116 VSS 0.00176f
C6249 VDD.n150 VSS 0.00177f
C6250 VDD.n151 VSS 0.00112f
C6251 VDD.n152 VSS 0.00428f
C6252 VDD.n153 VSS 7.34e-19
C6253 VDD.n154 VSS 0.00125f
C6254 VDD.n155 VSS 0.00207f
C6255 VDD.n156 VSS 0.00125f
C6256 VDD.n157 VSS 7.34e-19
C6257 VDD.n158 VSS 0.00415f
C6258 VDD.n159 VSS 7.34e-19
C6259 VDD.t118 VSS 6.5e-19
C6260 VDD.t702 VSS 0.00146f
C6261 VDD.n160 VSS 0.00234f
C6262 VDD.n161 VSS 0.00307f
C6263 VDD.n162 VSS 0.00207f
C6264 VDD.n163 VSS 7.89e-19
C6265 VDD.n164 VSS 7.34e-19
C6266 VDD.t703 VSS 0.00394f
C6267 VDD.n165 VSS 7.34e-19
C6268 VDD.n166 VSS 0.0012f
C6269 VDD.n167 VSS 0.00207f
C6270 VDD.n168 VSS 0.00101f
C6271 VDD.n169 VSS 7.34e-19
C6272 VDD.n170 VSS 0.00617f
C6273 VDD.n171 VSS 7.34e-19
C6274 VDD.n172 VSS 8.03e-19
C6275 VDD.t692 VSS 4.05e-19
C6276 VDD.t682 VSS 4.05e-19
C6277 VDD.n173 VSS 8.77e-19
C6278 VDD.n174 VSS 0.00101f
C6279 VDD.n175 VSS 7.34e-19
C6280 VDD.t85 VSS 0.00394f
C6281 VDD.n176 VSS 7.44e-19
C6282 VDD.n177 VSS 0.00134f
C6283 VDD.n178 VSS 0.00207f
C6284 VDD.n179 VSS 0.0012f
C6285 VDD.n180 VSS 7.34e-19
C6286 VDD.t109 VSS 0.00394f
C6287 VDD.n181 VSS 7.34e-19
C6288 VDD.t110 VSS 6.16e-19
C6289 VDD.t15 VSS -3.41e-19
C6290 VDD.n182 VSS 0.00241f
C6291 VDD.n183 VSS 0.00164f
C6292 VDD.n184 VSS 0.00207f
C6293 VDD.t438 VSS 0.00176f
C6294 VDD.n185 VSS 0.00177f
C6295 VDD.n186 VSS 0.00112f
C6296 VDD.n187 VSS 0.00428f
C6297 VDD.n188 VSS 7.34e-19
C6298 VDD.n189 VSS 0.00125f
C6299 VDD.n190 VSS 0.00207f
C6300 VDD.n191 VSS 0.00125f
C6301 VDD.n192 VSS 7.34e-19
C6302 VDD.n193 VSS 0.00415f
C6303 VDD.n194 VSS 7.34e-19
C6304 VDD.t440 VSS 6.5e-19
C6305 VDD.t276 VSS 0.00146f
C6306 VDD.n195 VSS 0.00234f
C6307 VDD.n196 VSS 0.00307f
C6308 VDD.n197 VSS 0.00207f
C6309 VDD.n198 VSS 7.89e-19
C6310 VDD.n199 VSS 7.34e-19
C6311 VDD.t273 VSS 0.00394f
C6312 VDD.n200 VSS 7.34e-19
C6313 VDD.n201 VSS 0.0012f
C6314 VDD.n202 VSS 0.00207f
C6315 VDD.n203 VSS 0.00101f
C6316 VDD.n204 VSS 7.34e-19
C6317 VDD.n205 VSS 0.00617f
C6318 VDD.n206 VSS 7.34e-19
C6319 VDD.n207 VSS 8.03e-19
C6320 VDD.t696 VSS 4.05e-19
C6321 VDD.t346 VSS 4.05e-19
C6322 VDD.n208 VSS 8.77e-19
C6323 VDD.n209 VSS 0.00101f
C6324 VDD.n210 VSS 7.34e-19
C6325 VDD.t6 VSS 0.00394f
C6326 VDD.n211 VSS 7.44e-19
C6327 VDD.n212 VSS 0.00134f
C6328 VDD.n213 VSS 0.00207f
C6329 VDD.n214 VSS 0.0012f
C6330 VDD.n215 VSS 7.34e-19
C6331 VDD.t288 VSS 0.00394f
C6332 VDD.n216 VSS 7.34e-19
C6333 VDD.t289 VSS 6.16e-19
C6334 VDD.t460 VSS -3.41e-19
C6335 VDD.n217 VSS 0.00241f
C6336 VDD.n218 VSS 0.00164f
C6337 VDD.n219 VSS 0.00207f
C6338 VDD.t278 VSS 0.00176f
C6339 VDD.n220 VSS 0.00177f
C6340 VDD.n221 VSS 0.00112f
C6341 VDD.n222 VSS 0.00428f
C6342 VDD.n223 VSS 7.34e-19
C6343 VDD.n224 VSS 0.00125f
C6344 VDD.n225 VSS 0.00207f
C6345 VDD.n226 VSS 0.00125f
C6346 VDD.n227 VSS 7.34e-19
C6347 VDD.n228 VSS 0.00415f
C6348 VDD.n229 VSS 7.34e-19
C6349 VDD.t280 VSS 6.5e-19
C6350 VDD.t389 VSS 0.00146f
C6351 VDD.n230 VSS 0.00234f
C6352 VDD.n231 VSS 0.00307f
C6353 VDD.n232 VSS 0.00207f
C6354 VDD.n233 VSS 7.89e-19
C6355 VDD.n234 VSS 7.34e-19
C6356 VDD.t390 VSS 0.00394f
C6357 VDD.n235 VSS 7.34e-19
C6358 VDD.n236 VSS 0.0012f
C6359 VDD.n237 VSS 0.00207f
C6360 VDD.n238 VSS 0.00101f
C6361 VDD.n239 VSS 7.34e-19
C6362 VDD.n240 VSS 0.00617f
C6363 VDD.n241 VSS 7.34e-19
C6364 VDD.n242 VSS 8.03e-19
C6365 VDD.t634 VSS 4.05e-19
C6366 VDD.t3 VSS 4.05e-19
C6367 VDD.n243 VSS 8.77e-19
C6368 VDD.n244 VSS 7.44e-19
C6369 VDD.t2 VSS 0.00394f
C6370 VDD.n245 VSS 0.0036f
C6371 VDD.t633 VSS 0.00317f
C6372 VDD.n246 VSS 0.00262f
C6373 VDD.n247 VSS 0.00103f
C6374 VDD.n248 VSS 0.00136f
C6375 VDD.n249 VSS 0.00182f
C6376 VDD.n250 VSS 0.00187f
C6377 VDD.n251 VSS 0.00207f
C6378 VDD.n252 VSS 0.00207f
C6379 VDD.t74 VSS 9.52e-19
C6380 VDD.n253 VSS 0.00207f
C6381 VDD.n254 VSS 0.00136f
C6382 VDD.n255 VSS 7.44e-19
C6383 VDD.n256 VSS 0.00582f
C6384 VDD.t73 VSS 0.00394f
C6385 VDD.n257 VSS 0.00398f
C6386 VDD.t503 VSS 0.00394f
C6387 VDD.n258 VSS 0.00514f
C6388 VDD.t1 VSS 0.00394f
C6389 VDD.n259 VSS 0.0036f
C6390 VDD.n260 VSS 7.34e-19
C6391 VDD.n261 VSS 0.00125f
C6392 VDD.n262 VSS 0.00207f
C6393 VDD.n263 VSS 0.00207f
C6394 VDD.n264 VSS 0.00207f
C6395 VDD.n265 VSS 0.00207f
C6396 VDD.t391 VSS 3.65e-19
C6397 VDD.t171 VSS 3.84e-19
C6398 VDD.n266 VSS 8.01e-19
C6399 VDD.n267 VSS 0.00187f
C6400 VDD.n268 VSS 0.00137f
C6401 VDD.n269 VSS 7.44e-19
C6402 VDD.n270 VSS 0.00454f
C6403 VDD.t170 VSS 0.00394f
C6404 VDD.n271 VSS 0.0045f
C6405 VDD.t279 VSS 0.00381f
C6406 VDD.t524 VSS 0.00372f
C6407 VDD.n272 VSS 0.00407f
C6408 VDD.n273 VSS 7.34e-19
C6409 VDD.n274 VSS 0.00125f
C6410 VDD.n275 VSS 6.94e-19
C6411 VDD.n276 VSS 0.00207f
C6412 VDD.n277 VSS 0.00207f
C6413 VDD.n278 VSS 7.35e-19
C6414 VDD.n279 VSS 7.34e-19
C6415 VDD.n280 VSS 0.00565f
C6416 VDD.t388 VSS 0.00394f
C6417 VDD.n281 VSS 0.00617f
C6418 VDD.t502 VSS 0.00394f
C6419 VDD.t0 VSS 0.00754f
C6420 VDD.n282 VSS 7.34e-19
C6421 VDD.n283 VSS 0.00125f
C6422 VDD.n284 VSS 0.00207f
C6423 VDD.n285 VSS 0.00207f
C6424 VDD.n286 VSS 0.00207f
C6425 VDD.n287 VSS 1.32e-19
C6426 VDD.t757 VSS 4.24e-19
C6427 VDD.t169 VSS 0.001f
C6428 VDD.n288 VSS 0.00209f
C6429 VDD.n289 VSS 3.57e-19
C6430 VDD.n290 VSS 7.07e-19
C6431 VDD.n291 VSS 0.00261f
C6432 VDD.n292 VSS 4.15e-19
C6433 VDD.n293 VSS 3.73e-19
C6434 VDD.t753 VSS 4.18e-19
C6435 VDD.n294 VSS 3.02e-19
C6436 VDD.n295 VSS 6.43e-19
C6437 VDD.n296 VSS 0.00133f
C6438 VDD.t145 VSS 0.00157f
C6439 VDD.n297 VSS 0.00118f
C6440 VDD.t462 VSS 3.84e-19
C6441 VDD.t147 VSS 3.84e-19
C6442 VDD.n298 VSS 8.1e-19
C6443 VDD.n299 VSS 0.00207f
C6444 VDD.n300 VSS 0.00105f
C6445 VDD.n301 VSS 0.00101f
C6446 VDD.n302 VSS 0.00207f
C6447 VDD.n303 VSS 0.00207f
C6448 VDD.n304 VSS 0.00172f
C6449 VDD.n305 VSS 9.71e-19
C6450 VDD.n306 VSS 8.91e-19
C6451 VDD.n307 VSS 9.41e-19
C6452 VDD.n308 VSS 0.00471f
C6453 VDD.t461 VSS 0.00539f
C6454 VDD.t146 VSS 0.00873f
C6455 VDD.t257 VSS 0.00642f
C6456 VDD.n309 VSS 0.00308f
C6457 VDD.t277 VSS 0.00394f
C6458 VDD.n310 VSS 0.00531f
C6459 VDD.n311 VSS 0.00711f
C6460 VDD.n312 VSS 7.34e-19
C6461 VDD.n313 VSS 0.00195f
C6462 VDD.n314 VSS 0.00281f
C6463 VDD.n315 VSS 0.00207f
C6464 VDD.n316 VSS 0.00207f
C6465 VDD.n317 VSS 0.00125f
C6466 VDD.n318 VSS 7.34e-19
C6467 VDD.n319 VSS 0.00415f
C6468 VDD.t459 VSS 0.00394f
C6469 VDD.n320 VSS 0.00629f
C6470 VDD.n321 VSS 0.00407f
C6471 VDD.t463 VSS 0.00394f
C6472 VDD.n322 VSS 0.00569f
C6473 VDD.n323 VSS 7.34e-19
C6474 VDD.n324 VSS 0.00109f
C6475 VDD.n325 VSS 0.00207f
C6476 VDD.t464 VSS 5.71e-19
C6477 VDD.t7 VSS -1.82e-19
C6478 VDD.n326 VSS 0.00268f
C6479 VDD.n327 VSS 0.00243f
C6480 VDD.n328 VSS 0.00207f
C6481 VDD.n329 VSS 7.21e-19
C6482 VDD.n330 VSS 0.00155f
C6483 VDD.n331 VSS 0.00101f
C6484 VDD.n332 VSS 7.34e-19
C6485 VDD.n333 VSS 0.00599f
C6486 VDD.n334 VSS 0.00398f
C6487 VDD.t695 VSS 0.00317f
C6488 VDD.t345 VSS 0.00394f
C6489 VDD.n335 VSS 0.0036f
C6490 VDD.n336 VSS 7.44e-19
C6491 VDD.n337 VSS 0.00136f
C6492 VDD.n338 VSS 0.00182f
C6493 VDD.n339 VSS 0.00187f
C6494 VDD.n340 VSS 0.00207f
C6495 VDD.n341 VSS 0.00207f
C6496 VDD.t114 VSS 9.52e-19
C6497 VDD.n342 VSS 0.00207f
C6498 VDD.n343 VSS 0.00136f
C6499 VDD.n344 VSS 7.44e-19
C6500 VDD.n345 VSS 0.00582f
C6501 VDD.t113 VSS 0.00394f
C6502 VDD.n346 VSS 0.00398f
C6503 VDD.t210 VSS 0.00394f
C6504 VDD.n347 VSS 0.00514f
C6505 VDD.t348 VSS 0.00394f
C6506 VDD.n348 VSS 0.0036f
C6507 VDD.n349 VSS 7.34e-19
C6508 VDD.n350 VSS 0.00125f
C6509 VDD.n351 VSS 0.00207f
C6510 VDD.n352 VSS 0.00207f
C6511 VDD.n353 VSS 0.00207f
C6512 VDD.n354 VSS 0.00207f
C6513 VDD.t274 VSS 3.65e-19
C6514 VDD.t177 VSS 3.84e-19
C6515 VDD.n355 VSS 8.01e-19
C6516 VDD.n356 VSS 0.00187f
C6517 VDD.n357 VSS 0.00137f
C6518 VDD.n358 VSS 7.44e-19
C6519 VDD.n359 VSS 0.00454f
C6520 VDD.t176 VSS 0.00394f
C6521 VDD.n360 VSS 0.0045f
C6522 VDD.t439 VSS 0.00381f
C6523 VDD.t30 VSS 0.00372f
C6524 VDD.n361 VSS 0.00407f
C6525 VDD.n362 VSS 7.34e-19
C6526 VDD.n363 VSS 0.00125f
C6527 VDD.n364 VSS 6.94e-19
C6528 VDD.n365 VSS 0.00207f
C6529 VDD.n366 VSS 0.00207f
C6530 VDD.n367 VSS 7.35e-19
C6531 VDD.n368 VSS 7.34e-19
C6532 VDD.n369 VSS 0.00565f
C6533 VDD.t275 VSS 0.00394f
C6534 VDD.n370 VSS 0.00617f
C6535 VDD.t209 VSS 0.00394f
C6536 VDD.t347 VSS 0.00754f
C6537 VDD.n371 VSS 7.34e-19
C6538 VDD.n372 VSS 0.00125f
C6539 VDD.n373 VSS 0.00207f
C6540 VDD.n374 VSS 0.00207f
C6541 VDD.n375 VSS 0.00207f
C6542 VDD.n376 VSS 1.32e-19
C6543 VDD.t745 VSS 4.24e-19
C6544 VDD.t175 VSS 0.001f
C6545 VDD.n377 VSS 0.00209f
C6546 VDD.n378 VSS 3.57e-19
C6547 VDD.n379 VSS 7.07e-19
C6548 VDD.n380 VSS 0.00261f
C6549 VDD.n381 VSS 4.15e-19
C6550 VDD.n382 VSS 3.73e-19
C6551 VDD.t744 VSS 4.18e-19
C6552 VDD.n383 VSS 3.02e-19
C6553 VDD.n384 VSS 6.43e-19
C6554 VDD.n385 VSS 0.00133f
C6555 VDD.t166 VSS 0.00157f
C6556 VDD.n386 VSS 0.00118f
C6557 VDD.t17 VSS 3.84e-19
C6558 VDD.t168 VSS 3.84e-19
C6559 VDD.n387 VSS 8.1e-19
C6560 VDD.n388 VSS 0.00207f
C6561 VDD.n389 VSS 0.00105f
C6562 VDD.n390 VSS 0.00101f
C6563 VDD.n391 VSS 0.00207f
C6564 VDD.n392 VSS 0.00207f
C6565 VDD.n393 VSS 0.00172f
C6566 VDD.n394 VSS 9.71e-19
C6567 VDD.n395 VSS 8.91e-19
C6568 VDD.n396 VSS 9.41e-19
C6569 VDD.n397 VSS 0.00471f
C6570 VDD.t16 VSS 0.00539f
C6571 VDD.t167 VSS 0.00873f
C6572 VDD.t57 VSS 0.00642f
C6573 VDD.n398 VSS 0.00308f
C6574 VDD.t437 VSS 0.00394f
C6575 VDD.n399 VSS 0.00531f
C6576 VDD.n400 VSS 0.00711f
C6577 VDD.n401 VSS 7.34e-19
C6578 VDD.n402 VSS 0.00195f
C6579 VDD.n403 VSS 0.00281f
C6580 VDD.n404 VSS 0.00207f
C6581 VDD.n405 VSS 0.00207f
C6582 VDD.n406 VSS 0.00125f
C6583 VDD.n407 VSS 7.34e-19
C6584 VDD.n408 VSS 0.00415f
C6585 VDD.t14 VSS 0.00394f
C6586 VDD.n409 VSS 0.00629f
C6587 VDD.n410 VSS 0.00407f
C6588 VDD.t18 VSS 0.00394f
C6589 VDD.n411 VSS 0.00569f
C6590 VDD.n412 VSS 7.34e-19
C6591 VDD.n413 VSS 0.00109f
C6592 VDD.n414 VSS 0.00207f
C6593 VDD.t19 VSS 5.71e-19
C6594 VDD.t86 VSS -1.82e-19
C6595 VDD.n415 VSS 0.00268f
C6596 VDD.n416 VSS 0.00243f
C6597 VDD.n417 VSS 0.00207f
C6598 VDD.n418 VSS 7.21e-19
C6599 VDD.n419 VSS 0.00155f
C6600 VDD.n420 VSS 0.00101f
C6601 VDD.n421 VSS 7.34e-19
C6602 VDD.n422 VSS 0.00599f
C6603 VDD.n423 VSS 0.00398f
C6604 VDD.t691 VSS 0.00317f
C6605 VDD.t681 VSS 0.00394f
C6606 VDD.n424 VSS 0.0036f
C6607 VDD.n425 VSS 7.44e-19
C6608 VDD.n426 VSS 0.00136f
C6609 VDD.n427 VSS 0.00182f
C6610 VDD.n428 VSS 0.00187f
C6611 VDD.n429 VSS 0.00207f
C6612 VDD.n430 VSS 0.00207f
C6613 VDD.t466 VSS 9.52e-19
C6614 VDD.n431 VSS 0.00207f
C6615 VDD.n432 VSS 0.00136f
C6616 VDD.n433 VSS 7.44e-19
C6617 VDD.n434 VSS 0.00582f
C6618 VDD.t465 VSS 0.00394f
C6619 VDD.n435 VSS 0.00398f
C6620 VDD.t482 VSS 0.00394f
C6621 VDD.n436 VSS 0.00514f
C6622 VDD.t680 VSS 0.00394f
C6623 VDD.n437 VSS 0.0036f
C6624 VDD.n438 VSS 7.34e-19
C6625 VDD.n439 VSS 0.00125f
C6626 VDD.n440 VSS 0.00207f
C6627 VDD.n441 VSS 0.00207f
C6628 VDD.n442 VSS 0.00207f
C6629 VDD.n443 VSS 0.00207f
C6630 VDD.t704 VSS 3.65e-19
C6631 VDD.t156 VSS 3.84e-19
C6632 VDD.n444 VSS 8.01e-19
C6633 VDD.n445 VSS 0.00187f
C6634 VDD.n446 VSS 0.00137f
C6635 VDD.n447 VSS 7.44e-19
C6636 VDD.n448 VSS 0.00454f
C6637 VDD.t155 VSS 0.00394f
C6638 VDD.n449 VSS 0.0045f
C6639 VDD.t117 VSS 0.00381f
C6640 VDD.t97 VSS 0.00372f
C6641 VDD.n450 VSS 0.00407f
C6642 VDD.n451 VSS 7.34e-19
C6643 VDD.n452 VSS 0.00125f
C6644 VDD.n453 VSS 6.94e-19
C6645 VDD.n454 VSS 0.00207f
C6646 VDD.n455 VSS 0.00207f
C6647 VDD.n456 VSS 7.35e-19
C6648 VDD.n457 VSS 7.34e-19
C6649 VDD.n458 VSS 0.00565f
C6650 VDD.t701 VSS 0.00394f
C6651 VDD.n459 VSS 0.00617f
C6652 VDD.t481 VSS 0.00394f
C6653 VDD.t679 VSS 0.00754f
C6654 VDD.n460 VSS 7.34e-19
C6655 VDD.n461 VSS 0.00125f
C6656 VDD.n462 VSS 0.00207f
C6657 VDD.n463 VSS 0.00207f
C6658 VDD.n464 VSS 0.00207f
C6659 VDD.n465 VSS 1.32e-19
C6660 VDD.t751 VSS 4.24e-19
C6661 VDD.t154 VSS 0.001f
C6662 VDD.n466 VSS 0.00209f
C6663 VDD.n467 VSS 3.57e-19
C6664 VDD.n468 VSS 7.07e-19
C6665 VDD.n469 VSS 0.00261f
C6666 VDD.n470 VSS 4.15e-19
C6667 VDD.n471 VSS 3.73e-19
C6668 VDD.t746 VSS 4.18e-19
C6669 VDD.n472 VSS 3.02e-19
C6670 VDD.n473 VSS 6.43e-19
C6671 VDD.n474 VSS 0.00133f
C6672 VDD.t163 VSS 0.00157f
C6673 VDD.n475 VSS 0.00118f
C6674 VDD.t432 VSS 3.84e-19
C6675 VDD.t165 VSS 3.84e-19
C6676 VDD.n476 VSS 8.1e-19
C6677 VDD.n477 VSS 0.00207f
C6678 VDD.n478 VSS 0.00105f
C6679 VDD.n479 VSS 0.00101f
C6680 VDD.n480 VSS 0.00207f
C6681 VDD.n481 VSS 0.00207f
C6682 VDD.n482 VSS 0.00172f
C6683 VDD.n483 VSS 9.71e-19
C6684 VDD.n484 VSS 8.91e-19
C6685 VDD.n485 VSS 9.41e-19
C6686 VDD.n486 VSS 0.00471f
C6687 VDD.t431 VSS 0.00539f
C6688 VDD.t164 VSS 0.00873f
C6689 VDD.t662 VSS 0.00642f
C6690 VDD.n487 VSS 0.00308f
C6691 VDD.t115 VSS 0.00394f
C6692 VDD.n488 VSS 0.00531f
C6693 VDD.n489 VSS 0.00711f
C6694 VDD.n490 VSS 7.34e-19
C6695 VDD.n491 VSS 0.00195f
C6696 VDD.n492 VSS 0.00281f
C6697 VDD.n493 VSS 0.00207f
C6698 VDD.n494 VSS 0.00207f
C6699 VDD.n495 VSS 0.00125f
C6700 VDD.n496 VSS 7.34e-19
C6701 VDD.n497 VSS 0.00415f
C6702 VDD.t429 VSS 0.00394f
C6703 VDD.n498 VSS 0.00629f
C6704 VDD.n499 VSS 0.00407f
C6705 VDD.t433 VSS 0.00394f
C6706 VDD.n500 VSS 0.00569f
C6707 VDD.n501 VSS 7.34e-19
C6708 VDD.n502 VSS 0.00109f
C6709 VDD.n503 VSS 0.00207f
C6710 VDD.t434 VSS 5.71e-19
C6711 VDD.t39 VSS -1.82e-19
C6712 VDD.n504 VSS 0.00268f
C6713 VDD.n505 VSS 0.00243f
C6714 VDD.n506 VSS 0.00207f
C6715 VDD.n507 VSS 7.21e-19
C6716 VDD.n508 VSS 0.00155f
C6717 VDD.n509 VSS 0.00101f
C6718 VDD.n510 VSS 7.34e-19
C6719 VDD.n511 VSS 0.00599f
C6720 VDD.n512 VSS 0.00398f
C6721 VDD.t687 VSS 0.00317f
C6722 VDD.t66 VSS 0.00394f
C6723 VDD.n513 VSS 0.0036f
C6724 VDD.n514 VSS 7.44e-19
C6725 VDD.n515 VSS 0.00136f
C6726 VDD.n516 VSS 0.00182f
C6727 VDD.n517 VSS 0.00187f
C6728 VDD.n518 VSS 0.00207f
C6729 VDD.n519 VSS 0.00207f
C6730 VDD.t428 VSS 9.52e-19
C6731 VDD.n520 VSS 0.00207f
C6732 VDD.n521 VSS 0.00136f
C6733 VDD.n522 VSS 7.44e-19
C6734 VDD.n523 VSS 0.00582f
C6735 VDD.t427 VSS 0.00394f
C6736 VDD.n524 VSS 0.00398f
C6737 VDD.t435 VSS 0.00394f
C6738 VDD.n525 VSS 0.00514f
C6739 VDD.t65 VSS 0.00394f
C6740 VDD.n526 VSS 0.0036f
C6741 VDD.n527 VSS 7.34e-19
C6742 VDD.n528 VSS 0.00125f
C6743 VDD.n529 VSS 0.00207f
C6744 VDD.n530 VSS 0.00207f
C6745 VDD.n531 VSS 0.00207f
C6746 VDD.n532 VSS 0.00207f
C6747 VDD.t511 VSS 3.65e-19
C6748 VDD.t141 VSS 3.84e-19
C6749 VDD.n533 VSS 8.01e-19
C6750 VDD.n534 VSS 0.00187f
C6751 VDD.n535 VSS 0.00137f
C6752 VDD.n536 VSS 7.44e-19
C6753 VDD.n537 VSS 0.00454f
C6754 VDD.t140 VSS 0.00394f
C6755 VDD.n538 VSS 0.0045f
C6756 VDD.t237 VSS 0.00381f
C6757 VDD.t283 VSS 0.00372f
C6758 VDD.n539 VSS 0.00407f
C6759 VDD.n540 VSS 7.34e-19
C6760 VDD.n541 VSS 0.00125f
C6761 VDD.n542 VSS 6.94e-19
C6762 VDD.n543 VSS 0.00207f
C6763 VDD.n544 VSS 0.00207f
C6764 VDD.n545 VSS 7.35e-19
C6765 VDD.n546 VSS 7.34e-19
C6766 VDD.n547 VSS 0.00565f
C6767 VDD.t512 VSS 0.00394f
C6768 VDD.n548 VSS 0.00617f
C6769 VDD.t436 VSS 0.00394f
C6770 VDD.t64 VSS 0.00754f
C6771 VDD.n549 VSS 7.34e-19
C6772 VDD.n550 VSS 0.00125f
C6773 VDD.n551 VSS 0.00207f
C6774 VDD.n552 VSS 0.00207f
C6775 VDD.n553 VSS 0.00207f
C6776 VDD.n554 VSS 1.32e-19
C6777 VDD.t756 VSS 4.24e-19
C6778 VDD.t139 VSS 0.001f
C6779 VDD.n555 VSS 0.00209f
C6780 VDD.n556 VSS 3.57e-19
C6781 VDD.n557 VSS 7.07e-19
C6782 VDD.n558 VSS 0.00261f
C6783 VDD.n559 VSS 4.15e-19
C6784 VDD.n560 VSS 3.73e-19
C6785 VDD.t752 VSS 4.18e-19
C6786 VDD.n561 VSS 3.02e-19
C6787 VDD.n562 VSS 6.43e-19
C6788 VDD.n563 VSS 0.00133f
C6789 VDD.t148 VSS 0.00157f
C6790 VDD.n564 VSS 0.00118f
C6791 VDD.t553 VSS 3.84e-19
C6792 VDD.t150 VSS 3.84e-19
C6793 VDD.n565 VSS 8.1e-19
C6794 VDD.n566 VSS 0.00207f
C6795 VDD.n567 VSS 0.00105f
C6796 VDD.n568 VSS 0.00101f
C6797 VDD.n569 VSS 0.00207f
C6798 VDD.n570 VSS 0.00207f
C6799 VDD.n571 VSS 0.00172f
C6800 VDD.n572 VSS 9.71e-19
C6801 VDD.n573 VSS 8.91e-19
C6802 VDD.n574 VSS 9.41e-19
C6803 VDD.n575 VSS 0.00471f
C6804 VDD.t552 VSS 0.00539f
C6805 VDD.t149 VSS 0.00873f
C6806 VDD.t675 VSS 0.00642f
C6807 VDD.n576 VSS 0.00308f
C6808 VDD.t239 VSS 0.00394f
C6809 VDD.n577 VSS 0.00531f
C6810 VDD.n578 VSS 0.00711f
C6811 VDD.n579 VSS 7.34e-19
C6812 VDD.n580 VSS 0.00195f
C6813 VDD.n581 VSS 0.00281f
C6814 VDD.n582 VSS 0.00207f
C6815 VDD.n583 VSS 0.00207f
C6816 VDD.n584 VSS 0.00207f
C6817 VDD.n585 VSS 0.00125f
C6818 VDD.n586 VSS 7.34e-19
C6819 VDD.n587 VSS 0.00415f
C6820 VDD.t550 VSS 0.00394f
C6821 VDD.n588 VSS 0.00629f
C6822 VDD.t125 VSS 0.00394f
C6823 VDD.n589 VSS 0.00407f
C6824 VDD.t554 VSS 0.00394f
C6825 VDD.n590 VSS 0.00569f
C6826 VDD.n591 VSS 7.34e-19
C6827 VDD.n592 VSS 0.00109f
C6828 VDD.n593 VSS 0.00134f
C6829 VDD.n594 VSS 0.00243f
C6830 VDD.n595 VSS 0.00207f
C6831 VDD.n596 VSS 0.00155f
C6832 VDD.n597 VSS 0.00155f
C6833 VDD.n598 VSS 0.00116f
C6834 VDD.n599 VSS 7.34e-19
C6835 VDD.n600 VSS 0.00788f
C6836 VDD.n601 VSS 0.00514f
C6837 VDD.t360 VSS 0.00394f
C6838 VDD.n602 VSS 0.0036f
C6839 VDD.t372 VSS 0.00394f
C6840 VDD.n603 VSS 0.0036f
C6841 VDD.n604 VSS 7.34e-19
C6842 VDD.t373 VSS 6.33e-19
C6843 VDD.t359 VSS 6.33e-19
C6844 VDD.n605 VSS 0.00144f
C6845 VDD.n606 VSS 0.00173f
C6846 VDD.n607 VSS 0.00105f
C6847 VDD.n608 VSS 0.00207f
C6848 VDD.n609 VSS 0.00207f
C6849 VDD.n610 VSS 0.00207f
C6850 VDD.n611 VSS 9.39e-19
C6851 VDD.n612 VSS 7.34e-19
C6852 VDD.n613 VSS 0.0036f
C6853 VDD.t380 VSS 0.00377f
C6854 VDD.t374 VSS 0.00377f
C6855 VDD.n614 VSS 0.0036f
C6856 VDD.t356 VSS 0.00394f
C6857 VDD.n615 VSS 0.0036f
C6858 VDD.t352 VSS 0.00394f
C6859 VDD.n616 VSS 0.0036f
C6860 VDD.t366 VSS 0.00394f
C6861 VDD.n617 VSS 0.0036f
C6862 VDD.n618 VSS 7.34e-19
C6863 VDD.t357 VSS 6.33e-19
C6864 VDD.t367 VSS 6.33e-19
C6865 VDD.n619 VSS 0.00144f
C6866 VDD.n620 VSS 0.00173f
C6867 VDD.n621 VSS 8.3e-19
C6868 VDD.n622 VSS 0.00207f
C6869 VDD.n623 VSS 0.00207f
C6870 VDD.n624 VSS 0.00207f
C6871 VDD.n625 VSS 7.21e-19
C6872 VDD.n626 VSS 0.00173f
C6873 VDD.n627 VSS 0.00114f
C6874 VDD.n628 VSS 7.34e-19
C6875 VDD.n629 VSS 0.0036f
C6876 VDD.t382 VSS 0.00394f
C6877 VDD.n630 VSS 0.0036f
C6878 VDD.t370 VSS 0.00278f
C6879 VDD.n631 VSS 0.0018f
C6880 VDD.n632 VSS 0.00116f
C6881 VDD.n633 VSS 0.0018f
C6882 VDD.n634 VSS 3.27e-19
C6883 VDD.n635 VSS 5.58e-19
C6884 VDD.n636 VSS 4.56e-19
C6885 VDD.n637 VSS 0.00207f
C6886 VDD.n638 VSS 0.00196f
C6887 VDD.n639 VSS 5.1e-19
C6888 VDD.n640 VSS 6.12e-20
C6889 VDD.n641 VSS 4.9e-19
C6890 VDD.n642 VSS 2.87e-19
C6891 VDD.n643 VSS 0.00171f
C6892 VDD.n644 VSS 7.28e-19
C6893 VDD.t368 VSS 0.00321f
C6894 VDD.n645 VSS 0.00188f
C6895 VDD.n646 VSS 3.39e-19
C6896 VDD.n647 VSS 1.22e-19
C6897 VDD.n648 VSS 1.16e-19
C6898 VDD.n649 VSS 4.42e-19
C6899 VDD.n650 VSS 9.23e-19
C6900 VDD.n651 VSS 9.57e-19
C6901 VDD.n652 VSS 1.36e-19
C6902 VDD.n653 VSS 1.16e-19
C6903 VDD.n654 VSS 6.78e-20
C6904 VDD.n655 VSS 7.28e-19
C6905 VDD.n656 VSS 0.00154f
C6906 VDD.t376 VSS 0.00321f
C6907 VDD.n657 VSS 0.0024f
C6908 VDD.n658 VSS 3.27e-19
C6909 VDD.n659 VSS 9.53e-20
C6910 VDD.n660 VSS 0.0015f
C6911 VDD.n661 VSS 3.95e-19
C6912 VDD.n662 VSS 9.23e-19
C6913 VDD.n663 VSS 1.91e-19
C6914 VDD.n664 VSS 9.57e-19
C6915 VDD.n665 VSS 1.36e-19
C6916 VDD.n666 VSS 3.39e-19
C6917 VDD.n667 VSS 0.0012f
C6918 VDD.t364 VSS 0.00321f
C6919 VDD.n668 VSS 0.00274f
C6920 VDD.n669 VSS 8.56e-19
C6921 VDD.n670 VSS 7.28e-19
C6922 VDD.n671 VSS 6.78e-20
C6923 VDD.n672 VSS 1.16e-19
C6924 VDD.n673 VSS 1.36e-19
C6925 VDD.n674 VSS 9.57e-19
C6926 VDD.n675 VSS 1.91e-19
C6927 VDD.n676 VSS 9.23e-19
C6928 VDD.n677 VSS 2.86e-19
C6929 VDD.n678 VSS 0.0015f
C6930 VDD.n679 VSS 2.04e-19
C6931 VDD.n680 VSS 3.27e-19
C6932 VDD.n681 VSS 0.00308f
C6933 VDD.n682 VSS 7.28e-19
C6934 VDD.t574 VSS 0.00321f
C6935 VDD.n683 VSS 5.14e-19
C6936 VDD.n684 VSS 3.39e-19
C6937 VDD.n685 VSS 1.36e-19
C6938 VDD.n686 VSS 1.16e-19
C6939 VDD.n687 VSS 4.42e-19
C6940 VDD.n688 VSS 9.23e-19
C6941 VDD.n689 VSS 9.57e-19
C6942 VDD.n690 VSS 1.36e-19
C6943 VDD.n691 VSS 1.16e-19
C6944 VDD.n692 VSS 6.78e-20
C6945 VDD.n693 VSS 4.71e-19
C6946 VDD.t568 VSS 4.28e-19
C6947 VDD.n694 VSS 0.00347f
C6948 VDD.t572 VSS 3e-19
C6949 VDD.n695 VSS 0.00334f
C6950 VDD.n696 VSS 3.27e-19
C6951 VDD.n697 VSS 3.13e-19
C6952 VDD.n698 VSS 0.0015f
C6953 VDD.n699 VSS 1.77e-19
C6954 VDD.n700 VSS 9.23e-19
C6955 VDD.n701 VSS 1.91e-19
C6956 VDD.n702 VSS 9.57e-19
C6957 VDD.n703 VSS 1.36e-19
C6958 VDD.n704 VSS 3.39e-19
C6959 VDD.n705 VSS 0.00343f
C6960 VDD.t566 VSS 0.00321f
C6961 VDD.n706 VSS 5.14e-19
C6962 VDD.n707 VSS 0.00308f
C6963 VDD.n708 VSS 7.28e-19
C6964 VDD.n709 VSS 6.78e-20
C6965 VDD.n710 VSS 1.16e-19
C6966 VDD.n711 VSS 1.36e-19
C6967 VDD.n712 VSS 9.57e-19
C6968 VDD.n713 VSS 1.91e-19
C6969 VDD.n714 VSS 9.23e-19
C6970 VDD.n715 VSS 6.8e-20
C6971 VDD.n716 VSS 0.0015f
C6972 VDD.n717 VSS 4.22e-19
C6973 VDD.n718 VSS 3.27e-19
C6974 VDD.n719 VSS 8.56e-19
C6975 VDD.n720 VSS 7.28e-19
C6976 VDD.t576 VSS 0.00321f
C6977 VDD.n721 VSS 0.00274f
C6978 VDD.n722 VSS 3.39e-19
C6979 VDD.n723 VSS 1.36e-19
C6980 VDD.n724 VSS 1.16e-19
C6981 VDD.n725 VSS 4.42e-19
C6982 VDD.n726 VSS 9.23e-19
C6983 VDD.n727 VSS 1.8e-19
C6984 VDD.n728 VSS 8.84e-20
C6985 VDD.n729 VSS 1.91e-19
C6986 VDD.n730 VSS 9.57e-19
C6987 VDD.n731 VSS 9.53e-20
C6988 VDD.n732 VSS 1.16e-19
C6989 VDD.n733 VSS 6.78e-20
C6990 VDD.n734 VSS 7.28e-19
C6991 VDD.n735 VSS 0.00154f
C6992 VDD.n736 VSS 0.0036f
C6993 VDD.t596 VSS 0.00394f
C6994 VDD.n737 VSS 0.00565f
C6995 VDD.n738 VSS 6.94e-19
C6996 VDD.t597 VSS 0.00265f
C6997 VDD.n739 VSS 0.00443f
C6998 VDD.n740 VSS 4.49e-19
C6999 VDD.n741 VSS 0.00133f
C7000 VDD.n742 VSS 0.00207f
C7001 VDD.n743 VSS 0.00207f
C7002 VDD.n744 VSS 0.00207f
C7003 VDD.n745 VSS 8.71e-19
C7004 VDD.n746 VSS 0.00136f
C7005 VDD.n747 VSS 7.44e-19
C7006 VDD.n748 VSS 0.0036f
C7007 VDD.t598 VSS 0.00394f
C7008 VDD.n749 VSS 0.0036f
C7009 VDD.t600 VSS 0.00394f
C7010 VDD.n750 VSS 0.00274f
C7011 VDD.t660 VSS 0.00394f
C7012 VDD.n751 VSS 0.0036f
C7013 VDD.n752 VSS 7.34e-19
C7014 VDD.n753 VSS 6.6e-19
C7015 VDD.n754 VSS 7.35e-19
C7016 VDD.n755 VSS 0.00155f
C7017 VDD.n756 VSS 0.00155f
C7018 VDD.n757 VSS 9.19e-19
C7019 VDD.n758 VSS 7.34e-19
C7020 VDD.n759 VSS 0.00531f
C7021 VDD.t211 VSS 0.00394f
C7022 VDD.n760 VSS 0.00377f
C7023 VDD.t235 VSS 0.00394f
C7024 VDD.n761 VSS 0.00278f
C7025 VDD.n762 VSS 7.34e-19
C7026 VDD.n763 VSS 5.17e-19
C7027 VDD.n764 VSS 0.00155f
C7028 VDD.n765 VSS 0.0743f
C7029 VDD.n766 VSS 0.0111f
C7030 VDD.n767 VSS 0.0111f
C7031 VDD.n768 VSS 0.00191f
C7032 VDD.t607 VSS 5.37e-19
C7033 VDD.t605 VSS 5.37e-19
C7034 VDD.n769 VSS 0.00125f
C7035 VDD.n770 VSS 0.0036f
C7036 VDD.n771 VSS 7.55e-19
C7037 VDD.n772 VSS 7.55e-19
C7038 VDD.n773 VSS 7.34e-19
C7039 VDD.n774 VSS 7.34e-19
C7040 VDD.n775 VSS 0.00496f
C7041 VDD.t710 VSS 6.33e-19
C7042 VDD.t454 VSS 6.33e-19
C7043 VDD.n776 VSS 0.00145f
C7044 VDD.n777 VSS 0.00235f
C7045 VDD.n778 VSS 7.51e-19
C7046 VDD.t711 VSS 0.00404f
C7047 VDD.n779 VSS 7.59e-19
C7048 VDD.n780 VSS 6.38e-19
C7049 VDD.t712 VSS 6.33e-19
C7050 VDD.t714 VSS 6.33e-19
C7051 VDD.n781 VSS 0.00145f
C7052 VDD.n782 VSS 6.94e-19
C7053 VDD.n783 VSS 4.59e-19
C7054 VDD.t716 VSS 0.00251f
C7055 VDD.n784 VSS 0.00419f
C7056 VDD.n785 VSS 0.00365f
C7057 VDD.t715 VSS 0.0074f
C7058 VDD.n786 VSS 0.00795f
C7059 VDD.n787 VSS 9.97e-19
C7060 VDD.n788 VSS 0.013f
C7061 VDD.n789 VSS 0.00248f
C7062 VDD.n790 VSS 4.63e-19
C7063 VDD.n791 VSS 1.36e-19
C7064 VDD.n792 VSS 7.34e-19
C7065 VDD.n793 VSS 0.00225f
C7066 VDD.n794 VSS 0.00199f
C7067 VDD.n795 VSS 0.00155f
C7068 VDD.n796 VSS 0.00174f
C7069 VDD.n797 VSS 0.00459f
C7070 VDD.n798 VSS 5.98e-19
C7071 VDD.n799 VSS 0.00302f
C7072 VDD.n800 VSS 1.44e-19
C7073 VDD.n801 VSS 7.59e-19
C7074 VDD.n802 VSS 0.00365f
C7075 VDD.t713 VSS 0.00399f
C7076 VDD.n803 VSS 0.00365f
C7077 VDD.t709 VSS 0.00395f
C7078 VDD.n804 VSS 0.00278f
C7079 VDD.t453 VSS 0.00399f
C7080 VDD.n805 VSS 0.00365f
C7081 VDD.n806 VSS 7.51e-19
C7082 VDD.n807 VSS 7.74e-19
C7083 VDD.n808 VSS 0.00138f
C7084 VDD.n809 VSS 0.00291f
C7085 VDD.n810 VSS 0.00124f
C7086 VDD.n811 VSS 0.00164f
C7087 VDD.n812 VSS 0.00226f
C7088 VDD.n813 VSS 0.00187f
C7089 VDD.n814 VSS 4.59e-19
C7090 VDD.n815 VSS 1.36e-19
C7091 VDD.n816 VSS 7.55e-19
C7092 VDD.n817 VSS 0.00538f
C7093 VDD.t606 VSS 0.00399f
C7094 VDD.n818 VSS 0.00382f
C7095 VDD.t604 VSS 0.00399f
C7096 VDD.n819 VSS 0.00282f
C7097 VDD.n820 VSS 7.55e-19
C7098 VDD.n821 VSS 0.00147f
C7099 VDD.n822 VSS 0.00261f
C7100 VDD.n823 VSS 0.00207f
C7101 VDD.t63 VSS 0.0025f
C7102 VDD.n824 VSS 0.00282f
C7103 VDD.n825 VSS 7.34e-19
C7104 VDD.n826 VSS 3.67e-19
C7105 VDD.n827 VSS 4.97e-19
C7106 VDD.n828 VSS 9.59e-19
C7107 VDD.n829 VSS 9.46e-19
C7108 VDD.n830 VSS 2.59e-19
C7109 VDD.n831 VSS 3.27e-19
C7110 VDD.n832 VSS 7.34e-19
C7111 VDD.n833 VSS 7.77e-20
C7112 VDD.n834 VSS 4.15e-19
C7113 VDD.n835 VSS 9.35e-19
C7114 VDD.n836 VSS 9.46e-19
C7115 VDD.n837 VSS 3.39e-19
C7116 VDD.n838 VSS 0.00354f
C7117 VDD.n839 VSS 3.27e-19
C7118 VDD.n840 VSS 2.59e-19
C7119 VDD.n841 VSS 1.16e-19
C7120 VDD.n842 VSS 1.91e-19
C7121 VDD.n843 VSS 3.88e-19
C7122 VDD.n845 VSS 9.46e-19
C7123 VDD.n846 VSS 3.39e-19
C7124 VDD.n847 VSS 7.77e-20
C7125 VDD.n848 VSS 0.00112f
C7126 VDD.n849 VSS 3.27e-19
C7127 VDD.n850 VSS 4.42e-19
C7128 VDD.n851 VSS 1.16e-19
C7129 VDD.n852 VSS 1.91e-19
C7130 VDD.n853 VSS 1.16e-19
C7131 VDD.n854 VSS 9.46e-19
C7132 VDD.n855 VSS 6.78e-20
C7133 VDD.t400 VSS 0.00324f
C7134 VDD.n856 VSS 3.39e-19
C7135 VDD.n857 VSS 1.16e-19
C7136 VDD.n858 VSS 9.35e-19
C7137 VDD.n859 VSS 4.42e-19
C7138 VDD.n860 VSS 3.27e-19
C7139 VDD.n861 VSS 7.34e-19
C7140 VDD.n862 VSS 7.77e-20
C7141 VDD.n863 VSS 1.63e-19
C7142 VDD.n864 VSS 9.46e-19
C7143 VDD.n865 VSS 3.39e-19
C7144 VDD.n866 VSS 0.00328f
C7145 VDD.n867 VSS 3.27e-19
C7146 VDD.n868 VSS 4.42e-19
C7147 VDD.n869 VSS 1.16e-19
C7148 VDD.n870 VSS 1.91e-19
C7149 VDD.n871 VSS 1.16e-19
C7150 VDD.n872 VSS 9.46e-19
C7151 VDD.n873 VSS 6.78e-20
C7152 VDD.t637 VSS 0.00324f
C7153 VDD.n874 VSS 3.39e-19
C7154 VDD.n875 VSS 1.16e-19
C7155 VDD.n876 VSS 9.35e-19
C7156 VDD.n877 VSS 1.09e-19
C7157 VDD.n878 VSS 7.77e-20
C7158 VDD.n879 VSS 3.39e-19
C7159 VDD.n880 VSS 9.07e-19
C7160 VDD.n881 VSS 3.27e-19
C7161 VDD.n882 VSS 4.42e-19
C7162 VDD.n883 VSS 1.16e-19
C7163 VDD.n884 VSS 1.91e-19
C7164 VDD.n885 VSS 1.16e-19
C7165 VDD.n886 VSS 9.46e-19
C7166 VDD.n887 VSS 6.78e-20
C7167 VDD.t401 VSS 0.00324f
C7168 VDD.n888 VSS 3.39e-19
C7169 VDD.n889 VSS 1.16e-19
C7170 VDD.n890 VSS 9.35e-19
C7171 VDD.n891 VSS 4.42e-19
C7172 VDD.n892 VSS 3.27e-19
C7173 VDD.n893 VSS 7.34e-19
C7174 VDD.n894 VSS 6.78e-20
C7175 VDD.n895 VSS 1.16e-19
C7176 VDD.n896 VSS 4.49e-19
C7177 VDD.n897 VSS 1.16e-19
C7178 VDD.n898 VSS 1.91e-19
C7179 VDD.n899 VSS 1.16e-19
C7180 VDD.n900 VSS 3.39e-19
C7181 VDD.n901 VSS 0.00354f
C7182 VDD.n902 VSS 3.27e-19
C7183 VDD.n903 VSS 1.36e-19
C7184 VDD.n904 VSS 1.91e-19
C7185 VDD.n905 VSS 4.69e-19
C7186 VDD.n907 VSS 0.00207f
C7187 VDD.n908 VSS 0.00105f
C7188 VDD.n909 VSS 7.34e-19
C7189 VDD.n910 VSS 2.91e-19
C7190 VDD.n911 VSS 0.00535f
C7191 VDD.n912 VSS 7.34e-19
C7192 VDD.n913 VSS 0.00281f
C7193 VDD.t640 VSS 0.00176f
C7194 VDD.n914 VSS 0.00177f
C7195 VDD.n915 VSS 0.00207f
C7196 VDD.n916 VSS 0.0012f
C7197 VDD.n917 VSS 7.34e-19
C7198 VDD.t43 VSS 0.00397f
C7199 VDD.n918 VSS 7.44e-19
C7200 VDD.n919 VSS 0.00134f
C7201 VDD.n920 VSS 0.00101f
C7202 VDD.n921 VSS 7.34e-19
C7203 VDD.t608 VSS 0.00397f
C7204 VDD.n922 VSS 7.34e-19
C7205 VDD.n923 VSS 8.03e-19
C7206 VDD.n924 VSS 0.00207f
C7207 VDD.t652 VSS 9.52e-19
C7208 VDD.n925 VSS 0.00101f
C7209 VDD.n926 VSS 7.34e-19
C7210 VDD.t610 VSS 0.00397f
C7211 VDD.n927 VSS 7.34e-19
C7212 VDD.n928 VSS 0.0012f
C7213 VDD.n929 VSS 0.00207f
C7214 VDD.t251 VSS 3.84e-19
C7215 VDD.t500 VSS 3.65e-19
C7216 VDD.n930 VSS 8.01e-19
C7217 VDD.n931 VSS 7.89e-19
C7218 VDD.n932 VSS 7.34e-19
C7219 VDD.t666 VSS 0.00376f
C7220 VDD.n933 VSS 7.34e-19
C7221 VDD.n934 VSS 6.94e-19
C7222 VDD.n935 VSS 0.00207f
C7223 VDD.n936 VSS 0.00125f
C7224 VDD.n937 VSS 7.34e-19
C7225 VDD.t272 VSS 0.00397f
C7226 VDD.n938 VSS 7.34e-19
C7227 VDD.n939 VSS 0.00125f
C7228 VDD.n940 VSS 0.00207f
C7229 VDD.t249 VSS 3.84e-19
C7230 VDD.t132 VSS 3.84e-19
C7231 VDD.n941 VSS 8.11e-19
C7232 VDD.n942 VSS 0.0017f
C7233 VDD.n943 VSS 0.00137f
C7234 VDD.n944 VSS 7.44e-19
C7235 VDD.t659 VSS 0.00397f
C7236 VDD.n945 VSS 7.34e-19
C7237 VDD.n946 VSS 0.00105f
C7238 VDD.n947 VSS 0.00207f
C7239 VDD.n948 VSS 0.00281f
C7240 VDD.n949 VSS 7.34e-19
C7241 VDD.t129 VSS 0.00397f
C7242 VDD.n950 VSS 7.34e-19
C7243 VDD.n951 VSS 0.0012f
C7244 VDD.t130 VSS -3.41e-19
C7245 VDD.t456 VSS 6.16e-19
C7246 VDD.n952 VSS 0.00241f
C7247 VDD.n953 VSS 0.00164f
C7248 VDD.n954 VSS 0.00207f
C7249 VDD.t468 VSS -1.82e-19
C7250 VDD.t128 VSS 5.71e-19
C7251 VDD.n955 VSS 0.00268f
C7252 VDD.n956 VSS 0.00243f
C7253 VDD.n957 VSS 0.00134f
C7254 VDD.n958 VSS 7.44e-19
C7255 VDD.n959 VSS 7.34e-19
C7256 VDD.n960 VSS 0.00101f
C7257 VDD.n961 VSS 0.00207f
C7258 VDD.t56 VSS 4.05e-19
C7259 VDD.t549 VSS 4.05e-19
C7260 VDD.n962 VSS 8.77e-19
C7261 VDD.n963 VSS 8.03e-19
C7262 VDD.n964 VSS 7.34e-19
C7263 VDD.t655 VSS 0.00397f
C7264 VDD.n965 VSS 7.34e-19
C7265 VDD.n966 VSS 0.00101f
C7266 VDD.n967 VSS 0.00207f
C7267 VDD.n968 VSS 0.0012f
C7268 VDD.n969 VSS 7.34e-19
C7269 VDD.t516 VSS 0.00397f
C7270 VDD.n970 VSS 7.34e-19
C7271 VDD.n971 VSS 7.89e-19
C7272 VDD.n972 VSS 0.00207f
C7273 VDD.n973 VSS 6.94e-19
C7274 VDD.n974 VSS 7.34e-19
C7275 VDD.t447 VSS 0.00397f
C7276 VDD.n975 VSS 7.34e-19
C7277 VDD.n976 VSS 0.00125f
C7278 VDD.t448 VSS 0.00146f
C7279 VDD.t313 VSS 6.5e-19
C7280 VDD.n977 VSS 0.00234f
C7281 VDD.n978 VSS 0.00307f
C7282 VDD.n979 VSS 0.00207f
C7283 VDD.n980 VSS 0.00125f
C7284 VDD.n981 VSS 7.34e-19
C7285 VDD.t20 VSS 0.00397f
C7286 VDD.n982 VSS 7.44e-19
C7287 VDD.n983 VSS 0.00137f
C7288 VDD.n984 VSS 0.00207f
C7289 VDD.n985 VSS 0.00105f
C7290 VDD.n986 VSS 7.34e-19
C7291 VDD.n987 VSS 0.00535f
C7292 VDD.n988 VSS 7.34e-19
C7293 VDD.n989 VSS 0.00281f
C7294 VDD.t311 VSS 0.00176f
C7295 VDD.n990 VSS 0.00177f
C7296 VDD.n991 VSS 0.00207f
C7297 VDD.n992 VSS 0.0012f
C7298 VDD.n993 VSS 7.34e-19
C7299 VDD.t22 VSS 0.00397f
C7300 VDD.n994 VSS 7.44e-19
C7301 VDD.n995 VSS 0.00134f
C7302 VDD.n996 VSS 0.00101f
C7303 VDD.n997 VSS 7.34e-19
C7304 VDD.t254 VSS 0.00397f
C7305 VDD.n998 VSS 7.34e-19
C7306 VDD.n999 VSS 8.03e-19
C7307 VDD.n1000 VSS 0.00207f
C7308 VDD.t646 VSS 9.52e-19
C7309 VDD.n1001 VSS 0.00101f
C7310 VDD.n1002 VSS 7.34e-19
C7311 VDD.t252 VSS 0.00397f
C7312 VDD.n1003 VSS 7.34e-19
C7313 VDD.n1004 VSS 0.0012f
C7314 VDD.n1005 VSS 0.00207f
C7315 VDD.t84 VSS 3.84e-19
C7316 VDD.t342 VSS 3.65e-19
C7317 VDD.n1006 VSS 8.01e-19
C7318 VDD.n1007 VSS 7.89e-19
C7319 VDD.n1008 VSS 7.34e-19
C7320 VDD.t68 VSS 0.00376f
C7321 VDD.n1009 VSS 7.34e-19
C7322 VDD.n1010 VSS 6.94e-19
C7323 VDD.n1011 VSS 0.00207f
C7324 VDD.n1012 VSS 0.00125f
C7325 VDD.n1013 VSS 7.34e-19
C7326 VDD.t520 VSS 0.00397f
C7327 VDD.n1014 VSS 7.34e-19
C7328 VDD.n1015 VSS 0.00125f
C7329 VDD.n1016 VSS 0.00207f
C7330 VDD.t82 VSS 3.84e-19
C7331 VDD.t265 VSS 3.84e-19
C7332 VDD.n1017 VSS 8.11e-19
C7333 VDD.n1018 VSS 0.0017f
C7334 VDD.n1019 VSS 0.00137f
C7335 VDD.n1020 VSS 7.44e-19
C7336 VDD.t270 VSS 0.00397f
C7337 VDD.n1021 VSS 7.34e-19
C7338 VDD.n1022 VSS 0.00105f
C7339 VDD.n1023 VSS 0.00207f
C7340 VDD.n1024 VSS 0.00281f
C7341 VDD.n1025 VSS 7.34e-19
C7342 VDD.t266 VSS 0.00397f
C7343 VDD.n1026 VSS 7.34e-19
C7344 VDD.n1027 VSS 0.0012f
C7345 VDD.t267 VSS -3.41e-19
C7346 VDD.t50 VSS 6.16e-19
C7347 VDD.n1028 VSS 0.00241f
C7348 VDD.n1029 VSS 0.00164f
C7349 VDD.n1030 VSS 0.0065f
C7350 VDD.t642 VSS -1.82e-19
C7351 VDD.t269 VSS 5.71e-19
C7352 VDD.n1031 VSS 0.00268f
C7353 VDD.n1032 VSS 0.00243f
C7354 VDD.n1033 VSS 0.00134f
C7355 VDD.n1034 VSS 7.44e-19
C7356 VDD.n1035 VSS 0.00118f
C7357 VDD.n1036 VSS 0.00922f
C7358 VDD.t641 VSS 0.00455f
C7359 VDD.n1037 VSS 0.0041f
C7360 VDD.t268 VSS 0.00397f
C7361 VDD.n1038 VSS 0.00635f
C7362 VDD.n1039 VSS 0.00574f
C7363 VDD.n1040 VSS 7.34e-19
C7364 VDD.n1041 VSS 0.00109f
C7365 VDD.n1042 VSS 0.00207f
C7366 VDD.n1043 VSS 0.00207f
C7367 VDD.n1044 VSS 0.00207f
C7368 VDD.n1045 VSS 0.00125f
C7369 VDD.n1046 VSS 7.34e-19
C7370 VDD.n1047 VSS 0.00419f
C7371 VDD.t49 VSS 0.00397f
C7372 VDD.n1048 VSS 0.00535f
C7373 VDD.n1049 VSS 0.00311f
C7374 VDD.t594 VSS 0.00397f
C7375 VDD.n1050 VSS 0.00717f
C7376 VDD.n1051 VSS 7.34e-19
C7377 VDD.t595 VSS 0.00176f
C7378 VDD.n1052 VSS 0.00177f
C7379 VDD.n1053 VSS 0.00195f
C7380 VDD.n1054 VSS 0.00207f
C7381 VDD.n1055 VSS 0.00207f
C7382 VDD.n1056 VSS 0.00207f
C7383 VDD.n1057 VSS 0.0011f
C7384 VDD.n1058 VSS 7.34e-19
C7385 VDD.n1059 VSS 0.00414f
C7386 VDD.t81 VSS 0.00397f
C7387 VDD.n1060 VSS 0.00466f
C7388 VDD.t264 VSS 0.00397f
C7389 VDD.n1061 VSS 0.00432f
C7390 VDD.n1062 VSS 0.00475f
C7391 VDD.n1063 VSS 7.34e-19
C7392 VDD.n1064 VSS 8.91e-19
C7393 VDD.n1065 VSS 0.00207f
C7394 VDD.n1066 VSS 0.00207f
C7395 VDD.n1067 VSS 0.00207f
C7396 VDD.n1068 VSS 0.00125f
C7397 VDD.n1069 VSS 7.34e-19
C7398 VDD.t253 VSS 0.0076f
C7399 VDD.n1070 VSS 0.00622f
C7400 VDD.t343 VSS 0.00397f
C7401 VDD.t592 VSS 0.00384f
C7402 VDD.n1071 VSS 0.00419f
C7403 VDD.n1072 VSS 0.0057f
C7404 VDD.n1073 VSS 7.34e-19
C7405 VDD.t344 VSS 0.00146f
C7406 VDD.t593 VSS 6.5e-19
C7407 VDD.n1074 VSS 0.00234f
C7408 VDD.n1075 VSS 0.00307f
C7409 VDD.n1076 VSS 7.35e-19
C7410 VDD.n1077 VSS 0.00207f
C7411 VDD.n1078 VSS 0.00207f
C7412 VDD.n1079 VSS 0.00207f
C7413 VDD.n1080 VSS 0.00125f
C7414 VDD.n1081 VSS 7.34e-19
C7415 VDD.n1082 VSS 0.0041f
C7416 VDD.n1083 VSS 0.00453f
C7417 VDD.t83 VSS 0.00397f
C7418 VDD.n1084 VSS 0.00518f
C7419 VDD.t341 VSS 0.00397f
C7420 VDD.n1085 VSS 0.00458f
C7421 VDD.n1086 VSS 7.44e-19
C7422 VDD.n1087 VSS 0.00137f
C7423 VDD.n1088 VSS 0.00187f
C7424 VDD.n1089 VSS 0.00207f
C7425 VDD.n1090 VSS 0.00207f
C7426 VDD.n1091 VSS 0.00207f
C7427 VDD.n1092 VSS 0.00125f
C7428 VDD.n1093 VSS 7.34e-19
C7429 VDD.n1094 VSS 0.00363f
C7430 VDD.t521 VSS 0.00397f
C7431 VDD.n1095 VSS 0.00401f
C7432 VDD.t645 VSS 0.00397f
C7433 VDD.n1096 VSS 0.00622f
C7434 VDD.n1097 VSS 0.00587f
C7435 VDD.n1098 VSS 7.44e-19
C7436 VDD.n1099 VSS 0.00136f
C7437 VDD.n1100 VSS 0.00207f
C7438 VDD.n1101 VSS 0.00207f
C7439 VDD.n1102 VSS 0.00207f
C7440 VDD.n1103 VSS 0.00122f
C7441 VDD.n1104 VSS 0.00207f
C7442 VDD.t255 VSS 4.05e-19
C7443 VDD.t523 VSS 4.05e-19
C7444 VDD.n1105 VSS 8.77e-19
C7445 VDD.n1106 VSS 0.00182f
C7446 VDD.n1107 VSS 0.00136f
C7447 VDD.n1108 VSS 7.44e-19
C7448 VDD.n1109 VSS 0.00363f
C7449 VDD.t522 VSS 0.00393f
C7450 VDD.n1110 VSS 7.34e-19
C7451 VDD.n1111 VSS 0.0041f
C7452 VDD.t664 VSS 0.00397f
C7453 VDD.n1112 VSS 0.00535f
C7454 VDD.n1113 VSS 7.34e-19
C7455 VDD.n1114 VSS 0.00101f
C7456 VDD.n1115 VSS 0.00155f
C7457 VDD.t665 VSS -1.82e-19
C7458 VDD.t23 VSS 5.71e-19
C7459 VDD.n1116 VSS 0.00268f
C7460 VDD.n1117 VSS 0.00243f
C7461 VDD.n1118 VSS 0.00207f
C7462 VDD.n1119 VSS 0.00207f
C7463 VDD.n1120 VSS 0.00109f
C7464 VDD.n1121 VSS 7.34e-19
C7465 VDD.n1122 VSS 0.00574f
C7466 VDD.n1123 VSS 0.00635f
C7467 VDD.t24 VSS 0.00397f
C7468 VDD.t296 VSS 0.00397f
C7469 VDD.n1124 VSS 0.00419f
C7470 VDD.n1125 VSS 7.34e-19
C7471 VDD.t25 VSS -3.41e-19
C7472 VDD.t297 VSS 6.16e-19
C7473 VDD.n1126 VSS 0.00241f
C7474 VDD.n1127 VSS 0.00164f
C7475 VDD.n1128 VSS 0.00125f
C7476 VDD.n1129 VSS 0.00207f
C7477 VDD.n1130 VSS 0.00207f
C7478 VDD.n1131 VSS 0.00207f
C7479 VDD.n1132 VSS 0.00195f
C7480 VDD.n1133 VSS 7.34e-19
C7481 VDD.n1134 VSS 0.00717f
C7482 VDD.t310 VSS 0.00397f
C7483 VDD.n1135 VSS 0.00311f
C7484 VDD.t321 VSS 0.00397f
C7485 VDD.n1136 VSS 0.00466f
C7486 VDD.t514 VSS 0.00397f
C7487 VDD.n1137 VSS 0.00414f
C7488 VDD.n1138 VSS 7.34e-19
C7489 VDD.n1139 VSS 0.0011f
C7490 VDD.n1140 VSS 0.00207f
C7491 VDD.t515 VSS 3.84e-19
C7492 VDD.t21 VSS 3.84e-19
C7493 VDD.n1141 VSS 8.11e-19
C7494 VDD.n1142 VSS 0.0017f
C7495 VDD.n1143 VSS 0.00207f
C7496 VDD.n1144 VSS 0.00207f
C7497 VDD.n1145 VSS 8.91e-19
C7498 VDD.n1146 VSS 7.34e-19
C7499 VDD.n1147 VSS 0.00475f
C7500 VDD.n1148 VSS 0.00432f
C7501 VDD.t700 VSS 0.00397f
C7502 VDD.n1149 VSS 0.00622f
C7503 VDD.t54 VSS 0.0076f
C7504 VDD.n1150 VSS 7.34e-19
C7505 VDD.n1151 VSS 0.00125f
C7506 VDD.n1152 VSS 0.00207f
C7507 VDD.n1153 VSS 0.00207f
C7508 VDD.n1154 VSS 0.00207f
C7509 VDD.n1155 VSS 7.35e-19
C7510 VDD.n1156 VSS 7.34e-19
C7511 VDD.n1157 VSS 0.0057f
C7512 VDD.n1158 VSS 0.00419f
C7513 VDD.t312 VSS 0.00384f
C7514 VDD.t11 VSS 0.00376f
C7515 VDD.n1159 VSS 0.00453f
C7516 VDD.n1160 VSS 0.0041f
C7517 VDD.n1161 VSS 7.34e-19
C7518 VDD.n1162 VSS 0.00125f
C7519 VDD.n1163 VSS 0.00207f
C7520 VDD.n1164 VSS 0.00207f
C7521 VDD.n1165 VSS 0.00207f
C7522 VDD.t517 VSS 3.84e-19
C7523 VDD.t446 VSS 3.65e-19
C7524 VDD.n1166 VSS 8.01e-19
C7525 VDD.n1167 VSS 0.00187f
C7526 VDD.n1168 VSS 0.00137f
C7527 VDD.n1169 VSS 7.44e-19
C7528 VDD.n1170 VSS 0.00458f
C7529 VDD.t445 VSS 0.00397f
C7530 VDD.n1171 VSS 0.00518f
C7531 VDD.t53 VSS 0.00397f
C7532 VDD.n1172 VSS 0.00401f
C7533 VDD.t699 VSS 0.00397f
C7534 VDD.n1173 VSS 0.00363f
C7535 VDD.n1174 VSS 7.34e-19
C7536 VDD.n1175 VSS 0.00125f
C7537 VDD.n1176 VSS 0.00207f
C7538 VDD.n1177 VSS 0.00207f
C7539 VDD.n1178 VSS 0.00207f
C7540 VDD.t656 VSS 9.52e-19
C7541 VDD.n1179 VSS 0.00207f
C7542 VDD.n1180 VSS 0.00136f
C7543 VDD.n1181 VSS 7.44e-19
C7544 VDD.n1182 VSS 0.00587f
C7545 VDD.n1183 VSS 0.00622f
C7546 VDD.t55 VSS 0.00397f
C7547 VDD.n1184 VSS 7.34e-19
C7548 VDD.t548 VSS 0.00393f
C7549 VDD.n1185 VSS 0.00363f
C7550 VDD.n1186 VSS 7.44e-19
C7551 VDD.n1187 VSS 0.00136f
C7552 VDD.n1188 VSS 0.00182f
C7553 VDD.n1189 VSS 0.00207f
C7554 VDD.n1190 VSS 0.00122f
C7555 VDD.n1191 VSS 0.00155f
C7556 VDD.n1192 VSS 0.00101f
C7557 VDD.n1193 VSS 7.34e-19
C7558 VDD.n1194 VSS 0.00535f
C7559 VDD.t467 VSS 0.00397f
C7560 VDD.n1195 VSS 0.0041f
C7561 VDD.t127 VSS 0.00397f
C7562 VDD.n1196 VSS 0.00635f
C7563 VDD.n1197 VSS 0.00574f
C7564 VDD.n1198 VSS 7.34e-19
C7565 VDD.n1199 VSS 0.00109f
C7566 VDD.n1200 VSS 0.00207f
C7567 VDD.n1201 VSS 0.00207f
C7568 VDD.n1202 VSS 0.00207f
C7569 VDD.n1203 VSS 0.00125f
C7570 VDD.n1204 VSS 7.34e-19
C7571 VDD.n1205 VSS 0.00419f
C7572 VDD.t455 VSS 0.00397f
C7573 VDD.n1206 VSS 0.00535f
C7574 VDD.n1207 VSS 0.00311f
C7575 VDD.t621 VSS 0.00397f
C7576 VDD.n1208 VSS 0.00717f
C7577 VDD.n1209 VSS 7.34e-19
C7578 VDD.t622 VSS 0.00176f
C7579 VDD.n1210 VSS 0.00177f
C7580 VDD.n1211 VSS 0.00195f
C7581 VDD.n1212 VSS 0.00207f
C7582 VDD.n1213 VSS 0.00207f
C7583 VDD.n1214 VSS 0.00207f
C7584 VDD.n1215 VSS 0.0011f
C7585 VDD.n1216 VSS 7.34e-19
C7586 VDD.n1217 VSS 0.00414f
C7587 VDD.t248 VSS 0.00397f
C7588 VDD.n1218 VSS 0.00466f
C7589 VDD.t131 VSS 0.00397f
C7590 VDD.n1219 VSS 0.00432f
C7591 VDD.n1220 VSS 0.00475f
C7592 VDD.n1221 VSS 7.34e-19
C7593 VDD.n1222 VSS 8.91e-19
C7594 VDD.n1223 VSS 0.00207f
C7595 VDD.n1224 VSS 0.00207f
C7596 VDD.n1225 VSS 0.00207f
C7597 VDD.n1226 VSS 0.00125f
C7598 VDD.n1227 VSS 7.34e-19
C7599 VDD.t611 VSS 0.0076f
C7600 VDD.n1228 VSS 0.00622f
C7601 VDD.t497 VSS 0.00397f
C7602 VDD.t619 VSS 0.00384f
C7603 VDD.n1229 VSS 0.00419f
C7604 VDD.n1230 VSS 0.0057f
C7605 VDD.n1231 VSS 7.34e-19
C7606 VDD.t498 VSS 0.00146f
C7607 VDD.t620 VSS 6.5e-19
C7608 VDD.n1232 VSS 0.00234f
C7609 VDD.n1233 VSS 0.00307f
C7610 VDD.n1234 VSS 7.35e-19
C7611 VDD.n1235 VSS 0.00207f
C7612 VDD.n1236 VSS 0.00207f
C7613 VDD.n1237 VSS 0.00207f
C7614 VDD.n1238 VSS 0.00125f
C7615 VDD.n1239 VSS 7.34e-19
C7616 VDD.n1240 VSS 0.0041f
C7617 VDD.n1241 VSS 0.00453f
C7618 VDD.t250 VSS 0.00397f
C7619 VDD.n1242 VSS 0.00518f
C7620 VDD.t499 VSS 0.00397f
C7621 VDD.n1243 VSS 0.00458f
C7622 VDD.n1244 VSS 7.44e-19
C7623 VDD.n1245 VSS 0.00137f
C7624 VDD.n1246 VSS 0.00187f
C7625 VDD.n1247 VSS 0.00207f
C7626 VDD.n1248 VSS 0.00207f
C7627 VDD.n1249 VSS 0.00207f
C7628 VDD.n1250 VSS 0.00125f
C7629 VDD.n1251 VSS 7.34e-19
C7630 VDD.n1252 VSS 0.00363f
C7631 VDD.t271 VSS 0.00397f
C7632 VDD.n1253 VSS 0.00401f
C7633 VDD.t651 VSS 0.00397f
C7634 VDD.n1254 VSS 0.00622f
C7635 VDD.n1255 VSS 0.00587f
C7636 VDD.n1256 VSS 7.44e-19
C7637 VDD.n1257 VSS 0.00136f
C7638 VDD.n1258 VSS 0.00207f
C7639 VDD.n1259 VSS 0.00207f
C7640 VDD.n1260 VSS 0.00207f
C7641 VDD.n1261 VSS 0.00122f
C7642 VDD.n1262 VSS 0.00207f
C7643 VDD.t609 VSS 4.05e-19
C7644 VDD.t10 VSS 4.05e-19
C7645 VDD.n1263 VSS 8.77e-19
C7646 VDD.n1264 VSS 0.00182f
C7647 VDD.n1265 VSS 0.00136f
C7648 VDD.n1266 VSS 7.44e-19
C7649 VDD.n1267 VSS 0.00363f
C7650 VDD.t9 VSS 0.00393f
C7651 VDD.n1268 VSS 7.34e-19
C7652 VDD.n1269 VSS 0.0041f
C7653 VDD.t58 VSS 0.00397f
C7654 VDD.n1270 VSS 0.00535f
C7655 VDD.n1271 VSS 7.34e-19
C7656 VDD.n1272 VSS 0.00101f
C7657 VDD.n1273 VSS 0.00155f
C7658 VDD.t59 VSS -1.82e-19
C7659 VDD.t44 VSS 5.71e-19
C7660 VDD.n1274 VSS 0.00268f
C7661 VDD.n1275 VSS 0.00243f
C7662 VDD.n1276 VSS 0.00207f
C7663 VDD.n1277 VSS 0.00207f
C7664 VDD.n1278 VSS 0.00109f
C7665 VDD.n1279 VSS 7.34e-19
C7666 VDD.n1280 VSS 0.00574f
C7667 VDD.n1281 VSS 0.00635f
C7668 VDD.t45 VSS 0.00397f
C7669 VDD.t449 VSS 0.00397f
C7670 VDD.n1282 VSS 0.00419f
C7671 VDD.n1283 VSS 7.34e-19
C7672 VDD.t46 VSS -3.41e-19
C7673 VDD.t450 VSS 6.16e-19
C7674 VDD.n1284 VSS 0.00241f
C7675 VDD.n1285 VSS 0.00164f
C7676 VDD.n1286 VSS 0.00125f
C7677 VDD.n1287 VSS 0.00207f
C7678 VDD.n1288 VSS 0.00207f
C7679 VDD.n1289 VSS 0.00207f
C7680 VDD.n1290 VSS 0.00195f
C7681 VDD.n1291 VSS 7.34e-19
C7682 VDD.n1292 VSS 0.00717f
C7683 VDD.t639 VSS 0.00397f
C7684 VDD.n1293 VSS 0.00311f
C7685 VDD.t740 VSS 0.00397f
C7686 VDD.n1294 VSS 3.39e-19
C7687 VDD.n1295 VSS 0.00367f
C7688 VDD.n1296 VSS 7.77e-20
C7689 VDD.n1297 VSS 7.34e-19
C7690 VDD.n1298 VSS 6.48e-19
C7691 VDD.t669 VSS 0.00285f
C7692 VDD.n1299 VSS 0.00414f
C7693 VDD.n1300 VSS 6.3e-19
C7694 VDD.n1301 VSS 0.00108f
C7695 VDD.n1302 VSS 0.00197f
C7696 VDD.n1303 VSS 0.00104f
C7697 VDD.t670 VSS 3.84e-19
C7698 VDD.t48 VSS 3.84e-19
C7699 VDD.n1304 VSS 8.07e-19
C7700 VDD.n1305 VSS 0.0017f
C7701 VDD.n1306 VSS 7.48e-19
C7702 VDD.n1307 VSS 9.35e-19
C7703 VDD.n1308 VSS 9.46e-19
C7704 VDD.n1309 VSS 1.29e-19
C7705 VDD.n1310 VSS 1.16e-19
C7706 VDD.n1311 VSS 6.78e-20
C7707 VDD.n1312 VSS 3.45e-19
C7708 VDD.t47 VSS 4.32e-19
C7709 VDD.n1313 VSS 0.00363f
C7710 VDD.n1314 VSS 0.00354f
C7711 VDD.n1315 VSS 3.27e-19
C7712 VDD.n1316 VSS 4.42e-19
C7713 VDD.n1317 VSS 4.49e-19
C7714 VDD.n1318 VSS 9.35e-19
C7715 VDD.n1319 VSS 1.91e-19
C7716 VDD.n1320 VSS 9.46e-19
C7717 VDD.n1321 VSS 1.29e-19
C7718 VDD.n1322 VSS 3.39e-19
C7719 VDD.n1323 VSS 0.00117f
C7720 VDD.t350 VSS 0.00324f
C7721 VDD.n1324 VSS 0.00281f
C7722 VDD.n1325 VSS 8.2e-19
C7723 VDD.n1326 VSS 7.34e-19
C7724 VDD.n1327 VSS 6.78e-20
C7725 VDD.n1328 VSS 1.16e-19
C7726 VDD.n1329 VSS 1.29e-19
C7727 VDD.n1330 VSS 9.46e-19
C7728 VDD.n1331 VSS 1.91e-19
C7729 VDD.n1332 VSS 9.35e-19
C7730 VDD.n1333 VSS 4.49e-19
C7731 VDD.n1334 VSS 4.42e-19
C7732 VDD.n1335 VSS 3.27e-19
C7733 VDD.n1336 VSS 0.00315f
C7734 VDD.n1337 VSS 7.34e-19
C7735 VDD.t77 VSS 0.00324f
C7736 VDD.n1338 VSS 0.00306f
C7737 VDD.n1339 VSS 3.39e-19
C7738 VDD.n1340 VSS 1.29e-19
C7739 VDD.n1341 VSS 1.16e-19
C7740 VDD.n1342 VSS 4.49e-19
C7741 VDD.n1343 VSS 9.35e-19
C7742 VDD.n1344 VSS 1.91e-19
C7743 VDD.n1345 VSS 9.46e-19
C7744 VDD.n1346 VSS 1.29e-19
C7745 VDD.n1347 VSS 1.16e-19
C7746 VDD.n1348 VSS 6.78e-20
C7747 VDD.n1349 VSS 7.34e-19
C7748 VDD.n1350 VSS 0.00367f
C7749 VDD.n1351 VSS 0.00104f
C7750 VDD.n1352 VSS 7.34e-19
C7751 VDD.n1353 VSS 0.00354f
C7752 VDD.n1354 VSS 3.27e-19
C7753 VDD.t78 VSS 0.00146f
C7754 VDD.t638 VSS 6.5e-19
C7755 VDD.n1356 VSS 0.00234f
C7756 VDD.n1357 VSS 0.00294f
C7757 VDD.n1358 VSS 6.8e-20
C7758 VDD.n1359 VSS 9.46e-19
C7759 VDD.n1360 VSS 1.91e-19
C7760 VDD.n1361 VSS 9.35e-19
C7761 VDD.n1362 VSS 4.49e-19
C7762 VDD.n1363 VSS 4.42e-19
C7763 VDD.n1364 VSS 3.27e-19
C7764 VDD.n1365 VSS 0.00294f
C7765 VDD.n1366 VSS 7.34e-19
C7766 VDD.t624 VSS 0.00324f
C7767 VDD.n1367 VSS 6.91e-19
C7768 VDD.n1368 VSS 3.39e-19
C7769 VDD.n1369 VSS 1.29e-19
C7770 VDD.n1370 VSS 1.16e-19
C7771 VDD.n1371 VSS 4.49e-19
C7772 VDD.n1372 VSS 9.35e-19
C7773 VDD.n1373 VSS 9.35e-19
C7774 VDD.n1374 VSS 1.91e-19
C7775 VDD.n1375 VSS 9.46e-19
C7776 VDD.n1376 VSS 1.29e-19
C7777 VDD.n1377 VSS 1.16e-19
C7778 VDD.n1378 VSS 6.78e-20
C7779 VDD.n1379 VSS 7.34e-19
C7780 VDD.n1380 VSS 0.00138f
C7781 VDD.t667 VSS 0.00324f
C7782 VDD.n1381 VSS 0.00259f
C7783 VDD.n1382 VSS 3.27e-19
C7784 VDD.t668 VSS 3.84e-19
C7785 VDD.t76 VSS 3.65e-19
C7786 VDD.n1383 VSS 7.97e-19
C7787 VDD.n1384 VSS 1.91e-19
C7788 VDD.n1385 VSS 0.00187f
C7789 VDD.n1386 VSS 0.00114f
C7790 VDD.n1388 VSS 3.39e-19
C7791 VDD.n1389 VSS 0.00199f
C7792 VDD.t75 VSS 0.00324f
C7793 VDD.n1390 VSS 0.00199f
C7794 VDD.n1391 VSS 0.00319f
C7795 VDD.n1392 VSS 7.34e-19
C7796 VDD.n1393 VSS 6.78e-20
C7797 VDD.n1394 VSS 1.16e-19
C7798 VDD.n1395 VSS 1.29e-19
C7799 VDD.n1396 VSS 9.46e-19
C7800 VDD.n1397 VSS 1.91e-19
C7801 VDD.n1398 VSS 9.35e-19
C7802 VDD.n1399 VSS 4.49e-19
C7803 VDD.n1400 VSS 4.42e-19
C7804 VDD.n1401 VSS 3.27e-19
C7805 VDD.n1402 VSS 7.77e-19
C7806 VDD.n1403 VSS 7.34e-19
C7807 VDD.t349 VSS 0.00324f
C7808 VDD.n1404 VSS 0.00285f
C7809 VDD.n1405 VSS 3.39e-19
C7810 VDD.n1406 VSS 1.29e-19
C7811 VDD.n1407 VSS 1.16e-19
C7812 VDD.n1408 VSS 4.49e-19
C7813 VDD.n1409 VSS 9.35e-19
C7814 VDD.n1410 VSS 9.35e-19
C7815 VDD.n1411 VSS 1.91e-19
C7816 VDD.n1412 VSS 9.46e-19
C7817 VDD.n1413 VSS 1.29e-19
C7818 VDD.n1414 VSS 1.16e-19
C7819 VDD.n1415 VSS 6.78e-20
C7820 VDD.n1416 VSS 7.34e-19
C7821 VDD.n1417 VSS 0.00289f
C7822 VDD.t580 VSS 0.00324f
C7823 VDD.n1418 VSS 3.39e-19
C7824 VDD.n1419 VSS 0.00367f
C7825 VDD.n1420 VSS 7.34e-19
C7826 VDD.n1421 VSS 0.00108f
C7827 VDD.n1422 VSS 3.27e-19
C7828 VDD.t581 VSS 9.48e-19
C7829 VDD.n1423 VSS 0.00207f
C7830 VDD.n1424 VSS 0.00113f
C7831 VDD.n1425 VSS 9.35e-19
C7832 VDD.n1426 VSS 9.35e-19
C7833 VDD.n1427 VSS 1.91e-19
C7834 VDD.n1428 VSS 9.46e-19
C7835 VDD.n1429 VSS 1.29e-19
C7836 VDD.n1430 VSS 1.16e-19
C7837 VDD.n1431 VSS 6.78e-20
C7838 VDD.n1432 VSS 7.34e-19
C7839 VDD.n1433 VSS 0.00306f
C7840 VDD.t398 VSS 0.00324f
C7841 VDD.n1434 VSS 9.07e-19
C7842 VDD.n1435 VSS 3.27e-19
C7843 VDD.t399 VSS 4.05e-19
C7844 VDD.t579 VSS 4.05e-19
C7845 VDD.n1436 VSS 8.73e-19
C7846 VDD.n1437 VSS 1.91e-19
C7847 VDD.n1438 VSS 0.00182f
C7848 VDD.n1439 VSS 0.00113f
C7849 VDD.n1441 VSS 3.39e-19
C7850 VDD.n1442 VSS 0.00272f
C7851 VDD.t578 VSS 0.00324f
C7852 VDD.n1443 VSS 0.00125f
C7853 VDD.n1444 VSS 7.77e-19
C7854 VDD.n1445 VSS 7.34e-19
C7855 VDD.n1446 VSS 6.78e-20
C7856 VDD.n1447 VSS 1.16e-19
C7857 VDD.n1448 VSS 1.29e-19
C7858 VDD.n1449 VSS 1.16e-19
C7859 VDD.n1450 VSS 1.91e-19
C7860 VDD.n1451 VSS 1.8e-19
C7861 VDD.n1452 VSS 0.00134f
C7862 VDD.n1453 VSS 0.00107f
C7863 VDD.n1454 VSS 6.94e-19
C7864 VDD.n1455 VSS 0.00643f
C7865 VDD.n1456 VSS 0.0041f
C7866 VDD.t62 VSS 0.00397f
C7867 VDD.n1457 VSS 0.00458f
C7868 VDD.n1458 VSS 7.34e-19
C7869 VDD.n1459 VSS 9.19e-19
C7870 VDD.n1460 VSS 0.00123f
C7871 VDD.n1461 VSS 0.0283f
C7872 VDD.n1462 VSS 0.00207f
C7873 VDD.t587 VSS 5.71e-19
C7874 VDD.t678 VSS -1.82e-19
C7875 VDD.n1463 VSS 0.00268f
C7876 VDD.n1464 VSS 0.00243f
C7877 VDD.n1465 VSS 0.00134f
C7878 VDD.n1466 VSS 7.44e-19
C7879 VDD.n1467 VSS 0.00621f
C7880 VDD.n1468 VSS 7.34e-19
C7881 VDD.n1469 VSS 0.0012f
C7882 VDD.n1470 VSS 0.00207f
C7883 VDD.t426 VSS 6.16e-19
C7884 VDD.t589 VSS -3.41e-19
C7885 VDD.n1471 VSS 0.00241f
C7886 VDD.n1472 VSS 0.00164f
C7887 VDD.n1473 VSS 7.34e-19
C7888 VDD.t485 VSS 0.00389f
C7889 VDD.n1474 VSS 7.34e-19
C7890 VDD.t486 VSS 0.00176f
C7891 VDD.n1475 VSS 0.00177f
C7892 VDD.n1476 VSS 0.00281f
C7893 VDD.n1477 VSS 0.00207f
C7894 VDD.n1478 VSS 0.00137f
C7895 VDD.n1479 VSS 7.44e-19
C7896 VDD.n1480 VSS 0.00422f
C7897 VDD.n1481 VSS 7.34e-19
C7898 VDD.n1482 VSS 0.00125f
C7899 VDD.n1483 VSS 0.00207f
C7900 VDD.n1484 VSS 0.00125f
C7901 VDD.n1485 VSS 7.34e-19
C7902 VDD.n1486 VSS 0.0041f
C7903 VDD.n1487 VSS 7.34e-19
C7904 VDD.t488 VSS 6.5e-19
C7905 VDD.t244 VSS 0.00146f
C7906 VDD.n1488 VSS 0.00234f
C7907 VDD.n1489 VSS 0.00307f
C7908 VDD.n1490 VSS 0.00207f
C7909 VDD.n1491 VSS 7.89e-19
C7910 VDD.n1492 VSS 7.34e-19
C7911 VDD.t245 VSS 0.00389f
C7912 VDD.n1493 VSS 7.34e-19
C7913 VDD.n1494 VSS 0.0012f
C7914 VDD.n1495 VSS 0.00207f
C7915 VDD.n1496 VSS 0.00101f
C7916 VDD.n1497 VSS 7.34e-19
C7917 VDD.n1498 VSS 0.00608f
C7918 VDD.n1499 VSS 7.34e-19
C7919 VDD.n1500 VSS 8.03e-19
C7920 VDD.t632 VSS 4.05e-19
C7921 VDD.t532 VSS 4.05e-19
C7922 VDD.n1501 VSS 8.77e-19
C7923 VDD.n1502 VSS 0.00101f
C7924 VDD.n1503 VSS 7.34e-19
C7925 VDD.t741 VSS 0.00389f
C7926 VDD.n1504 VSS 7.44e-19
C7927 VDD.n1505 VSS 0.00134f
C7928 VDD.n1506 VSS 0.00207f
C7929 VDD.n1507 VSS 0.0012f
C7930 VDD.n1508 VSS 7.34e-19
C7931 VDD.t423 VSS 0.00389f
C7932 VDD.n1509 VSS 7.34e-19
C7933 VDD.t424 VSS 6.16e-19
C7934 VDD.t32 VSS -3.41e-19
C7935 VDD.n1510 VSS 0.00241f
C7936 VDD.n1511 VSS 0.00164f
C7937 VDD.n1512 VSS 0.00207f
C7938 VDD.t92 VSS 0.00176f
C7939 VDD.n1513 VSS 0.00177f
C7940 VDD.n1514 VSS 7.34e-19
C7941 VDD.t386 VSS 0.00389f
C7942 VDD.n1515 VSS 7.44e-19
C7943 VDD.n1516 VSS 0.00137f
C7944 VDD.n1517 VSS 0.00105f
C7945 VDD.n1518 VSS 0.00207f
C7946 VDD.n1519 VSS 0.00125f
C7947 VDD.n1520 VSS 7.34e-19
C7948 VDD.n1521 VSS 0.00608f
C7949 VDD.n1522 VSS 7.34e-19
C7950 VDD.n1523 VSS 0.00125f
C7951 VDD.n1524 VSS 0.00207f
C7952 VDD.t90 VSS 6.5e-19
C7953 VDD.t122 VSS 0.00146f
C7954 VDD.n1525 VSS 0.00234f
C7955 VDD.n1526 VSS 0.00307f
C7956 VDD.n1527 VSS 7.34e-19
C7957 VDD.n1528 VSS 0.00443f
C7958 VDD.n1529 VSS 7.34e-19
C7959 VDD.n1530 VSS 7.89e-19
C7960 VDD.n1531 VSS 6.94e-19
C7961 VDD.n1532 VSS 0.00207f
C7962 VDD.t120 VSS 3.65e-19
C7963 VDD.t385 VSS 3.84e-19
C7964 VDD.n1533 VSS 8.01e-19
C7965 VDD.n1534 VSS 0.0012f
C7966 VDD.n1535 VSS 7.34e-19
C7967 VDD.t200 VSS 0.00389f
C7968 VDD.n1536 VSS 7.34e-19
C7969 VDD.n1537 VSS 0.00101f
C7970 VDD.n1538 VSS 0.00207f
C7971 VDD.t644 VSS 9.52e-19
C7972 VDD.n1539 VSS 8.03e-19
C7973 VDD.n1540 VSS 7.34e-19
C7974 VDD.t409 VSS 0.00313f
C7975 VDD.n1541 VSS 7.34e-19
C7976 VDD.n1542 VSS 0.00101f
C7977 VDD.n1543 VSS 0.00207f
C7978 VDD.t234 VSS 5.71e-19
C7979 VDD.t340 VSS -1.82e-19
C7980 VDD.n1544 VSS 0.00268f
C7981 VDD.n1545 VSS 0.00243f
C7982 VDD.n1546 VSS 0.00134f
C7983 VDD.n1547 VSS 7.44e-19
C7984 VDD.n1548 VSS 0.00621f
C7985 VDD.n1549 VSS 7.34e-19
C7986 VDD.n1550 VSS 0.0012f
C7987 VDD.n1551 VSS 0.00207f
C7988 VDD.t442 VSS 6.16e-19
C7989 VDD.t232 VSS -3.41e-19
C7990 VDD.n1552 VSS 0.00241f
C7991 VDD.n1553 VSS 0.00164f
C7992 VDD.n1554 VSS 7.34e-19
C7993 VDD.t203 VSS 0.00389f
C7994 VDD.n1555 VSS 7.34e-19
C7995 VDD.t204 VSS 0.00176f
C7996 VDD.n1556 VSS 0.00177f
C7997 VDD.n1557 VSS 0.00281f
C7998 VDD.n1558 VSS 0.00207f
C7999 VDD.n1559 VSS 0.00137f
C8000 VDD.n1560 VSS 7.44e-19
C8001 VDD.n1561 VSS 0.00422f
C8002 VDD.n1562 VSS 7.34e-19
C8003 VDD.n1563 VSS 0.00125f
C8004 VDD.n1564 VSS 0.00207f
C8005 VDD.n1565 VSS 0.00125f
C8006 VDD.n1566 VSS 7.34e-19
C8007 VDD.n1567 VSS 0.0041f
C8008 VDD.n1568 VSS 7.34e-19
C8009 VDD.t202 VSS 6.5e-19
C8010 VDD.t94 VSS 0.00146f
C8011 VDD.n1569 VSS 0.00234f
C8012 VDD.n1570 VSS 0.00307f
C8013 VDD.n1571 VSS 0.00207f
C8014 VDD.n1572 VSS 7.89e-19
C8015 VDD.n1573 VSS 7.34e-19
C8016 VDD.t95 VSS 0.00389f
C8017 VDD.n1574 VSS 7.34e-19
C8018 VDD.n1575 VSS 0.0012f
C8019 VDD.n1576 VSS 0.00207f
C8020 VDD.n1577 VSS 0.00101f
C8021 VDD.n1578 VSS 7.34e-19
C8022 VDD.n1579 VSS 0.00608f
C8023 VDD.n1580 VSS 7.34e-19
C8024 VDD.n1581 VSS 8.03e-19
C8025 VDD.t403 VSS 4.05e-19
C8026 VDD.t324 VSS 4.05e-19
C8027 VDD.n1582 VSS 8.77e-19
C8028 VDD.n1583 VSS 0.00101f
C8029 VDD.n1584 VSS 7.34e-19
C8030 VDD.t221 VSS 0.00389f
C8031 VDD.n1585 VSS 7.44e-19
C8032 VDD.n1586 VSS 0.00134f
C8033 VDD.n1587 VSS 0.00207f
C8034 VDD.n1588 VSS 0.0012f
C8035 VDD.n1589 VSS 7.34e-19
C8036 VDD.t51 VSS 0.00389f
C8037 VDD.n1590 VSS 7.34e-19
C8038 VDD.t52 VSS 6.16e-19
C8039 VDD.t728 VSS -3.41e-19
C8040 VDD.n1591 VSS 0.00241f
C8041 VDD.n1592 VSS 0.00164f
C8042 VDD.n1593 VSS 0.00207f
C8043 VDD.t557 VSS 0.00176f
C8044 VDD.n1594 VSS 0.00177f
C8045 VDD.n1595 VSS 7.34e-19
C8046 VDD.t615 VSS 0.00389f
C8047 VDD.n1596 VSS 7.44e-19
C8048 VDD.n1597 VSS 0.00137f
C8049 VDD.n1598 VSS 0.00105f
C8050 VDD.n1599 VSS 0.00207f
C8051 VDD.n1600 VSS 0.00125f
C8052 VDD.n1601 VSS 7.34e-19
C8053 VDD.n1602 VSS 0.00608f
C8054 VDD.n1603 VSS 7.34e-19
C8055 VDD.n1604 VSS 0.00125f
C8056 VDD.n1605 VSS 0.00207f
C8057 VDD.t559 VSS 6.5e-19
C8058 VDD.t27 VSS 0.00146f
C8059 VDD.n1606 VSS 0.00234f
C8060 VDD.n1607 VSS 0.00307f
C8061 VDD.n1608 VSS 7.34e-19
C8062 VDD.n1609 VSS 0.00443f
C8063 VDD.n1610 VSS 7.34e-19
C8064 VDD.n1611 VSS 7.89e-19
C8065 VDD.n1612 VSS 6.94e-19
C8066 VDD.n1613 VSS 0.00207f
C8067 VDD.t29 VSS 3.65e-19
C8068 VDD.t618 VSS 3.84e-19
C8069 VDD.n1614 VSS 8.01e-19
C8070 VDD.n1615 VSS 0.0012f
C8071 VDD.n1616 VSS 7.34e-19
C8072 VDD.t330 VSS 0.00389f
C8073 VDD.n1617 VSS 7.34e-19
C8074 VDD.n1618 VSS 0.00101f
C8075 VDD.n1619 VSS 0.00207f
C8076 VDD.t648 VSS 9.52e-19
C8077 VDD.n1620 VSS 8.03e-19
C8078 VDD.n1621 VSS 7.34e-19
C8079 VDD.t213 VSS 0.00313f
C8080 VDD.n1622 VSS 7.34e-19
C8081 VDD.n1623 VSS 0.00101f
C8082 VDD.n1624 VSS 0.00207f
C8083 VDD.t492 VSS 5.71e-19
C8084 VDD.t61 VSS -1.82e-19
C8085 VDD.n1625 VSS 0.00268f
C8086 VDD.n1626 VSS 0.00243f
C8087 VDD.n1627 VSS 0.00134f
C8088 VDD.n1628 VSS 7.44e-19
C8089 VDD.n1629 VSS 0.00621f
C8090 VDD.n1630 VSS 7.34e-19
C8091 VDD.n1631 VSS 0.0012f
C8092 VDD.n1632 VSS 0.00207f
C8093 VDD.t565 VSS 6.16e-19
C8094 VDD.t496 VSS -3.41e-19
C8095 VDD.n1633 VSS 0.00241f
C8096 VDD.n1634 VSS 0.00164f
C8097 VDD.n1635 VSS 7.34e-19
C8098 VDD.t205 VSS 0.00389f
C8099 VDD.n1636 VSS 7.34e-19
C8100 VDD.t206 VSS 0.00176f
C8101 VDD.n1637 VSS 0.00177f
C8102 VDD.n1638 VSS 0.00281f
C8103 VDD.n1639 VSS 0.00207f
C8104 VDD.n1640 VSS 0.00137f
C8105 VDD.n1641 VSS 7.44e-19
C8106 VDD.n1642 VSS 0.00422f
C8107 VDD.n1643 VSS 7.34e-19
C8108 VDD.n1644 VSS 0.00125f
C8109 VDD.n1645 VSS 0.00207f
C8110 VDD.n1646 VSS 0.00125f
C8111 VDD.n1647 VSS 7.34e-19
C8112 VDD.n1648 VSS 0.0041f
C8113 VDD.n1649 VSS 7.34e-19
C8114 VDD.t208 VSS 6.5e-19
C8115 VDD.t474 VSS 0.00146f
C8116 VDD.n1650 VSS 0.00234f
C8117 VDD.n1651 VSS 0.00307f
C8118 VDD.n1652 VSS 0.00207f
C8119 VDD.n1653 VSS 7.89e-19
C8120 VDD.n1654 VSS 7.34e-19
C8121 VDD.t475 VSS 0.00389f
C8122 VDD.n1655 VSS 7.34e-19
C8123 VDD.n1656 VSS 0.0012f
C8124 VDD.n1657 VSS 0.00207f
C8125 VDD.n1658 VSS 0.00101f
C8126 VDD.n1659 VSS 7.34e-19
C8127 VDD.n1660 VSS 0.00608f
C8128 VDD.n1661 VSS 7.34e-19
C8129 VDD.n1662 VSS 8.03e-19
C8130 VDD.t291 VSS 4.05e-19
C8131 VDD.t307 VSS 4.05e-19
C8132 VDD.n1663 VSS 8.77e-19
C8133 VDD.n1664 VSS 7.44e-19
C8134 VDD.t306 VSS 0.00389f
C8135 VDD.n1665 VSS 0.00355f
C8136 VDD.t290 VSS 0.00313f
C8137 VDD.n1666 VSS 0.00243f
C8138 VDD.n1667 VSS 0.00106f
C8139 VDD.n1668 VSS 0.00136f
C8140 VDD.n1669 VSS 0.00182f
C8141 VDD.n1670 VSS 0.00187f
C8142 VDD.n1671 VSS 0.00207f
C8143 VDD.n1672 VSS 0.00207f
C8144 VDD.t658 VSS 9.52e-19
C8145 VDD.n1673 VSS 0.00207f
C8146 VDD.n1674 VSS 0.00136f
C8147 VDD.n1675 VSS 7.44e-19
C8148 VDD.n1676 VSS 0.00574f
C8149 VDD.t657 VSS 0.00389f
C8150 VDD.n1677 VSS 0.00393f
C8151 VDD.t71 VSS 0.00389f
C8152 VDD.n1678 VSS 0.00507f
C8153 VDD.t305 VSS 0.00389f
C8154 VDD.n1679 VSS 0.00355f
C8155 VDD.n1680 VSS 7.34e-19
C8156 VDD.n1681 VSS 0.00125f
C8157 VDD.n1682 VSS 0.00207f
C8158 VDD.n1683 VSS 0.00207f
C8159 VDD.n1684 VSS 0.00207f
C8160 VDD.n1685 VSS 0.00207f
C8161 VDD.t476 VSS 3.65e-19
C8162 VDD.t732 VSS 3.84e-19
C8163 VDD.n1686 VSS 8.01e-19
C8164 VDD.n1687 VSS 0.00187f
C8165 VDD.n1688 VSS 0.00137f
C8166 VDD.n1689 VSS 7.44e-19
C8167 VDD.n1690 VSS 0.00448f
C8168 VDD.t731 VSS 0.00389f
C8169 VDD.n1691 VSS 0.00443f
C8170 VDD.t207 VSS 0.00376f
C8171 VDD.t190 VSS 0.00367f
C8172 VDD.n1692 VSS 0.00401f
C8173 VDD.n1693 VSS 7.34e-19
C8174 VDD.n1694 VSS 0.00125f
C8175 VDD.n1695 VSS 6.94e-19
C8176 VDD.n1696 VSS 0.00207f
C8177 VDD.n1697 VSS 0.00207f
C8178 VDD.n1698 VSS 7.35e-19
C8179 VDD.n1699 VSS 7.34e-19
C8180 VDD.n1700 VSS 0.00557f
C8181 VDD.t473 VSS 0.00389f
C8182 VDD.n1701 VSS 0.00608f
C8183 VDD.t72 VSS 0.00389f
C8184 VDD.t304 VSS 0.00743f
C8185 VDD.n1702 VSS 7.34e-19
C8186 VDD.n1703 VSS 0.00125f
C8187 VDD.n1704 VSS 0.00207f
C8188 VDD.n1705 VSS 0.00207f
C8189 VDD.t494 VSS 3.84e-19
C8190 VDD.t734 VSS 3.84e-19
C8191 VDD.n1706 VSS 8.11e-19
C8192 VDD.n1707 VSS 0.0017f
C8193 VDD.n1708 VSS 0.00207f
C8194 VDD.n1709 VSS 0.00207f
C8195 VDD.n1710 VSS 8.91e-19
C8196 VDD.n1711 VSS 7.34e-19
C8197 VDD.n1712 VSS 0.00465f
C8198 VDD.t493 VSS 0.00389f
C8199 VDD.n1713 VSS 0.00456f
C8200 VDD.t733 VSS 0.00389f
C8201 VDD.n1714 VSS 0.00304f
C8202 VDD.t483 VSS 0.00389f
C8203 VDD.n1715 VSS 0.00405f
C8204 VDD.n1716 VSS 7.34e-19
C8205 VDD.n1717 VSS 0.0011f
C8206 VDD.n1718 VSS 0.00105f
C8207 VDD.n1719 VSS 0.00207f
C8208 VDD.n1720 VSS 0.00207f
C8209 VDD.n1721 VSS 0.00195f
C8210 VDD.n1722 VSS 7.34e-19
C8211 VDD.n1723 VSS 0.00701f
C8212 VDD.n1724 VSS 0.00524f
C8213 VDD.t564 VSS 0.00389f
C8214 VDD.t495 VSS 0.00389f
C8215 VDD.n1725 VSS 0.0041f
C8216 VDD.n1726 VSS 7.34e-19
C8217 VDD.n1727 VSS 0.00125f
C8218 VDD.n1728 VSS 0.00207f
C8219 VDD.n1729 VSS 0.00207f
C8220 VDD.n1730 VSS 0.00207f
C8221 VDD.n1731 VSS 0.00109f
C8222 VDD.n1732 VSS 7.34e-19
C8223 VDD.n1733 VSS 0.00562f
C8224 VDD.t491 VSS 0.00389f
C8225 VDD.n1734 VSS 0.00401f
C8226 VDD.t60 VSS 0.00389f
C8227 VDD.n1735 VSS 0.00393f
C8228 VDD.n1736 VSS 0.00591f
C8229 VDD.n1737 VSS 7.34e-19
C8230 VDD.n1738 VSS 0.00101f
C8231 VDD.n1739 VSS 0.00155f
C8232 VDD.n1740 VSS 7.21e-19
C8233 VDD.n1741 VSS 0.00187f
C8234 VDD.t214 VSS 4.05e-19
C8235 VDD.t528 VSS 4.05e-19
C8236 VDD.n1742 VSS 8.77e-19
C8237 VDD.n1743 VSS 0.00182f
C8238 VDD.n1744 VSS 0.00136f
C8239 VDD.n1745 VSS 7.44e-19
C8240 VDD.n1746 VSS 0.00355f
C8241 VDD.t527 VSS 0.00389f
C8242 VDD.n1747 VSS 0.00608f
C8243 VDD.n1748 VSS 0.00393f
C8244 VDD.t647 VSS 0.00389f
C8245 VDD.n1749 VSS 0.00574f
C8246 VDD.n1750 VSS 7.44e-19
C8247 VDD.n1751 VSS 0.00136f
C8248 VDD.n1752 VSS 0.00207f
C8249 VDD.n1753 VSS 0.00207f
C8250 VDD.n1754 VSS 0.00207f
C8251 VDD.n1755 VSS 0.00207f
C8252 VDD.n1756 VSS 0.00125f
C8253 VDD.n1757 VSS 7.34e-19
C8254 VDD.n1758 VSS 0.00355f
C8255 VDD.t526 VSS 0.00389f
C8256 VDD.n1759 VSS 0.00507f
C8257 VDD.t28 VSS 0.00389f
C8258 VDD.t617 VSS 0.00389f
C8259 VDD.n1760 VSS 0.00448f
C8260 VDD.n1761 VSS 7.44e-19
C8261 VDD.n1762 VSS 0.00137f
C8262 VDD.n1763 VSS 0.00187f
C8263 VDD.n1764 VSS 0.00207f
C8264 VDD.n1765 VSS 0.00207f
C8265 VDD.n1766 VSS 0.00207f
C8266 VDD.n1767 VSS 0.00125f
C8267 VDD.n1768 VSS 7.34e-19
C8268 VDD.n1769 VSS 0.00401f
C8269 VDD.t739 VSS 0.00367f
C8270 VDD.t558 VSS 0.00376f
C8271 VDD.n1770 VSS 0.0041f
C8272 VDD.t26 VSS 0.00389f
C8273 VDD.n1771 VSS 0.00557f
C8274 VDD.n1772 VSS 7.34e-19
C8275 VDD.n1773 VSS 7.35e-19
C8276 VDD.n1774 VSS 0.00207f
C8277 VDD.n1775 VSS 0.00207f
C8278 VDD.n1776 VSS 0.00207f
C8279 VDD.n1777 VSS 0.00125f
C8280 VDD.n1778 VSS 7.34e-19
C8281 VDD.t525 VSS 0.00743f
C8282 VDD.t331 VSS 0.00389f
C8283 VDD.n1779 VSS 0.00422f
C8284 VDD.n1780 VSS 0.00456f
C8285 VDD.t725 VSS 0.00389f
C8286 VDD.n1781 VSS 0.00465f
C8287 VDD.n1782 VSS 7.34e-19
C8288 VDD.n1783 VSS 8.91e-19
C8289 VDD.n1784 VSS 0.00207f
C8290 VDD.t726 VSS 3.84e-19
C8291 VDD.t616 VSS 3.84e-19
C8292 VDD.n1785 VSS 8.11e-19
C8293 VDD.n1786 VSS 0.0017f
C8294 VDD.n1787 VSS 0.00207f
C8295 VDD.n1788 VSS 0.00207f
C8296 VDD.n1789 VSS 0.00207f
C8297 VDD.n1790 VSS 0.0011f
C8298 VDD.n1791 VSS 7.34e-19
C8299 VDD.n1792 VSS 0.00405f
C8300 VDD.t406 VSS 0.00389f
C8301 VDD.n1793 VSS 0.00304f
C8302 VDD.t556 VSS 0.00389f
C8303 VDD.n1794 VSS 0.00524f
C8304 VDD.n1795 VSS 0.00701f
C8305 VDD.n1796 VSS 7.34e-19
C8306 VDD.n1797 VSS 0.00195f
C8307 VDD.n1798 VSS 0.00281f
C8308 VDD.n1799 VSS 0.00207f
C8309 VDD.n1800 VSS 0.00207f
C8310 VDD.n1801 VSS 0.00125f
C8311 VDD.n1802 VSS 7.34e-19
C8312 VDD.n1803 VSS 0.0041f
C8313 VDD.t727 VSS 0.00389f
C8314 VDD.n1804 VSS 0.00621f
C8315 VDD.n1805 VSS 0.00401f
C8316 VDD.t729 VSS 0.00389f
C8317 VDD.n1806 VSS 0.00562f
C8318 VDD.n1807 VSS 7.34e-19
C8319 VDD.n1808 VSS 0.00109f
C8320 VDD.n1809 VSS 0.00207f
C8321 VDD.t730 VSS 5.71e-19
C8322 VDD.t222 VSS -1.82e-19
C8323 VDD.n1810 VSS 0.00268f
C8324 VDD.n1811 VSS 0.00243f
C8325 VDD.n1812 VSS 0.00207f
C8326 VDD.n1813 VSS 7.21e-19
C8327 VDD.n1814 VSS 0.00155f
C8328 VDD.n1815 VSS 0.00101f
C8329 VDD.n1816 VSS 7.34e-19
C8330 VDD.n1817 VSS 0.00591f
C8331 VDD.n1818 VSS 0.00393f
C8332 VDD.t402 VSS 0.00313f
C8333 VDD.t323 VSS 0.00389f
C8334 VDD.n1819 VSS 0.00355f
C8335 VDD.n1820 VSS 7.44e-19
C8336 VDD.n1821 VSS 0.00136f
C8337 VDD.n1822 VSS 0.00182f
C8338 VDD.n1823 VSS 0.00187f
C8339 VDD.n1824 VSS 0.00207f
C8340 VDD.n1825 VSS 0.00207f
C8341 VDD.t650 VSS 9.52e-19
C8342 VDD.n1826 VSS 0.00207f
C8343 VDD.n1827 VSS 0.00136f
C8344 VDD.n1828 VSS 7.44e-19
C8345 VDD.n1829 VSS 0.00574f
C8346 VDD.t649 VSS 0.00389f
C8347 VDD.n1830 VSS 0.00393f
C8348 VDD.t88 VSS 0.00389f
C8349 VDD.n1831 VSS 0.00507f
C8350 VDD.t325 VSS 0.00389f
C8351 VDD.n1832 VSS 0.00355f
C8352 VDD.n1833 VSS 7.34e-19
C8353 VDD.n1834 VSS 0.00125f
C8354 VDD.n1835 VSS 0.00207f
C8355 VDD.n1836 VSS 0.00207f
C8356 VDD.n1837 VSS 0.00207f
C8357 VDD.n1838 VSS 0.00207f
C8358 VDD.t96 VSS 3.65e-19
C8359 VDD.t630 VSS 3.84e-19
C8360 VDD.n1839 VSS 8.01e-19
C8361 VDD.n1840 VSS 0.00187f
C8362 VDD.n1841 VSS 0.00137f
C8363 VDD.n1842 VSS 7.44e-19
C8364 VDD.n1843 VSS 0.00448f
C8365 VDD.t629 VSS 0.00389f
C8366 VDD.n1844 VSS 0.00443f
C8367 VDD.t201 VSS 0.00376f
C8368 VDD.t314 VSS 0.00367f
C8369 VDD.n1845 VSS 0.00401f
C8370 VDD.n1846 VSS 7.34e-19
C8371 VDD.n1847 VSS 0.00125f
C8372 VDD.n1848 VSS 6.94e-19
C8373 VDD.n1849 VSS 0.00207f
C8374 VDD.n1850 VSS 0.00207f
C8375 VDD.n1851 VSS 7.35e-19
C8376 VDD.n1852 VSS 7.34e-19
C8377 VDD.n1853 VSS 0.00557f
C8378 VDD.t93 VSS 0.00389f
C8379 VDD.n1854 VSS 0.00608f
C8380 VDD.t87 VSS 0.00389f
C8381 VDD.t322 VSS 0.00743f
C8382 VDD.n1855 VSS 7.34e-19
C8383 VDD.n1856 VSS 0.00125f
C8384 VDD.n1857 VSS 0.00207f
C8385 VDD.n1858 VSS 0.00207f
C8386 VDD.t230 VSS 3.84e-19
C8387 VDD.t628 VSS 3.84e-19
C8388 VDD.n1859 VSS 8.11e-19
C8389 VDD.n1860 VSS 0.0017f
C8390 VDD.n1861 VSS 0.00207f
C8391 VDD.n1862 VSS 0.00207f
C8392 VDD.n1863 VSS 8.91e-19
C8393 VDD.n1864 VSS 7.34e-19
C8394 VDD.n1865 VSS 0.00465f
C8395 VDD.t229 VSS 0.00389f
C8396 VDD.n1866 VSS 0.00456f
C8397 VDD.t627 VSS 0.00389f
C8398 VDD.n1867 VSS 0.00304f
C8399 VDD.t397 VSS 0.00389f
C8400 VDD.n1868 VSS 0.00405f
C8401 VDD.n1869 VSS 7.34e-19
C8402 VDD.n1870 VSS 0.0011f
C8403 VDD.n1871 VSS 0.00105f
C8404 VDD.n1872 VSS 0.00207f
C8405 VDD.n1873 VSS 0.00207f
C8406 VDD.n1874 VSS 0.00195f
C8407 VDD.n1875 VSS 7.34e-19
C8408 VDD.n1876 VSS 0.00701f
C8409 VDD.n1877 VSS 0.00524f
C8410 VDD.t441 VSS 0.00389f
C8411 VDD.t231 VSS 0.00389f
C8412 VDD.n1878 VSS 0.0041f
C8413 VDD.n1879 VSS 7.34e-19
C8414 VDD.n1880 VSS 0.00125f
C8415 VDD.n1881 VSS 0.00207f
C8416 VDD.n1882 VSS 0.00207f
C8417 VDD.n1883 VSS 0.00207f
C8418 VDD.n1884 VSS 0.00109f
C8419 VDD.n1885 VSS 7.34e-19
C8420 VDD.n1886 VSS 0.00562f
C8421 VDD.t233 VSS 0.00389f
C8422 VDD.n1887 VSS 0.00401f
C8423 VDD.t339 VSS 0.00389f
C8424 VDD.n1888 VSS 0.00393f
C8425 VDD.n1889 VSS 0.00591f
C8426 VDD.n1890 VSS 7.34e-19
C8427 VDD.n1891 VSS 0.00101f
C8428 VDD.n1892 VSS 0.00155f
C8429 VDD.n1893 VSS 7.21e-19
C8430 VDD.n1894 VSS 0.00187f
C8431 VDD.t410 VSS 4.05e-19
C8432 VDD.t219 VSS 4.05e-19
C8433 VDD.n1895 VSS 8.77e-19
C8434 VDD.n1896 VSS 0.00182f
C8435 VDD.n1897 VSS 0.00136f
C8436 VDD.n1898 VSS 7.44e-19
C8437 VDD.n1899 VSS 0.00355f
C8438 VDD.t218 VSS 0.00389f
C8439 VDD.n1900 VSS 0.00608f
C8440 VDD.n1901 VSS 0.00393f
C8441 VDD.t643 VSS 0.00389f
C8442 VDD.n1902 VSS 0.00574f
C8443 VDD.n1903 VSS 7.44e-19
C8444 VDD.n1904 VSS 0.00136f
C8445 VDD.n1905 VSS 0.00207f
C8446 VDD.n1906 VSS 0.00207f
C8447 VDD.n1907 VSS 0.00207f
C8448 VDD.n1908 VSS 0.00207f
C8449 VDD.n1909 VSS 0.00125f
C8450 VDD.n1910 VSS 7.34e-19
C8451 VDD.n1911 VSS 0.00355f
C8452 VDD.t217 VSS 0.00389f
C8453 VDD.n1912 VSS 0.00507f
C8454 VDD.t119 VSS 0.00389f
C8455 VDD.t384 VSS 0.00389f
C8456 VDD.n1913 VSS 0.00448f
C8457 VDD.n1914 VSS 7.44e-19
C8458 VDD.n1915 VSS 0.00137f
C8459 VDD.n1916 VSS 0.00187f
C8460 VDD.n1917 VSS 0.00207f
C8461 VDD.n1918 VSS 0.00207f
C8462 VDD.n1919 VSS 0.00207f
C8463 VDD.n1920 VSS 0.00125f
C8464 VDD.n1921 VSS 7.34e-19
C8465 VDD.n1922 VSS 0.00401f
C8466 VDD.t484 VSS 0.00367f
C8467 VDD.t89 VSS 0.00376f
C8468 VDD.n1923 VSS 0.0041f
C8469 VDD.t121 VSS 0.00389f
C8470 VDD.n1924 VSS 0.00557f
C8471 VDD.n1925 VSS 7.34e-19
C8472 VDD.n1926 VSS 7.35e-19
C8473 VDD.n1927 VSS 0.00207f
C8474 VDD.n1928 VSS 0.00207f
C8475 VDD.n1929 VSS 0.00207f
C8476 VDD.n1930 VSS 0.00125f
C8477 VDD.n1931 VSS 7.34e-19
C8478 VDD.t220 VSS 0.00743f
C8479 VDD.t199 VSS 0.00389f
C8480 VDD.n1932 VSS 0.00422f
C8481 VDD.n1933 VSS 0.00456f
C8482 VDD.t35 VSS 0.00389f
C8483 VDD.n1934 VSS 0.00465f
C8484 VDD.n1935 VSS 7.34e-19
C8485 VDD.n1936 VSS 8.91e-19
C8486 VDD.n1937 VSS 0.00207f
C8487 VDD.t36 VSS 3.84e-19
C8488 VDD.t387 VSS 3.84e-19
C8489 VDD.n1938 VSS 8.11e-19
C8490 VDD.n1939 VSS 0.0017f
C8491 VDD.n1940 VSS 0.00207f
C8492 VDD.n1941 VSS 0.00207f
C8493 VDD.n1942 VSS 0.00207f
C8494 VDD.n1943 VSS 0.0011f
C8495 VDD.n1944 VSS 7.34e-19
C8496 VDD.n1945 VSS 0.00405f
C8497 VDD.t8 VSS 0.00389f
C8498 VDD.n1946 VSS 0.00304f
C8499 VDD.t91 VSS 0.00389f
C8500 VDD.n1947 VSS 0.00524f
C8501 VDD.n1948 VSS 0.00701f
C8502 VDD.n1949 VSS 7.34e-19
C8503 VDD.n1950 VSS 0.00195f
C8504 VDD.n1951 VSS 0.00281f
C8505 VDD.n1952 VSS 0.00207f
C8506 VDD.n1953 VSS 0.00207f
C8507 VDD.n1954 VSS 0.00125f
C8508 VDD.n1955 VSS 7.34e-19
C8509 VDD.n1956 VSS 0.0041f
C8510 VDD.t31 VSS 0.00389f
C8511 VDD.n1957 VSS 0.00621f
C8512 VDD.n1958 VSS 0.00401f
C8513 VDD.t33 VSS 0.00389f
C8514 VDD.n1959 VSS 0.00562f
C8515 VDD.n1960 VSS 7.34e-19
C8516 VDD.n1961 VSS 0.00109f
C8517 VDD.n1962 VSS 0.00207f
C8518 VDD.t34 VSS 5.71e-19
C8519 VDD.t742 VSS -1.82e-19
C8520 VDD.n1963 VSS 0.00268f
C8521 VDD.n1964 VSS 0.00243f
C8522 VDD.n1965 VSS 0.00207f
C8523 VDD.n1966 VSS 7.21e-19
C8524 VDD.n1967 VSS 0.00155f
C8525 VDD.n1968 VSS 0.00101f
C8526 VDD.n1969 VSS 7.34e-19
C8527 VDD.n1970 VSS 0.00591f
C8528 VDD.n1971 VSS 0.00393f
C8529 VDD.t631 VSS 0.00313f
C8530 VDD.t531 VSS 0.00389f
C8531 VDD.n1972 VSS 0.00355f
C8532 VDD.n1973 VSS 7.44e-19
C8533 VDD.n1974 VSS 0.00136f
C8534 VDD.n1975 VSS 0.00182f
C8535 VDD.n1976 VSS 0.00187f
C8536 VDD.n1977 VSS 0.00207f
C8537 VDD.n1978 VSS 0.00207f
C8538 VDD.t654 VSS 9.52e-19
C8539 VDD.n1979 VSS 0.00207f
C8540 VDD.n1980 VSS 0.00136f
C8541 VDD.n1981 VSS 7.44e-19
C8542 VDD.n1982 VSS 0.00574f
C8543 VDD.t653 VSS 0.00389f
C8544 VDD.n1983 VSS 0.00393f
C8545 VDD.t215 VSS 0.00389f
C8546 VDD.n1984 VSS 0.00507f
C8547 VDD.t529 VSS 0.00389f
C8548 VDD.n1985 VSS 0.00355f
C8549 VDD.n1986 VSS 7.34e-19
C8550 VDD.n1987 VSS 0.00125f
C8551 VDD.n1988 VSS 0.00207f
C8552 VDD.n1989 VSS 0.00207f
C8553 VDD.n1990 VSS 0.00207f
C8554 VDD.n1991 VSS 0.00207f
C8555 VDD.t246 VSS 3.65e-19
C8556 VDD.t106 VSS 3.84e-19
C8557 VDD.n1992 VSS 8.01e-19
C8558 VDD.n1993 VSS 0.00187f
C8559 VDD.n1994 VSS 0.00137f
C8560 VDD.n1995 VSS 7.44e-19
C8561 VDD.n1996 VSS 0.00448f
C8562 VDD.t105 VSS 0.00389f
C8563 VDD.n1997 VSS 0.00443f
C8564 VDD.t487 VSS 0.00376f
C8565 VDD.t332 VSS 0.00367f
C8566 VDD.n1998 VSS 0.00401f
C8567 VDD.n1999 VSS 7.34e-19
C8568 VDD.n2000 VSS 0.00125f
C8569 VDD.n2001 VSS 6.94e-19
C8570 VDD.n2002 VSS 0.00207f
C8571 VDD.n2003 VSS 0.00207f
C8572 VDD.n2004 VSS 7.35e-19
C8573 VDD.n2005 VSS 7.34e-19
C8574 VDD.n2006 VSS 0.00557f
C8575 VDD.t243 VSS 0.00389f
C8576 VDD.n2007 VSS 0.00608f
C8577 VDD.t216 VSS 0.00389f
C8578 VDD.t530 VSS 0.00743f
C8579 VDD.n2008 VSS 7.34e-19
C8580 VDD.n2009 VSS 0.00125f
C8581 VDD.n2010 VSS 0.00207f
C8582 VDD.n2011 VSS 0.00207f
C8583 VDD.t591 VSS 3.84e-19
C8584 VDD.t108 VSS 3.84e-19
C8585 VDD.n2012 VSS 8.11e-19
C8586 VDD.n2013 VSS 0.0017f
C8587 VDD.n2014 VSS 0.00207f
C8588 VDD.n2015 VSS 0.00207f
C8589 VDD.n2016 VSS 8.91e-19
C8590 VDD.n2017 VSS 7.34e-19
C8591 VDD.n2018 VSS 0.00465f
C8592 VDD.t590 VSS 0.00389f
C8593 VDD.n2019 VSS 0.00456f
C8594 VDD.t107 VSS 0.00389f
C8595 VDD.n2020 VSS 0.00304f
C8596 VDD.t612 VSS 0.00389f
C8597 VDD.n2021 VSS 0.00405f
C8598 VDD.n2022 VSS 7.34e-19
C8599 VDD.n2023 VSS 0.0011f
C8600 VDD.n2024 VSS 0.00105f
C8601 VDD.n2025 VSS 0.00207f
C8602 VDD.n2026 VSS 0.00207f
C8603 VDD.n2027 VSS 0.00195f
C8604 VDD.n2028 VSS 7.34e-19
C8605 VDD.n2029 VSS 0.00701f
C8606 VDD.n2030 VSS 0.00524f
C8607 VDD.t425 VSS 0.00389f
C8608 VDD.t588 VSS 0.00389f
C8609 VDD.n2031 VSS 0.0041f
C8610 VDD.n2032 VSS 7.34e-19
C8611 VDD.n2033 VSS 0.00125f
C8612 VDD.n2034 VSS 0.00207f
C8613 VDD.n2035 VSS 0.00207f
C8614 VDD.n2036 VSS 0.00207f
C8615 VDD.n2037 VSS 0.00109f
C8616 VDD.n2038 VSS 7.34e-19
C8617 VDD.n2039 VSS 0.00562f
C8618 VDD.t586 VSS 0.00389f
C8619 VDD.n2040 VSS 0.00401f
C8620 VDD.t677 VSS 0.00445f
C8621 VDD.n2041 VSS 0.00914f
C8622 VDD.n2042 VSS 0.00101f
C8623 VDD.n2043 VSS 0.00155f
C8624 VDD.n2044 VSS 1.19f
C8625 VDD.n2045 VSS 0.0312f
C8626 VDD.n2046 VSS 0.00786f
C8627 VDD.n2047 VSS 0.365f
C8628 VDD.n2048 VSS 0.67f
C8629 VDD.n2049 VSS 0.00207f
C8630 VDD.t563 VSS 5.37e-19
C8631 VDD.t282 VSS 5.37e-19
C8632 VDD.n2050 VSS 0.0013f
C8633 VDD.n2051 VSS 0.00246f
C8634 VDD.n2052 VSS 0.00136f
C8635 VDD.n2053 VSS 7.44e-19
C8636 VDD.n2054 VSS 7.34e-19
C8637 VDD.n2055 VSS 0.00207f
C8638 VDD.t192 VSS 6.33e-19
C8639 VDD.t561 VSS 6.33e-19
C8640 VDD.n2056 VSS 0.00145f
C8641 VDD.n2057 VSS 0.00225f
C8642 VDD.n2058 VSS 7.34e-19
C8643 VDD.t193 VSS 0.00459f
C8644 VDD.n2059 VSS 3.95e-19
C8645 VDD.t194 VSS 6.33e-19
C8646 VDD.t196 VSS 6.33e-19
C8647 VDD.n2060 VSS 0.0015f
C8648 VDD.n2061 VSS 0.00257f
C8649 VDD.n2062 VSS 0.00207f
C8650 VDD.n2063 VSS 0.00123f
C8651 VDD.t416 VSS 0.00295f
C8652 VDD.n2064 VSS 7.34e-19
C8653 VDD.t413 VSS 0.00391f
C8654 VDD.n2065 VSS 7.34e-19
C8655 VDD.n2066 VSS 0.00125f
C8656 VDD.t414 VSS 0.00101f
C8657 VDD.t412 VSS 6.33e-19
C8658 VDD.n2067 VSS 0.00211f
C8659 VDD.n2068 VSS 0.00283f
C8660 VDD.n2069 VSS 0.00207f
C8661 VDD.t80 VSS 6.01e-19
C8662 VDD.t418 VSS 2.93e-19
C8663 VDD.n2070 VSS 0.00217f
C8664 VDD.n2071 VSS 0.00173f
C8665 VDD.n2072 VSS 7.34e-19
C8666 VDD.t698 VSS 0.00391f
C8667 VDD.n2073 VSS 7.34e-19
C8668 VDD.n2074 VSS 0.00125f
C8669 VDD.n2075 VSS 0.00122f
C8670 VDD.n2076 VSS 0.00207f
C8671 VDD.t539 VSS 0.00151f
C8672 VDD.n2077 VSS 0.00244f
C8673 VDD.n2078 VSS 0.00136f
C8674 VDD.n2079 VSS 7.44e-19
C8675 VDD.t501 VSS 0.00391f
C8676 VDD.n2080 VSS 7.34e-19
C8677 VDD.n2081 VSS 0.00125f
C8678 VDD.n2082 VSS 0.00207f
C8679 VDD.n2083 VSS 0.001f
C8680 VDD.n2084 VSS 7.34e-19
C8681 VDD.t308 VSS 0.00391f
C8682 VDD.n2085 VSS 7.34e-19
C8683 VDD.n2086 VSS 0.00125f
C8684 VDD.t309 VSS 4.05e-19
C8685 VDD.t5 VSS 4.05e-19
C8686 VDD.n2087 VSS 8.7e-19
C8687 VDD.n2088 VSS 0.00182f
C8688 VDD.n2089 VSS 0.00207f
C8689 VDD.n2090 VSS 0.00104f
C8690 VDD.n2091 VSS 7.34e-19
C8691 VDD.t404 VSS 0.00314f
C8692 VDD.n2092 VSS 0.00708f
C8693 VDD.n2093 VSS 0.00105f
C8694 VDD.n2094 VSS 0.00187f
C8695 VDD.t405 VSS 4.05e-19
C8696 VDD.t519 VSS 4.05e-19
C8697 VDD.n2095 VSS 8.53e-19
C8698 VDD.n2096 VSS 0.00147f
C8699 VDD.n2097 VSS 0.00136f
C8700 VDD.n2098 VSS 7.44e-19
C8701 VDD.n2099 VSS 0.00357f
C8702 VDD.t518 VSS 0.00391f
C8703 VDD.n2100 VSS 0.00408f
C8704 VDD.t623 VSS 0.00391f
C8705 VDD.n2101 VSS 0.00611f
C8706 VDD.t697 VSS 0.00391f
C8707 VDD.n2102 VSS 0.00357f
C8708 VDD.n2103 VSS 7.34e-19
C8709 VDD.n2104 VSS 0.00125f
C8710 VDD.n2105 VSS 0.00207f
C8711 VDD.n2106 VSS 0.00207f
C8712 VDD.n2107 VSS 0.00207f
C8713 VDD.n2108 VSS 8.78e-19
C8714 VDD.n2109 VSS 7.34e-19
C8715 VDD.n2110 VSS 0.00357f
C8716 VDD.t4 VSS 0.00391f
C8717 VDD.n2111 VSS 0.00442f
C8718 VDD.n2112 VSS 0.00357f
C8719 VDD.t247 VSS 0.00391f
C8720 VDD.n2113 VSS 0.00747f
C8721 VDD.n2114 VSS 7.34e-19
C8722 VDD.n2115 VSS 0.00125f
C8723 VDD.n2116 VSS 0.00207f
C8724 VDD.n2117 VSS 0.00207f
C8725 VDD.n2118 VSS 0.00207f
C8726 VDD.n2119 VSS 0.00116f
C8727 VDD.n2120 VSS 7.34e-19
C8728 VDD.n2121 VSS 0.00459f
C8729 VDD.n2122 VSS 0.0073f
C8730 VDD.t538 VSS 0.00391f
C8731 VDD.n2123 VSS 0.00522f
C8732 VDD.n2124 VSS 0.00442f
C8733 VDD.n2125 VSS 7.34e-19
C8734 VDD.n2126 VSS 8.78e-19
C8735 VDD.n2127 VSS 0.00207f
C8736 VDD.n2128 VSS 0.00207f
C8737 VDD.n2129 VSS 0.00207f
C8738 VDD.n2130 VSS 0.00125f
C8739 VDD.n2131 VSS 7.34e-19
C8740 VDD.n2132 VSS 0.00357f
C8741 VDD.t537 VSS 0.00391f
C8742 VDD.n2133 VSS 0.00429f
C8743 VDD.t79 VSS 0.00391f
C8744 VDD.n2134 VSS 0.00357f
C8745 VDD.t417 VSS 0.00391f
C8746 VDD.n2135 VSS 0.00412f
C8747 VDD.n2136 VSS 7.34e-19
C8748 VDD.n2137 VSS 6.6e-19
C8749 VDD.n2138 VSS 0.00207f
C8750 VDD.n2139 VSS 0.00207f
C8751 VDD.n2140 VSS 0.00207f
C8752 VDD.n2141 VSS 6.46e-19
C8753 VDD.n2142 VSS 7.34e-19
C8754 VDD.n2143 VSS 0.00425f
C8755 VDD.t411 VSS 0.00391f
C8756 VDD.n2144 VSS 0.00357f
C8757 VDD.t415 VSS 0.00391f
C8758 VDD.t197 VSS 0.029f
C8759 VDD.n2145 VSS 0.0282f
C8760 VDD.n2146 VSS 7.34e-19
C8761 VDD.n2147 VSS 0.00412f
C8762 VDD.n2148 VSS 0.00155f
C8763 VDD.t198 VSS 0.00259f
C8764 VDD.n2149 VSS 0.00438f
C8765 VDD.n2150 VSS 0.00645f
C8766 VDD.n2151 VSS 0.00207f
C8767 VDD.n2152 VSS 0.00207f
C8768 VDD.n2153 VSS 0.00207f
C8769 VDD.n2154 VSS 8.71e-19
C8770 VDD.n2155 VSS 0.00133f
C8771 VDD.n2156 VSS 7.44e-19
C8772 VDD.n2157 VSS 0.00357f
C8773 VDD.t195 VSS 0.00391f
C8774 VDD.n2158 VSS 0.00357f
C8775 VDD.t191 VSS 0.00391f
C8776 VDD.n2159 VSS 0.00272f
C8777 VDD.t560 VSS 0.00391f
C8778 VDD.n2160 VSS 0.00357f
C8779 VDD.n2161 VSS 7.34e-19
C8780 VDD.n2162 VSS 6.6e-19
C8781 VDD.n2163 VSS 7.35e-19
C8782 VDD.n2164 VSS 0.00155f
C8783 VDD.n2165 VSS 0.00155f
C8784 VDD.n2166 VSS 9.19e-19
C8785 VDD.n2167 VSS 7.34e-19
C8786 VDD.n2168 VSS 0.00527f
C8787 VDD.t562 VSS 0.00391f
C8788 VDD.n2169 VSS 0.00374f
C8789 VDD.t281 VSS 0.00391f
C8790 VDD.n2170 VSS 0.00276f
C8791 VDD.n2171 VSS 7.34e-19
C8792 VDD.n2172 VSS 0.00103f
C8793 VDD.n2173 VSS 0.00123f
C8794 VDD.n2174 VSS 0.336f
C8795 VDD.n2175 VSS 0.00122f
C8796 VDD.t507 VSS 4.05e-19
C8797 VDD.t694 VSS 4.05e-19
C8798 VDD.n2176 VSS 8.77e-19
C8799 VDD.t506 VSS 0.0039f
C8800 VDD.n2177 VSS 0.00101f
C8801 VDD.n2178 VSS 7.34e-19
C8802 VDD.n2179 VSS 7.2e-19
C8803 VDD.t693 VSS 0.00385f
C8804 VDD.n2180 VSS 0.00356f
C8805 VDD.n2181 VSS 7.44e-19
C8806 VDD.n2182 VSS 0.00136f
C8807 VDD.n2183 VSS 0.00182f
C8808 VDD.n2184 VSS 0.00207f
C8809 VDD.n2185 VSS 0.0061f
C8810 VDD.n2186 VSS 7.34e-19
C8811 VDD.n2187 VSS 8.03e-19
C8812 VDD.n2188 VSS 0.00207f
C8813 VDD.t138 VSS 9.52e-19
C8814 VDD.t137 VSS 0.0039f
C8815 VDD.n2189 VSS 0.00576f
C8816 VDD.n2190 VSS 7.44e-19
C8817 VDD.n2191 VSS 0.00136f
C8818 VDD.n2192 VSS 0.00207f
C8819 VDD.n2193 VSS 0.00207f
C8820 VDD.t723 VSS 0.0039f
C8821 VDD.n2194 VSS 0.00394f
C8822 VDD.n2195 VSS 7.34e-19
C8823 VDD.n2196 VSS 0.00101f
C8824 VDD.n2197 VSS 0.00207f
C8825 VDD.t508 VSS 0.0039f
C8826 VDD.n2198 VSS 0.00356f
C8827 VDD.n2199 VSS 7.34e-19
C8828 VDD.n2200 VSS 0.00125f
C8829 VDD.n2201 VSS 0.00207f
C8830 VDD.n2202 VSS 0.00508f
C8831 VDD.n2203 VSS 7.34e-19
C8832 VDD.n2204 VSS 0.0012f
C8833 VDD.n2205 VSS 0.00207f
C8834 VDD.t444 VSS 3.84e-19
C8835 VDD.t393 VSS 3.65e-19
C8836 VDD.n2206 VSS 8.01e-19
C8837 VDD.t392 VSS 0.0039f
C8838 VDD.n2207 VSS 0.00449f
C8839 VDD.n2208 VSS 7.44e-19
C8840 VDD.n2209 VSS 0.00137f
C8841 VDD.n2210 VSS 0.00187f
C8842 VDD.n2211 VSS 0.00207f
C8843 VDD.t443 VSS 0.0039f
C8844 VDD.n2212 VSS 0.00445f
C8845 VDD.n2213 VSS 7.34e-19
C8846 VDD.n2214 VSS 7.89e-19
C8847 VDD.n2215 VSS 0.00207f
C8848 VDD.t98 VSS 0.00368f
C8849 VDD.n2216 VSS 0.00402f
C8850 VDD.n2217 VSS 7.34e-19
C8851 VDD.n2218 VSS 0.00125f
C8852 VDD.n2219 VSS 0.00207f
C8853 VDD.t395 VSS 0.00146f
C8854 VDD.t534 VSS 6.5e-19
C8855 VDD.n2220 VSS 0.00234f
C8856 VDD.n2221 VSS 0.00307f
C8857 VDD.t533 VSS 0.00377f
C8858 VDD.n2222 VSS 0.00411f
C8859 VDD.n2223 VSS 7.34e-19
C8860 VDD.n2224 VSS 6.94e-19
C8861 VDD.n2225 VSS 0.00207f
C8862 VDD.t394 VSS 0.0039f
C8863 VDD.n2226 VSS 0.00559f
C8864 VDD.n2227 VSS 7.34e-19
C8865 VDD.n2228 VSS 7.35e-19
C8866 VDD.n2229 VSS 0.00207f
C8867 VDD.n2230 VSS 0.0061f
C8868 VDD.n2231 VSS 7.34e-19
C8869 VDD.n2232 VSS 0.00125f
C8870 VDD.n2233 VSS 0.00207f
C8871 VDD.t509 VSS 0.00745f
C8872 VDD.n2234 VSS 7.34e-19
C8873 VDD.n2235 VSS 0.00125f
C8874 VDD.n2236 VSS 0.00207f
C8875 VDD.t724 VSS 0.0039f
C8876 VDD.n2237 VSS 0.00423f
C8877 VDD.n2238 VSS 7.34e-19
C8878 VDD.n2239 VSS 0.00125f
C8879 VDD.n2240 VSS 0.00207f
C8880 VDD.t225 VSS 0.0039f
C8881 VDD.n2241 VSS 0.00466f
C8882 VDD.n2242 VSS 7.34e-19
C8883 VDD.n2243 VSS 8.91e-19
C8884 VDD.n2244 VSS 0.00207f
C8885 VDD.t672 VSS 3.84e-19
C8886 VDD.t226 VSS 3.84e-19
C8887 VDD.n2245 VSS 8.11e-19
C8888 VDD.t671 VSS 0.0039f
C8889 VDD.n2246 VSS 0.00457f
C8890 VDD.n2247 VSS 7.44e-19
C8891 VDD.n2248 VSS 0.00137f
C8892 VDD.n2249 VSS 0.0017f
C8893 VDD.n2250 VSS 0.00207f
C8894 VDD.t663 VSS 0.0039f
C8895 VDD.n2251 VSS 0.00407f
C8896 VDD.n2252 VSS 7.34e-19
C8897 VDD.n2253 VSS 0.0011f
C8898 VDD.n2254 VSS 0.00207f
C8899 VDD.t535 VSS 0.0039f
C8900 VDD.n2255 VSS 0.00305f
C8901 VDD.n2256 VSS 7.34e-19
C8902 VDD.n2257 VSS 0.00105f
C8903 VDD.n2258 VSS 0.00207f
C8904 VDD.t185 VSS 0.00936f
C8905 VDD.n2259 VSS 0.00838f
C8906 VDD.n2260 VSS 9.01e-19
C8907 VDD.t536 VSS 0.00176f
C8908 VDD.n2261 VSS 0.00177f
C8909 VDD.n2262 VSS 0.00192f
C8910 VDD.n2263 VSS 0.00205f
C8911 VDD.n2264 VSS 0.00104f
C8912 VDD.t750 VSS 5.91e-19
C8913 VDD.n2265 VSS 0.00165f
C8914 VDD.t184 VSS 0.00108f
C8915 VDD.n2266 VSS 0.00225f
C8916 VDD.n2267 VSS 4.94e-19
C8917 VDD.n2268 VSS 0.00145f
C8918 VDD.n2269 VSS 2.67e-19
C8919 VDD.n2270 VSS 1.91e-19
C8920 VDD.n2271 VSS 0.00104f
C8921 VDD.t224 VSS -3.41e-19
C8922 VDD.t186 VSS 6.16e-19
C8923 VDD.n2272 VSS 0.00241f
C8924 VDD.n2273 VSS 0.00138f
C8925 VDD.n2274 VSS 0.00125f
C8926 VDD.n2275 VSS 0.0019f
C8927 VDD.t223 VSS 0.00644f
C8928 VDD.n2276 VSS 0.00622f
C8929 VDD.n2277 VSS 0.00114f
C8930 VDD.n2278 VSS 0.0012f
C8931 VDD.n2279 VSS 0.00207f
C8932 VDD.t227 VSS 0.0039f
C8933 VDD.n2280 VSS 0.00563f
C8934 VDD.n2281 VSS 7.34e-19
C8935 VDD.n2282 VSS 0.00109f
C8936 VDD.n2283 VSS 0.00207f
C8937 VDD.t718 VSS -1.82e-19
C8938 VDD.t228 VSS 5.71e-19
C8939 VDD.n2284 VSS 0.00268f
C8940 VDD.t717 VSS 0.0039f
C8941 VDD.n2285 VSS 0.00402f
C8942 VDD.n2286 VSS 7.44e-19
C8943 VDD.n2287 VSS 0.00134f
C8944 VDD.n2288 VSS 0.00243f
C8945 VDD.n2289 VSS 0.00207f
C8946 VDD.n2290 VSS 0.00155f
C8947 VDD.n2291 VSS 0.00101f
C8948 VDD.n2292 VSS 0.00101f
C8949 VDD.n2293 VSS 7.34e-19
C8950 VDD.n2294 VSS 7.2e-19
C8951 VDD.t685 VSS 0.00385f
C8952 VDD.n2295 VSS 0.00356f
C8953 VDD.n2296 VSS 7.44e-19
C8954 VDD.n2297 VSS 0.00124f
C8955 VDD.n2298 VSS 0.00182f
C8956 VDD.n2299 VSS 0.00188f
C8957 VDD.n2300 VSS 0.00104f
C8958 VDD.n2301 VSS 3.81e-19
C8959 VDD.n2302 VSS 1.16e-19
C8960 VDD.n2303 VSS 3.63e-19
C8961 VDD.n2304 VSS 6.78e-20
C8962 VDD.n2305 VSS 0.00385f
C8963 VDD.n2306 VSS 7.2e-19
C8964 VDD.n2307 VSS 0.00224f
C8965 VDD.n2308 VSS 3.71e-19
C8966 VDD.n2309 VSS 4.15e-19
C8967 VDD.n2310 VSS 1.22e-19
C8968 VDD.n2311 VSS 0.00123f
C8969 VDD.t614 VSS 9.52e-19
C8970 VDD.t613 VSS 0.0039f
C8971 VDD.n2312 VSS 0.00504f
C8972 VDD.n2313 VSS 6.76e-19
C8973 VDD.n2314 VSS 0.00125f
C8974 VDD.n2315 VSS 0.00207f
C8975 VDD.n2316 VSS 0.00207f
C8976 VDD.t504 VSS 0.0039f
C8977 VDD.n2317 VSS 0.00394f
C8978 VDD.n2318 VSS 7.34e-19
C8979 VDD.n2319 VSS 0.00101f
C8980 VDD.n2320 VSS 0.00207f
C8981 VDD.t302 VSS 0.0039f
C8982 VDD.n2321 VSS 0.00356f
C8983 VDD.n2322 VSS 7.34e-19
C8984 VDD.n2323 VSS 0.00125f
C8985 VDD.n2324 VSS 0.00207f
C8986 VDD.t582 VSS 0.00724f
C8987 VDD.n2325 VSS 0.00508f
C8988 VDD.n2326 VSS 0.00128f
C8989 VDD.n2327 VSS 0.0012f
C8990 VDD.n2328 VSS 0.00207f
C8991 VDD.n2329 VSS 0.00133f
C8992 VDD.t180 VSS 3.84e-19
C8993 VDD.t583 VSS 3.65e-19
C8994 VDD.n2330 VSS 7.99e-19
C8995 VDD.n2331 VSS 0.00189f
C8996 VDD.n2332 VSS 0.00199f
C8997 VDD.n2333 VSS 0.00104f
C8998 VDD.n2334 VSS 6.26e-19
C8999 VDD.t181 VSS 9.98e-19
C9000 VDD.t743 VSS 4.23e-19
C9001 VDD.n2335 VSS 0.00203f
C9002 VDD.n2336 VSS 8.3e-19
C9003 VDD.n2337 VSS 0.00257f
C9004 VDD.n2338 VSS 1.89e-19
C9005 VDD.n2339 VSS 1.56e-19
C9006 VDD.n2340 VSS 9.17e-20
C9007 VDD.n2341 VSS 1.15e-19
C9008 VDD.n2342 VSS 2.17e-19
C9009 VDD.n2343 VSS 5.52e-19
C9010 VDD.t759 VSS 4.24e-19
C9011 VDD.n2344 VSS 0.00188f
C9012 VDD.t178 VSS 0.00126f
C9013 VDD.n2345 VSS 0.00102f
C9014 VDD.n2346 VSS 1.51e-19
C9015 VDD.n2347 VSS 1.16e-19
C9016 VDD.n2348 VSS 1.91e-19
C9017 VDD.n2349 VSS 0.00104f
C9018 VDD.t37 VSS 0.00368f
C9019 VDD.t179 VSS 0.00894f
C9020 VDD.n2350 VSS 0.00457f
C9021 VDD.n2351 VSS 7.74e-19
C9022 VDD.n2352 VSS 0.00118f
C9023 VDD.n2353 VSS 0.00196f
C9024 VDD.t585 VSS 0.00146f
C9025 VDD.t420 VSS 6.5e-19
C9026 VDD.n2354 VSS 0.00234f
C9027 VDD.n2355 VSS 0.00307f
C9028 VDD.t419 VSS 0.00377f
C9029 VDD.n2356 VSS 0.00411f
C9030 VDD.n2357 VSS 7.34e-19
C9031 VDD.n2358 VSS 6.94e-19
C9032 VDD.n2359 VSS 0.00207f
C9033 VDD.t584 VSS 0.0039f
C9034 VDD.n2360 VSS 0.00559f
C9035 VDD.n2361 VSS 7.34e-19
C9036 VDD.n2362 VSS 7.35e-19
C9037 VDD.n2363 VSS 0.00207f
C9038 VDD.n2364 VSS 0.0061f
C9039 VDD.n2365 VSS 7.34e-19
C9040 VDD.n2366 VSS 0.00125f
C9041 VDD.n2367 VSS 0.00207f
C9042 VDD.t303 VSS 0.00745f
C9043 VDD.n2368 VSS 7.34e-19
C9044 VDD.n2369 VSS 0.00125f
C9045 VDD.n2370 VSS 0.00207f
C9046 VDD.t505 VSS 0.0039f
C9047 VDD.n2371 VSS 0.00423f
C9048 VDD.n2372 VSS 7.34e-19
C9049 VDD.n2373 VSS 0.00125f
C9050 VDD.n2374 VSS 0.00207f
C9051 VDD.t103 VSS 0.0039f
C9052 VDD.n2375 VSS 0.00466f
C9053 VDD.n2376 VSS 7.34e-19
C9054 VDD.n2377 VSS 8.91e-19
C9055 VDD.n2378 VSS 0.00207f
C9056 VDD.t183 VSS 3.84e-19
C9057 VDD.t104 VSS 3.84e-19
C9058 VDD.n2379 VSS 8.11e-19
C9059 VDD.t182 VSS 0.0039f
C9060 VDD.n2380 VSS 0.00457f
C9061 VDD.n2381 VSS 7.44e-19
C9062 VDD.n2382 VSS 0.00137f
C9063 VDD.n2383 VSS 0.0017f
C9064 VDD.n2384 VSS 0.00207f
C9065 VDD.t256 VSS 0.0039f
C9066 VDD.n2385 VSS 0.00407f
C9067 VDD.n2386 VSS 7.34e-19
C9068 VDD.n2387 VSS 0.0011f
C9069 VDD.n2388 VSS 0.00207f
C9070 VDD.t421 VSS 0.0039f
C9071 VDD.n2389 VSS 0.00305f
C9072 VDD.n2390 VSS 7.34e-19
C9073 VDD.n2391 VSS 0.00105f
C9074 VDD.n2392 VSS 0.00207f
C9075 VDD.n2393 VSS 0.00703f
C9076 VDD.n2394 VSS 7.34e-19
C9077 VDD.t422 VSS 0.00176f
C9078 VDD.n2395 VSS 0.00177f
C9079 VDD.n2396 VSS 0.00195f
C9080 VDD.n2397 VSS 0.00207f
C9081 VDD.t111 VSS 0.0039f
C9082 VDD.n2398 VSS 0.00525f
C9083 VDD.n2399 VSS 7.34e-19
C9084 VDD.n2400 VSS 0.00281f
C9085 VDD.n2401 VSS 0.00207f
C9086 VDD.t101 VSS 0.0039f
C9087 VDD.n2402 VSS 0.00411f
C9088 VDD.n2403 VSS 7.34e-19
C9089 VDD.t102 VSS -3.41e-19
C9090 VDD.t112 VSS 6.16e-19
C9091 VDD.n2404 VSS 0.00241f
C9092 VDD.n2405 VSS 0.00164f
C9093 VDD.n2406 VSS 0.00125f
C9094 VDD.n2407 VSS 0.00207f
C9095 VDD.n2408 VSS 0.00622f
C9096 VDD.n2409 VSS 7.34e-19
C9097 VDD.n2410 VSS 0.0012f
C9098 VDD.n2411 VSS 0.00207f
C9099 VDD.t99 VSS 0.0039f
C9100 VDD.n2412 VSS 0.00563f
C9101 VDD.n2413 VSS 7.34e-19
C9102 VDD.n2414 VSS 0.00109f
C9103 VDD.n2415 VSS 0.00207f
C9104 VDD.t720 VSS -1.82e-19
C9105 VDD.t100 VSS 5.71e-19
C9106 VDD.n2416 VSS 0.00268f
C9107 VDD.t719 VSS 0.0039f
C9108 VDD.n2417 VSS 0.00402f
C9109 VDD.n2418 VSS 7.44e-19
C9110 VDD.n2419 VSS 0.00134f
C9111 VDD.n2420 VSS 0.00243f
C9112 VDD.n2421 VSS 0.00207f
C9113 VDD.n2422 VSS 0.00155f
C9114 VDD.n2423 VSS 0.00101f
C9115 VDD.n2424 VSS 0.00101f
C9116 VDD.n2425 VSS 7.34e-19
C9117 VDD.n2426 VSS 7.2e-19
C9118 VDD.t683 VSS 0.00385f
C9119 VDD.n2427 VSS 0.00356f
C9120 VDD.n2428 VSS 7.44e-19
C9121 VDD.n2429 VSS 0.00136f
C9122 VDD.n2430 VSS 0.00182f
C9123 VDD.n2431 VSS 0.00207f
C9124 VDD.n2432 VSS 0.0061f
C9125 VDD.n2433 VSS 7.34e-19
C9126 VDD.n2434 VSS 8.03e-19
C9127 VDD.n2435 VSS 0.00207f
C9128 VDD.t70 VSS 9.52e-19
C9129 VDD.t69 VSS 0.0039f
C9130 VDD.n2436 VSS 0.00576f
C9131 VDD.n2437 VSS 7.44e-19
C9132 VDD.n2438 VSS 0.00136f
C9133 VDD.n2439 VSS 0.00207f
C9134 VDD.n2440 VSS 0.00207f
C9135 VDD.t407 VSS 0.0039f
C9136 VDD.n2441 VSS 0.00394f
C9137 VDD.n2442 VSS 7.34e-19
C9138 VDD.n2443 VSS 0.00101f
C9139 VDD.n2444 VSS 0.00207f
C9140 VDD.t737 VSS 0.0039f
C9141 VDD.n2445 VSS 0.00356f
C9142 VDD.n2446 VSS 7.34e-19
C9143 VDD.n2447 VSS 0.00125f
C9144 VDD.n2448 VSS 0.00207f
C9145 VDD.t328 VSS 0.00724f
C9146 VDD.n2449 VSS 0.00508f
C9147 VDD.n2450 VSS 0.00128f
C9148 VDD.n2451 VSS 0.0012f
C9149 VDD.n2452 VSS 0.00207f
C9150 VDD.n2453 VSS 0.00133f
C9151 VDD.t144 VSS 3.84e-19
C9152 VDD.t329 VSS 3.65e-19
C9153 VDD.n2454 VSS 7.99e-19
C9154 VDD.n2455 VSS 0.00189f
C9155 VDD.n2456 VSS 0.00199f
C9156 VDD.n2457 VSS 0.00104f
C9157 VDD.n2458 VSS 6.26e-19
C9158 VDD.t187 VSS 9.98e-19
C9159 VDD.t758 VSS 4.23e-19
C9160 VDD.n2459 VSS 0.00203f
C9161 VDD.n2460 VSS 8.3e-19
C9162 VDD.n2461 VSS 0.00257f
C9163 VDD.n2462 VSS 1.89e-19
C9164 VDD.n2463 VSS 1.56e-19
C9165 VDD.n2464 VSS 9.17e-20
C9166 VDD.n2465 VSS 1.15e-19
C9167 VDD.n2466 VSS 2.17e-19
C9168 VDD.n2467 VSS 5.52e-19
C9169 VDD.t755 VSS 4.24e-19
C9170 VDD.n2468 VSS 0.00188f
C9171 VDD.t142 VSS 0.00127f
C9172 VDD.n2469 VSS 0.00103f
C9173 VDD.n2470 VSS 1.52e-19
C9174 VDD.n2471 VSS 1.16e-19
C9175 VDD.n2472 VSS 1.91e-19
C9176 VDD.n2473 VSS 0.00104f
C9177 VDD.t676 VSS 0.00368f
C9178 VDD.t143 VSS 0.00894f
C9179 VDD.n2474 VSS 0.00457f
C9180 VDD.n2475 VSS 7.74e-19
C9181 VDD.n2476 VSS 0.00118f
C9182 VDD.n2477 VSS 0.00196f
C9183 VDD.t327 VSS 0.00146f
C9184 VDD.t545 VSS 6.5e-19
C9185 VDD.n2478 VSS 0.00234f
C9186 VDD.n2479 VSS 0.00307f
C9187 VDD.t544 VSS 0.00377f
C9188 VDD.n2480 VSS 0.00411f
C9189 VDD.n2481 VSS 7.34e-19
C9190 VDD.n2482 VSS 6.94e-19
C9191 VDD.n2483 VSS 0.00207f
C9192 VDD.t326 VSS 0.0039f
C9193 VDD.n2484 VSS 0.00559f
C9194 VDD.n2485 VSS 7.34e-19
C9195 VDD.n2486 VSS 7.35e-19
C9196 VDD.n2487 VSS 0.00207f
C9197 VDD.n2488 VSS 0.0061f
C9198 VDD.n2489 VSS 7.34e-19
C9199 VDD.n2490 VSS 0.00125f
C9200 VDD.n2491 VSS 0.00207f
C9201 VDD.t738 VSS 0.00745f
C9202 VDD.n2492 VSS 7.34e-19
C9203 VDD.n2493 VSS 0.00125f
C9204 VDD.n2494 VSS 0.00207f
C9205 VDD.t408 VSS 0.0039f
C9206 VDD.n2495 VSS 0.00423f
C9207 VDD.n2496 VSS 7.34e-19
C9208 VDD.n2497 VSS 0.00125f
C9209 VDD.n2498 VSS 0.00207f
C9210 VDD.t319 VSS 0.0039f
C9211 VDD.n2499 VSS 0.00466f
C9212 VDD.n2500 VSS 7.34e-19
C9213 VDD.n2501 VSS 8.91e-19
C9214 VDD.n2502 VSS 0.00207f
C9215 VDD.t189 VSS 3.84e-19
C9216 VDD.t320 VSS 3.84e-19
C9217 VDD.n2503 VSS 8.11e-19
C9218 VDD.t188 VSS 0.0039f
C9219 VDD.n2504 VSS 0.00457f
C9220 VDD.n2505 VSS 7.44e-19
C9221 VDD.n2506 VSS 0.00137f
C9222 VDD.n2507 VSS 0.0017f
C9223 VDD.n2508 VSS 0.00207f
C9224 VDD.t635 VSS 0.0039f
C9225 VDD.n2509 VSS 0.00407f
C9226 VDD.n2510 VSS 7.34e-19
C9227 VDD.n2511 VSS 0.0011f
C9228 VDD.n2512 VSS 0.00207f
C9229 VDD.t546 VSS 0.0039f
C9230 VDD.n2513 VSS 0.00305f
C9231 VDD.n2514 VSS 7.34e-19
C9232 VDD.n2515 VSS 0.00105f
C9233 VDD.n2516 VSS 0.00207f
C9234 VDD.n2517 VSS 0.00703f
C9235 VDD.n2518 VSS 7.34e-19
C9236 VDD.t547 VSS 0.00176f
C9237 VDD.n2519 VSS 0.00177f
C9238 VDD.n2520 VSS 0.00195f
C9239 VDD.n2521 VSS 0.00207f
C9240 VDD.t298 VSS 0.0039f
C9241 VDD.n2522 VSS 0.00525f
C9242 VDD.n2523 VSS 7.34e-19
C9243 VDD.n2524 VSS 0.00281f
C9244 VDD.n2525 VSS 0.00207f
C9245 VDD.t315 VSS 0.0039f
C9246 VDD.n2526 VSS 0.00411f
C9247 VDD.n2527 VSS 7.34e-19
C9248 VDD.t316 VSS -3.41e-19
C9249 VDD.t299 VSS 6.16e-19
C9250 VDD.n2528 VSS 0.00241f
C9251 VDD.n2529 VSS 0.00164f
C9252 VDD.n2530 VSS 0.00125f
C9253 VDD.n2531 VSS 0.00207f
C9254 VDD.n2532 VSS 0.00622f
C9255 VDD.n2533 VSS 7.34e-19
C9256 VDD.n2534 VSS 0.0012f
C9257 VDD.n2535 VSS 0.00207f
C9258 VDD.t317 VSS 0.0039f
C9259 VDD.n2536 VSS 0.00563f
C9260 VDD.n2537 VSS 7.34e-19
C9261 VDD.n2538 VSS 0.00109f
C9262 VDD.n2539 VSS 0.00207f
C9263 VDD.t452 VSS -1.82e-19
C9264 VDD.t318 VSS 5.71e-19
C9265 VDD.n2540 VSS 0.00268f
C9266 VDD.t451 VSS 0.0039f
C9267 VDD.n2541 VSS 0.00402f
C9268 VDD.n2542 VSS 7.44e-19
C9269 VDD.n2543 VSS 0.00134f
C9270 VDD.n2544 VSS 0.00243f
C9271 VDD.n2545 VSS 0.00207f
C9272 VDD.n2546 VSS 0.00155f
C9273 VDD.n2547 VSS 0.00101f
C9274 VDD.n2548 VSS 0.00101f
C9275 VDD.n2549 VSS 7.34e-19
C9276 VDD.n2550 VSS 7.2e-19
C9277 VDD.t625 VSS 0.00385f
C9278 VDD.n2551 VSS 0.00356f
C9279 VDD.n2552 VSS 7.44e-19
C9280 VDD.n2553 VSS 0.00136f
C9281 VDD.n2554 VSS 0.00182f
C9282 VDD.n2555 VSS 0.00207f
C9283 VDD.n2556 VSS 0.0061f
C9284 VDD.n2557 VSS 7.34e-19
C9285 VDD.n2558 VSS 8.03e-19
C9286 VDD.n2559 VSS 0.00207f
C9287 VDD.t674 VSS 9.52e-19
C9288 VDD.t673 VSS 0.0039f
C9289 VDD.n2560 VSS 0.00576f
C9290 VDD.n2561 VSS 7.44e-19
C9291 VDD.n2562 VSS 0.00136f
C9292 VDD.n2563 VSS 0.00207f
C9293 VDD.n2564 VSS 0.00207f
C9294 VDD.t489 VSS 0.0039f
C9295 VDD.n2565 VSS 0.00394f
C9296 VDD.n2566 VSS 7.34e-19
C9297 VDD.n2567 VSS 0.00101f
C9298 VDD.n2568 VSS 0.00207f
C9299 VDD.t705 VSS 0.0039f
C9300 VDD.n2569 VSS 0.00356f
C9301 VDD.n2570 VSS 7.34e-19
C9302 VDD.n2571 VSS 0.00125f
C9303 VDD.n2572 VSS 0.00207f
C9304 VDD.t477 VSS 0.00724f
C9305 VDD.n2573 VSS 0.00508f
C9306 VDD.n2574 VSS 0.00128f
C9307 VDD.n2575 VSS 0.0012f
C9308 VDD.n2576 VSS 0.00207f
C9309 VDD.n2577 VSS 0.00133f
C9310 VDD.t162 VSS 3.84e-19
C9311 VDD.t478 VSS 3.65e-19
C9312 VDD.n2578 VSS 7.99e-19
C9313 VDD.n2579 VSS 0.00189f
C9314 VDD.n2580 VSS 0.00199f
C9315 VDD.n2581 VSS 0.00104f
C9316 VDD.n2582 VSS 6.26e-19
C9317 VDD.t151 VSS 9.98e-19
C9318 VDD.t754 VSS 4.23e-19
C9319 VDD.n2583 VSS 0.00203f
C9320 VDD.n2584 VSS 8.3e-19
C9321 VDD.n2585 VSS 0.00257f
C9322 VDD.n2586 VSS 1.89e-19
C9323 VDD.n2587 VSS 1.56e-19
C9324 VDD.n2588 VSS 9.17e-20
C9325 VDD.n2589 VSS 1.15e-19
C9326 VDD.n2590 VSS 2.17e-19
C9327 VDD.n2591 VSS 5.52e-19
C9328 VDD.t747 VSS 4.24e-19
C9329 VDD.n2592 VSS 0.00188f
C9330 VDD.t160 VSS 0.00127f
C9331 VDD.n2593 VSS 0.00103f
C9332 VDD.n2594 VSS 1.52e-19
C9333 VDD.n2595 VSS 1.16e-19
C9334 VDD.n2596 VSS 1.91e-19
C9335 VDD.n2597 VSS 0.00104f
C9336 VDD.t351 VSS 0.00368f
C9337 VDD.t161 VSS 0.00894f
C9338 VDD.n2598 VSS 0.00457f
C9339 VDD.n2599 VSS 7.74e-19
C9340 VDD.n2600 VSS 0.00118f
C9341 VDD.n2601 VSS 0.00196f
C9342 VDD.t480 VSS 0.00146f
C9343 VDD.t136 VSS 6.5e-19
C9344 VDD.n2602 VSS 0.00234f
C9345 VDD.n2603 VSS 0.00307f
C9346 VDD.t135 VSS 0.00377f
C9347 VDD.n2604 VSS 0.00411f
C9348 VDD.n2605 VSS 7.34e-19
C9349 VDD.n2606 VSS 6.94e-19
C9350 VDD.n2607 VSS 0.00207f
C9351 VDD.t479 VSS 0.0039f
C9352 VDD.n2608 VSS 0.00559f
C9353 VDD.n2609 VSS 7.34e-19
C9354 VDD.n2610 VSS 7.35e-19
C9355 VDD.n2611 VSS 0.00207f
C9356 VDD.n2612 VSS 0.0061f
C9357 VDD.n2613 VSS 7.34e-19
C9358 VDD.n2614 VSS 0.00125f
C9359 VDD.n2615 VSS 0.00207f
C9360 VDD.t706 VSS 0.00745f
C9361 VDD.n2616 VSS 7.34e-19
C9362 VDD.n2617 VSS 0.00125f
C9363 VDD.n2618 VSS 0.00207f
C9364 VDD.t490 VSS 0.0039f
C9365 VDD.n2619 VSS 0.00423f
C9366 VDD.n2620 VSS 7.34e-19
C9367 VDD.n2621 VSS 0.00125f
C9368 VDD.n2622 VSS 0.00207f
C9369 VDD.t335 VSS 0.0039f
C9370 VDD.n2623 VSS 0.00466f
C9371 VDD.n2624 VSS 7.34e-19
C9372 VDD.n2625 VSS 8.91e-19
C9373 VDD.n2626 VSS 0.00207f
C9374 VDD.t153 VSS 3.84e-19
C9375 VDD.t336 VSS 3.84e-19
C9376 VDD.n2627 VSS 8.11e-19
C9377 VDD.t152 VSS 0.0039f
C9378 VDD.n2628 VSS 0.00457f
C9379 VDD.n2629 VSS 7.44e-19
C9380 VDD.n2630 VSS 0.00137f
C9381 VDD.n2631 VSS 0.0017f
C9382 VDD.n2632 VSS 0.00207f
C9383 VDD.t636 VSS 0.0039f
C9384 VDD.n2633 VSS 0.00407f
C9385 VDD.n2634 VSS 7.34e-19
C9386 VDD.n2635 VSS 0.0011f
C9387 VDD.n2636 VSS 0.00207f
C9388 VDD.t133 VSS 0.0039f
C9389 VDD.n2637 VSS 0.00305f
C9390 VDD.n2638 VSS 7.34e-19
C9391 VDD.n2639 VSS 0.00105f
C9392 VDD.n2640 VSS 0.00207f
C9393 VDD.n2641 VSS 0.00703f
C9394 VDD.n2642 VSS 7.34e-19
C9395 VDD.t134 VSS 0.00176f
C9396 VDD.n2643 VSS 0.00177f
C9397 VDD.n2644 VSS 0.00195f
C9398 VDD.n2645 VSS 0.00207f
C9399 VDD.t12 VSS 0.0039f
C9400 VDD.n2646 VSS 0.00525f
C9401 VDD.n2647 VSS 7.34e-19
C9402 VDD.n2648 VSS 0.00281f
C9403 VDD.n2649 VSS 0.00207f
C9404 VDD.t333 VSS 0.0039f
C9405 VDD.n2650 VSS 0.00411f
C9406 VDD.n2651 VSS 7.34e-19
C9407 VDD.t334 VSS -3.41e-19
C9408 VDD.t13 VSS 6.16e-19
C9409 VDD.n2652 VSS 0.00241f
C9410 VDD.n2653 VSS 0.00164f
C9411 VDD.n2654 VSS 0.00125f
C9412 VDD.n2655 VSS 0.00207f
C9413 VDD.n2656 VSS 0.00622f
C9414 VDD.n2657 VSS 7.34e-19
C9415 VDD.n2658 VSS 0.0012f
C9416 VDD.n2659 VSS 0.00207f
C9417 VDD.t337 VSS 0.0039f
C9418 VDD.n2660 VSS 0.00563f
C9419 VDD.n2661 VSS 7.34e-19
C9420 VDD.n2662 VSS 0.00109f
C9421 VDD.n2663 VSS 0.00207f
C9422 VDD.t242 VSS -1.82e-19
C9423 VDD.t338 VSS 5.71e-19
C9424 VDD.n2664 VSS 0.00268f
C9425 VDD.t241 VSS 0.0039f
C9426 VDD.n2665 VSS 0.00402f
C9427 VDD.n2666 VSS 7.44e-19
C9428 VDD.n2667 VSS 0.00134f
C9429 VDD.n2668 VSS 0.00243f
C9430 VDD.n2669 VSS 0.00207f
C9431 VDD.n2670 VSS 0.00101f
C9432 VDD.t285 VSS 0.0039f
C9433 VDD.n2671 VSS 0.00994f
C9434 VDD.n2672 VSS 0.00112f
C9435 VDD.t458 VSS -1.82e-19
C9436 VDD.t263 VSS 5.71e-19
C9437 VDD.n2673 VSS 0.00268f
C9438 VDD.t457 VSS 0.00451f
C9439 VDD.n2674 VSS 0.00402f
C9440 VDD.n2675 VSS 7.44e-19
C9441 VDD.n2676 VSS 0.00134f
C9442 VDD.n2677 VSS 0.00243f
C9443 VDD.n2678 VSS 0.00484f
C9444 VDD.t262 VSS 0.0039f
C9445 VDD.n2679 VSS 0.00563f
C9446 VDD.n2680 VSS 7.34e-19
C9447 VDD.n2681 VSS 0.00109f
C9448 VDD.n2682 VSS 0.00207f
C9449 VDD.n2683 VSS 0.00622f
C9450 VDD.n2684 VSS 7.34e-19
C9451 VDD.n2685 VSS 0.0012f
C9452 VDD.n2686 VSS 0.00207f
C9453 VDD.t260 VSS 0.0039f
C9454 VDD.n2687 VSS 0.00411f
C9455 VDD.n2688 VSS 7.34e-19
C9456 VDD.t261 VSS -3.41e-19
C9457 VDD.t293 VSS 6.16e-19
C9458 VDD.n2689 VSS 0.00241f
C9459 VDD.n2690 VSS 0.00164f
C9460 VDD.n2691 VSS 0.00125f
C9461 VDD.n2692 VSS 0.00207f
C9462 VDD.t292 VSS 0.0039f
C9463 VDD.n2693 VSS 0.00525f
C9464 VDD.n2694 VSS 7.34e-19
C9465 VDD.n2695 VSS 0.00281f
C9466 VDD.n2696 VSS 0.00207f
C9467 VDD.n2697 VSS 0.00703f
C9468 VDD.n2698 VSS 7.34e-19
C9469 VDD.t472 VSS 0.00176f
C9470 VDD.n2699 VSS 0.00177f
C9471 VDD.n2700 VSS 0.00195f
C9472 VDD.n2701 VSS 0.00207f
C9473 VDD.t471 VSS 0.0039f
C9474 VDD.n2702 VSS 0.00305f
C9475 VDD.n2703 VSS 7.34e-19
C9476 VDD.n2704 VSS 0.00105f
C9477 VDD.n2705 VSS 0.00207f
C9478 VDD.t42 VSS 0.0039f
C9479 VDD.n2706 VSS 0.00407f
C9480 VDD.n2707 VSS 7.34e-19
C9481 VDD.n2708 VSS 0.0011f
C9482 VDD.n2709 VSS 0.00207f
C9483 VDD.t159 VSS 3.84e-19
C9484 VDD.t259 VSS 3.84e-19
C9485 VDD.n2710 VSS 8.11e-19
C9486 VDD.t158 VSS 0.0039f
C9487 VDD.n2711 VSS 0.00457f
C9488 VDD.n2712 VSS 7.44e-19
C9489 VDD.n2713 VSS 0.00137f
C9490 VDD.n2714 VSS 0.0017f
C9491 VDD.n2715 VSS 0.00207f
C9492 VDD.t258 VSS 0.0039f
C9493 VDD.n2716 VSS 0.00466f
C9494 VDD.n2717 VSS 7.34e-19
C9495 VDD.n2718 VSS 8.91e-19
C9496 VDD.n2719 VSS 0.00207f
C9497 VDD.t123 VSS 0.0039f
C9498 VDD.n2720 VSS 0.00423f
C9499 VDD.n2721 VSS 7.34e-19
C9500 VDD.n2722 VSS 0.00125f
C9501 VDD.n2723 VSS 0.00207f
C9502 VDD.t287 VSS 0.00745f
C9503 VDD.n2724 VSS 7.34e-19
C9504 VDD.n2725 VSS 0.00125f
C9505 VDD.n2726 VSS 0.00207f
C9506 VDD.n2727 VSS 0.0061f
C9507 VDD.n2728 VSS 7.34e-19
C9508 VDD.n2729 VSS 0.00125f
C9509 VDD.n2730 VSS 0.00207f
C9510 VDD.t540 VSS 0.0039f
C9511 VDD.n2731 VSS 0.00559f
C9512 VDD.n2732 VSS 7.34e-19
C9513 VDD.n2733 VSS 7.35e-19
C9514 VDD.n2734 VSS 0.00207f
C9515 VDD.t541 VSS 0.00146f
C9516 VDD.t470 VSS 6.5e-19
C9517 VDD.n2735 VSS 0.00234f
C9518 VDD.n2736 VSS 0.00307f
C9519 VDD.t469 VSS 0.00377f
C9520 VDD.n2737 VSS 0.00411f
C9521 VDD.n2738 VSS 7.34e-19
C9522 VDD.n2739 VSS 6.94e-19
C9523 VDD.n2740 VSS 0.00207f
C9524 VDD.t396 VSS 0.00368f
C9525 VDD.t173 VSS 0.00894f
C9526 VDD.n2741 VSS 0.00457f
C9527 VDD.n2742 VSS 7.74e-19
C9528 VDD.n2743 VSS 0.00118f
C9529 VDD.n2744 VSS 0.00196f
C9530 VDD.n2745 VSS 0.00104f
C9531 VDD.n2746 VSS 6.26e-19
C9532 VDD.t157 VSS 9.98e-19
C9533 VDD.t749 VSS 4.23e-19
C9534 VDD.n2747 VSS 0.00203f
C9535 VDD.n2748 VSS 8.3e-19
C9536 VDD.n2749 VSS 0.00257f
C9537 VDD.n2750 VSS 1.89e-19
C9538 VDD.n2751 VSS 1.56e-19
C9539 VDD.n2752 VSS 9.17e-20
C9540 VDD.n2753 VSS 1.15e-19
C9541 VDD.n2754 VSS 2.17e-19
C9542 VDD.n2755 VSS 5.52e-19
C9543 VDD.t748 VSS 4.24e-19
C9544 VDD.n2756 VSS 0.00188f
C9545 VDD.t172 VSS 0.00127f
C9546 VDD.n2757 VSS 0.00103f
C9547 VDD.n2758 VSS 1.53e-19
C9548 VDD.n2759 VSS 1.16e-19
C9549 VDD.n2760 VSS 1.91e-19
C9550 VDD.n2761 VSS 0.00104f
C9551 VDD.n2762 VSS 0.00133f
C9552 VDD.t174 VSS 3.84e-19
C9553 VDD.t543 VSS 3.65e-19
C9554 VDD.n2763 VSS 7.99e-19
C9555 VDD.n2764 VSS 0.00189f
C9556 VDD.n2765 VSS 0.00199f
C9557 VDD.t542 VSS 0.00724f
C9558 VDD.n2766 VSS 0.00508f
C9559 VDD.n2767 VSS 0.00128f
C9560 VDD.n2768 VSS 0.0012f
C9561 VDD.n2769 VSS 0.00207f
C9562 VDD.t284 VSS 0.0039f
C9563 VDD.n2770 VSS 0.00356f
C9564 VDD.n2771 VSS 7.34e-19
C9565 VDD.n2772 VSS 0.00125f
C9566 VDD.n2773 VSS 0.00207f
C9567 VDD.t124 VSS 0.0039f
C9568 VDD.n2774 VSS 0.00394f
C9569 VDD.n2775 VSS 7.34e-19
C9570 VDD.n2776 VSS 0.00101f
C9571 VDD.n2777 VSS 0.00207f
C9572 VDD.t722 VSS 9.52e-19
C9573 VDD.t721 VSS 0.0039f
C9574 VDD.n2778 VSS 0.00576f
C9575 VDD.n2779 VSS 7.44e-19
C9576 VDD.n2780 VSS 0.00136f
C9577 VDD.n2781 VSS 0.00207f
C9578 VDD.n2782 VSS 0.00207f
C9579 VDD.n2783 VSS 0.0061f
C9580 VDD.n2784 VSS 7.34e-19
C9581 VDD.n2785 VSS 8.03e-19
C9582 VDD.n2786 VSS 0.00207f
C9583 VDD.n2787 VSS 0.00122f
C9584 VDD.n2788 VSS 0.00207f
C9585 VDD.t286 VSS 4.05e-19
C9586 VDD.t690 VSS 4.05e-19
C9587 VDD.n2789 VSS 8.77e-19
C9588 VDD.n2790 VSS 0.00182f
C9589 VDD.n2791 VSS 0.00136f
C9590 VDD.n2792 VSS 7.44e-19
C9591 VDD.n2793 VSS 0.00356f
C9592 VDD.t689 VSS 0.00385f
C9593 VDD.n2794 VSS 7.34e-19
C9594 VDD.n2795 VSS 7.2e-19
C9595 VDD.n2796 VSS 0.00525f
C9596 VDD.n2797 VSS 7.34e-19
C9597 VDD.n2798 VSS 0.00101f
C9598 VDD.n2799 VSS 0.00155f
.ends

