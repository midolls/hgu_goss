magic
tech sky130A
magscale 1 2
timestamp 1699184830
<< nwell >>
rect 6688 3781 7508 3812
rect 553 3184 13468 3781
rect 504 3183 13468 3184
rect 24 2816 13468 3183
rect 553 2487 6759 2816
rect 7262 2487 13468 2816
rect 1198 2421 1416 2487
rect 1930 2424 2274 2487
rect 3142 2424 3486 2487
rect 4354 2424 4698 2487
rect 5566 2424 5910 2487
rect 6340 2439 6751 2487
rect 6340 2438 6559 2439
rect 7907 2421 8125 2487
rect 8639 2424 8983 2487
rect 9851 2424 10195 2487
rect 11063 2424 11407 2487
rect 12275 2424 12619 2487
rect 13049 2439 13460 2487
rect 13049 2438 13268 2439
rect 196 -1118 415 -1117
rect 4 -1166 415 -1118
rect 845 -1166 1189 -1103
rect 2057 -1166 2401 -1103
rect 3269 -1166 3613 -1103
rect 4481 -1166 4825 -1103
rect 5339 -1166 5557 -1100
rect 6905 -1118 7124 -1117
rect 6713 -1166 7124 -1118
rect 7554 -1166 7898 -1103
rect 8766 -1166 9110 -1103
rect 9978 -1166 10322 -1103
rect 11190 -1166 11534 -1103
rect 12048 -1166 12266 -1100
rect -4 -1495 6202 -1166
rect 6705 -1495 12911 -1166
rect -4 -1862 13440 -1495
rect -4 -1863 12960 -1862
rect -4 -2460 12911 -1863
rect 6188 -2464 6992 -2460
rect 6221 -2467 6992 -2464
<< pwell >>
rect 104 2576 290 2758
rect 294 2576 480 2758
rect 104 2572 125 2576
rect 91 2538 125 2572
rect 459 2572 480 2576
rect 459 2538 493 2572
rect 6813 2576 6999 2758
rect 7003 2576 7189 2758
rect 6813 2572 6834 2576
rect 6800 2538 6834 2572
rect 7168 2572 7189 2576
rect 7168 2538 7202 2572
rect 24 -606 13310 1820
rect 6262 -1251 6296 -1217
rect 6275 -1255 6296 -1251
rect 6630 -1251 6664 -1217
rect 6630 -1255 6651 -1251
rect 6275 -1437 6461 -1255
rect 6465 -1437 6651 -1255
rect 12971 -1251 13005 -1217
rect 12984 -1255 13005 -1251
rect 13339 -1251 13373 -1217
rect 13339 -1255 13360 -1251
rect 12984 -1437 13170 -1255
rect 13174 -1437 13360 -1255
<< nmos >>
rect 1645 2272 1675 2356
rect 2377 2272 2407 2356
rect 2499 2272 2529 2356
rect 3589 2272 3619 2356
rect 3711 2272 3741 2356
rect 4927 2272 4957 2356
rect 5049 2272 5079 2356
rect 5783 2272 5813 2356
rect 6435 2273 6465 2357
rect 6527 2273 6557 2357
rect 6623 2273 6653 2357
rect 8354 2272 8384 2356
rect 9086 2272 9116 2356
rect 9208 2272 9238 2356
rect 10298 2272 10328 2356
rect 10420 2272 10450 2356
rect 11636 2272 11666 2356
rect 11758 2272 11788 2356
rect 12492 2272 12522 2356
rect 13144 2273 13174 2357
rect 13236 2273 13266 2357
rect 13332 2273 13362 2357
rect 625 2088 655 2172
rect 697 2088 727 2172
rect 6435 2135 6465 2219
rect 7334 2088 7364 2172
rect 7406 2088 7436 2172
rect 13144 2135 13174 2219
rect 625 1950 655 2034
rect 697 1950 727 2034
rect 7334 1950 7364 2034
rect 7406 1950 7436 2034
rect 625 1812 655 1896
rect 697 1812 727 1896
rect 7334 1812 7364 1896
rect 7406 1812 7436 1896
rect 625 1674 655 1758
rect 697 1674 727 1758
rect 7334 1674 7364 1758
rect 7406 1674 7436 1758
rect 625 1536 655 1620
rect 697 1536 727 1620
rect 7334 1536 7364 1620
rect 7406 1536 7436 1620
rect 625 1398 655 1482
rect 697 1398 727 1482
rect 7334 1398 7364 1482
rect 7406 1398 7436 1482
rect 625 1260 655 1344
rect 697 1260 727 1344
rect 7334 1260 7364 1344
rect 7406 1260 7436 1344
rect 625 1122 655 1206
rect 697 1122 727 1206
rect 7334 1122 7364 1206
rect 7406 1122 7436 1206
rect 6028 115 6058 199
rect 6100 115 6130 199
rect 12737 115 12767 199
rect 12809 115 12839 199
rect 6028 -23 6058 61
rect 6100 -23 6130 61
rect 12737 -23 12767 61
rect 12809 -23 12839 61
rect 6028 -161 6058 -77
rect 6100 -161 6130 -77
rect 12737 -161 12767 -77
rect 12809 -161 12839 -77
rect 6028 -299 6058 -215
rect 6100 -299 6130 -215
rect 12737 -299 12767 -215
rect 12809 -299 12839 -215
rect 6028 -437 6058 -353
rect 6100 -437 6130 -353
rect 12737 -437 12767 -353
rect 12809 -437 12839 -353
rect 6028 -575 6058 -491
rect 6100 -575 6130 -491
rect 12737 -575 12767 -491
rect 12809 -575 12839 -491
rect 6028 -713 6058 -629
rect 6100 -713 6130 -629
rect 12737 -713 12767 -629
rect 12809 -713 12839 -629
rect 290 -898 320 -814
rect 6028 -851 6058 -767
rect 6100 -851 6130 -767
rect 6999 -898 7029 -814
rect 12737 -851 12767 -767
rect 12809 -851 12839 -767
rect 102 -1036 132 -952
rect 198 -1036 228 -952
rect 290 -1036 320 -952
rect 942 -1035 972 -951
rect 1676 -1035 1706 -951
rect 1798 -1035 1828 -951
rect 3014 -1035 3044 -951
rect 3136 -1035 3166 -951
rect 4226 -1035 4256 -951
rect 4348 -1035 4378 -951
rect 5080 -1035 5110 -951
rect 6811 -1036 6841 -952
rect 6907 -1036 6937 -952
rect 6999 -1036 7029 -952
rect 7651 -1035 7681 -951
rect 8385 -1035 8415 -951
rect 8507 -1035 8537 -951
rect 9723 -1035 9753 -951
rect 9845 -1035 9875 -951
rect 10935 -1035 10965 -951
rect 11057 -1035 11087 -951
rect 11789 -1035 11819 -951
<< scnmos >>
rect 182 2602 212 2732
rect 372 2602 402 2732
rect 6891 2602 6921 2732
rect 7081 2602 7111 2732
rect 6353 -1411 6383 -1281
rect 6543 -1411 6573 -1281
rect 13062 -1411 13092 -1281
rect 13252 -1411 13282 -1281
<< pmos >>
rect 1292 2470 1322 2554
rect 2024 2473 2054 2557
rect 2150 2473 2180 2557
rect 3236 2473 3266 2557
rect 3362 2473 3392 2557
rect 4448 2473 4478 2557
rect 4574 2473 4604 2557
rect 5660 2473 5690 2557
rect 5786 2473 5816 2557
rect 8001 2470 8031 2554
rect 8733 2473 8763 2557
rect 8859 2473 8889 2557
rect 9945 2473 9975 2557
rect 10071 2473 10101 2557
rect 11157 2473 11187 2557
rect 11283 2473 11313 2557
rect 12369 2473 12399 2557
rect 12495 2473 12525 2557
rect 939 -1236 969 -1152
rect 1065 -1236 1095 -1152
rect 2151 -1236 2181 -1152
rect 2277 -1236 2307 -1152
rect 3363 -1236 3393 -1152
rect 3489 -1236 3519 -1152
rect 4575 -1236 4605 -1152
rect 4701 -1236 4731 -1152
rect 5433 -1233 5463 -1149
rect 7648 -1236 7678 -1152
rect 7774 -1236 7804 -1152
rect 8860 -1236 8890 -1152
rect 8986 -1236 9016 -1152
rect 10072 -1236 10102 -1152
rect 10198 -1236 10228 -1152
rect 11284 -1236 11314 -1152
rect 11410 -1236 11440 -1152
rect 12142 -1233 12172 -1149
<< scpmoshvt >>
rect 182 2852 212 3052
rect 372 2852 402 3052
rect 6891 2852 6921 3052
rect 7081 2852 7111 3052
rect 6353 -1731 6383 -1531
rect 6543 -1731 6573 -1531
rect 13062 -1731 13092 -1531
rect 13252 -1731 13282 -1531
<< pmoshvt >>
rect 650 3615 680 3699
rect 7359 3615 7389 3699
rect 650 3477 680 3561
rect 7359 3477 7389 3561
rect 650 3339 680 3423
rect 7359 3339 7389 3423
rect 650 3201 680 3285
rect 7359 3201 7389 3285
rect 650 3063 680 3147
rect 7359 3063 7389 3147
rect 650 2925 680 3009
rect 7359 2925 7389 3009
rect 6435 2614 6465 2698
rect 13144 2614 13174 2698
rect 6435 2476 6465 2560
rect 6527 2476 6557 2560
rect 6623 2476 6653 2560
rect 13144 2476 13174 2560
rect 13236 2476 13266 2560
rect 13332 2476 13362 2560
rect 102 -1239 132 -1155
rect 198 -1239 228 -1155
rect 290 -1239 320 -1155
rect 6811 -1239 6841 -1155
rect 6907 -1239 6937 -1155
rect 6999 -1239 7029 -1155
rect 290 -1377 320 -1293
rect 6999 -1377 7029 -1293
rect 6075 -1688 6105 -1604
rect 12784 -1688 12814 -1604
rect 6075 -1826 6105 -1742
rect 12784 -1826 12814 -1742
rect 6075 -1964 6105 -1880
rect 12784 -1964 12814 -1880
rect 6075 -2102 6105 -2018
rect 12784 -2102 12814 -2018
rect 6075 -2240 6105 -2156
rect 12784 -2240 12814 -2156
rect 6075 -2378 6105 -2294
rect 12784 -2378 12814 -2294
<< ndiff >>
rect 130 2720 182 2732
rect 130 2686 138 2720
rect 172 2686 182 2720
rect 130 2652 182 2686
rect 130 2618 138 2652
rect 172 2618 182 2652
rect 130 2602 182 2618
rect 212 2720 264 2732
rect 212 2686 222 2720
rect 256 2686 264 2720
rect 212 2652 264 2686
rect 212 2618 222 2652
rect 256 2618 264 2652
rect 212 2602 264 2618
rect 320 2720 372 2732
rect 320 2686 328 2720
rect 362 2686 372 2720
rect 320 2652 372 2686
rect 320 2618 328 2652
rect 362 2618 372 2652
rect 320 2602 372 2618
rect 402 2720 454 2732
rect 402 2686 412 2720
rect 446 2686 454 2720
rect 6839 2720 6891 2732
rect 402 2652 454 2686
rect 402 2618 412 2652
rect 446 2618 454 2652
rect 402 2602 454 2618
rect 6839 2686 6847 2720
rect 6881 2686 6891 2720
rect 6839 2652 6891 2686
rect 6839 2618 6847 2652
rect 6881 2618 6891 2652
rect 6839 2602 6891 2618
rect 6921 2720 6973 2732
rect 6921 2686 6931 2720
rect 6965 2686 6973 2720
rect 6921 2652 6973 2686
rect 6921 2618 6931 2652
rect 6965 2618 6973 2652
rect 6921 2602 6973 2618
rect 7029 2720 7081 2732
rect 7029 2686 7037 2720
rect 7071 2686 7081 2720
rect 7029 2652 7081 2686
rect 7029 2618 7037 2652
rect 7071 2618 7081 2652
rect 7029 2602 7081 2618
rect 7111 2720 7163 2732
rect 7111 2686 7121 2720
rect 7155 2686 7163 2720
rect 7111 2652 7163 2686
rect 7111 2618 7121 2652
rect 7155 2618 7163 2652
rect 7111 2602 7163 2618
rect 1587 2344 1645 2356
rect 1587 2284 1599 2344
rect 1633 2284 1645 2344
rect 1587 2272 1645 2284
rect 1675 2344 1733 2356
rect 1675 2284 1689 2344
rect 1723 2284 1733 2344
rect 1675 2272 1733 2284
rect 2319 2344 2377 2356
rect 2319 2284 2331 2344
rect 2365 2284 2377 2344
rect 2319 2272 2377 2284
rect 2407 2344 2499 2356
rect 2407 2284 2438 2344
rect 2472 2284 2499 2344
rect 2407 2272 2499 2284
rect 2529 2344 2587 2356
rect 2529 2284 2541 2344
rect 2575 2284 2587 2344
rect 2529 2272 2587 2284
rect 3531 2344 3589 2356
rect 3531 2284 3543 2344
rect 3577 2284 3589 2344
rect 3531 2272 3589 2284
rect 3619 2344 3711 2356
rect 3619 2284 3649 2344
rect 3683 2284 3711 2344
rect 3619 2272 3711 2284
rect 3741 2344 3799 2356
rect 3741 2284 3753 2344
rect 3787 2284 3799 2344
rect 3741 2272 3799 2284
rect 4869 2344 4927 2356
rect 4869 2284 4881 2344
rect 4915 2284 4927 2344
rect 4869 2272 4927 2284
rect 4957 2344 5049 2356
rect 4957 2284 4989 2344
rect 5023 2284 5049 2344
rect 4957 2272 5049 2284
rect 5079 2344 5137 2356
rect 5079 2284 5091 2344
rect 5125 2284 5137 2344
rect 5079 2272 5137 2284
rect 5724 2344 5783 2356
rect 5724 2284 5736 2344
rect 5770 2284 5783 2344
rect 5724 2272 5783 2284
rect 5813 2344 5871 2356
rect 5813 2284 5825 2344
rect 5859 2284 5871 2344
rect 5813 2272 5871 2284
rect 6377 2345 6435 2357
rect 6377 2285 6389 2345
rect 6423 2285 6435 2345
rect 6377 2273 6435 2285
rect 6465 2345 6527 2357
rect 6465 2285 6477 2345
rect 6511 2285 6527 2345
rect 6465 2273 6527 2285
rect 6557 2345 6623 2357
rect 6557 2285 6573 2345
rect 6607 2285 6623 2345
rect 6557 2273 6623 2285
rect 6653 2345 6715 2357
rect 6653 2285 6669 2345
rect 6703 2285 6715 2345
rect 6653 2273 6715 2285
rect 8296 2344 8354 2356
rect 8296 2284 8308 2344
rect 8342 2284 8354 2344
rect 8296 2272 8354 2284
rect 8384 2344 8442 2356
rect 8384 2284 8398 2344
rect 8432 2284 8442 2344
rect 8384 2272 8442 2284
rect 9028 2344 9086 2356
rect 9028 2284 9040 2344
rect 9074 2284 9086 2344
rect 9028 2272 9086 2284
rect 9116 2344 9208 2356
rect 9116 2284 9147 2344
rect 9181 2284 9208 2344
rect 9116 2272 9208 2284
rect 9238 2344 9296 2356
rect 9238 2284 9250 2344
rect 9284 2284 9296 2344
rect 9238 2272 9296 2284
rect 10240 2344 10298 2356
rect 10240 2284 10252 2344
rect 10286 2284 10298 2344
rect 10240 2272 10298 2284
rect 10328 2344 10420 2356
rect 10328 2284 10358 2344
rect 10392 2284 10420 2344
rect 10328 2272 10420 2284
rect 10450 2344 10508 2356
rect 10450 2284 10462 2344
rect 10496 2284 10508 2344
rect 10450 2272 10508 2284
rect 11578 2344 11636 2356
rect 11578 2284 11590 2344
rect 11624 2284 11636 2344
rect 11578 2272 11636 2284
rect 11666 2344 11758 2356
rect 11666 2284 11698 2344
rect 11732 2284 11758 2344
rect 11666 2272 11758 2284
rect 11788 2344 11846 2356
rect 11788 2284 11800 2344
rect 11834 2284 11846 2344
rect 11788 2272 11846 2284
rect 12433 2344 12492 2356
rect 12433 2284 12445 2344
rect 12479 2284 12492 2344
rect 12433 2272 12492 2284
rect 12522 2344 12580 2356
rect 12522 2284 12534 2344
rect 12568 2284 12580 2344
rect 12522 2272 12580 2284
rect 13086 2345 13144 2357
rect 13086 2285 13098 2345
rect 13132 2285 13144 2345
rect 13086 2273 13144 2285
rect 13174 2345 13236 2357
rect 13174 2285 13186 2345
rect 13220 2285 13236 2345
rect 13174 2273 13236 2285
rect 13266 2345 13332 2357
rect 13266 2285 13282 2345
rect 13316 2285 13332 2345
rect 13266 2273 13332 2285
rect 13362 2345 13424 2357
rect 13362 2285 13378 2345
rect 13412 2285 13424 2345
rect 13362 2273 13424 2285
rect 6377 2207 6435 2219
rect 567 2160 625 2172
rect 567 2100 579 2160
rect 613 2100 625 2160
rect 567 2088 625 2100
rect 655 2088 697 2172
rect 727 2160 785 2172
rect 727 2100 739 2160
rect 773 2100 785 2160
rect 6377 2147 6389 2207
rect 6423 2147 6435 2207
rect 6377 2135 6435 2147
rect 6465 2207 6523 2219
rect 6465 2147 6477 2207
rect 6511 2147 6523 2207
rect 13086 2207 13144 2219
rect 6465 2135 6523 2147
rect 7276 2160 7334 2172
rect 727 2088 785 2100
rect 7276 2100 7288 2160
rect 7322 2100 7334 2160
rect 7276 2088 7334 2100
rect 7364 2088 7406 2172
rect 7436 2160 7494 2172
rect 7436 2100 7448 2160
rect 7482 2100 7494 2160
rect 13086 2147 13098 2207
rect 13132 2147 13144 2207
rect 13086 2135 13144 2147
rect 13174 2207 13232 2219
rect 13174 2147 13186 2207
rect 13220 2147 13232 2207
rect 13174 2135 13232 2147
rect 7436 2088 7494 2100
rect 567 2022 625 2034
rect 567 1962 579 2022
rect 613 1962 625 2022
rect 567 1950 625 1962
rect 655 1950 697 2034
rect 727 2022 785 2034
rect 727 1962 739 2022
rect 773 1962 785 2022
rect 727 1950 785 1962
rect 7276 2022 7334 2034
rect 7276 1962 7288 2022
rect 7322 1962 7334 2022
rect 7276 1950 7334 1962
rect 7364 1950 7406 2034
rect 7436 2022 7494 2034
rect 7436 1962 7448 2022
rect 7482 1962 7494 2022
rect 7436 1950 7494 1962
rect 567 1884 625 1896
rect 567 1824 579 1884
rect 613 1824 625 1884
rect 567 1812 625 1824
rect 655 1812 697 1896
rect 727 1884 785 1896
rect 727 1824 739 1884
rect 773 1824 785 1884
rect 727 1812 785 1824
rect 7276 1884 7334 1896
rect 7276 1824 7288 1884
rect 7322 1824 7334 1884
rect 7276 1812 7334 1824
rect 7364 1812 7406 1896
rect 7436 1884 7494 1896
rect 7436 1824 7448 1884
rect 7482 1824 7494 1884
rect 7436 1812 7494 1824
rect 567 1746 625 1758
rect 567 1686 579 1746
rect 613 1686 625 1746
rect 567 1674 625 1686
rect 655 1674 697 1758
rect 727 1746 785 1758
rect 727 1686 739 1746
rect 773 1686 785 1746
rect 727 1674 785 1686
rect 7276 1746 7334 1758
rect 7276 1686 7288 1746
rect 7322 1686 7334 1746
rect 7276 1674 7334 1686
rect 7364 1674 7406 1758
rect 7436 1746 7494 1758
rect 7436 1686 7448 1746
rect 7482 1686 7494 1746
rect 7436 1674 7494 1686
rect 567 1608 625 1620
rect 567 1548 579 1608
rect 613 1548 625 1608
rect 567 1536 625 1548
rect 655 1536 697 1620
rect 727 1608 785 1620
rect 727 1548 739 1608
rect 773 1548 785 1608
rect 727 1536 785 1548
rect 7276 1608 7334 1620
rect 7276 1548 7288 1608
rect 7322 1548 7334 1608
rect 7276 1536 7334 1548
rect 7364 1536 7406 1620
rect 7436 1608 7494 1620
rect 7436 1548 7448 1608
rect 7482 1548 7494 1608
rect 7436 1536 7494 1548
rect 567 1470 625 1482
rect 567 1410 579 1470
rect 613 1410 625 1470
rect 567 1398 625 1410
rect 655 1398 697 1482
rect 727 1470 785 1482
rect 727 1410 739 1470
rect 773 1410 785 1470
rect 727 1398 785 1410
rect 7276 1470 7334 1482
rect 7276 1410 7288 1470
rect 7322 1410 7334 1470
rect 7276 1398 7334 1410
rect 7364 1398 7406 1482
rect 7436 1470 7494 1482
rect 7436 1410 7448 1470
rect 7482 1410 7494 1470
rect 7436 1398 7494 1410
rect 567 1332 625 1344
rect 567 1272 579 1332
rect 613 1272 625 1332
rect 567 1260 625 1272
rect 655 1260 697 1344
rect 727 1332 785 1344
rect 727 1272 739 1332
rect 773 1272 785 1332
rect 727 1260 785 1272
rect 7276 1332 7334 1344
rect 7276 1272 7288 1332
rect 7322 1272 7334 1332
rect 7276 1260 7334 1272
rect 7364 1260 7406 1344
rect 7436 1332 7494 1344
rect 7436 1272 7448 1332
rect 7482 1272 7494 1332
rect 7436 1260 7494 1272
rect 567 1194 625 1206
rect 567 1134 579 1194
rect 613 1134 625 1194
rect 567 1122 625 1134
rect 655 1122 697 1206
rect 727 1194 785 1206
rect 727 1134 739 1194
rect 773 1134 785 1194
rect 7276 1194 7334 1206
rect 727 1122 785 1134
rect 7276 1134 7288 1194
rect 7322 1134 7334 1194
rect 7276 1122 7334 1134
rect 7364 1122 7406 1206
rect 7436 1194 7494 1206
rect 7436 1134 7448 1194
rect 7482 1134 7494 1194
rect 7436 1122 7494 1134
rect 5970 187 6028 199
rect 5970 127 5982 187
rect 6016 127 6028 187
rect 5970 115 6028 127
rect 6058 115 6100 199
rect 6130 187 6188 199
rect 6130 127 6142 187
rect 6176 127 6188 187
rect 12679 187 12737 199
rect 6130 115 6188 127
rect 12679 127 12691 187
rect 12725 127 12737 187
rect 12679 115 12737 127
rect 12767 115 12809 199
rect 12839 187 12897 199
rect 12839 127 12851 187
rect 12885 127 12897 187
rect 12839 115 12897 127
rect 5970 49 6028 61
rect 5970 -11 5982 49
rect 6016 -11 6028 49
rect 5970 -23 6028 -11
rect 6058 -23 6100 61
rect 6130 49 6188 61
rect 6130 -11 6142 49
rect 6176 -11 6188 49
rect 6130 -23 6188 -11
rect 12679 49 12737 61
rect 12679 -11 12691 49
rect 12725 -11 12737 49
rect 12679 -23 12737 -11
rect 12767 -23 12809 61
rect 12839 49 12897 61
rect 12839 -11 12851 49
rect 12885 -11 12897 49
rect 12839 -23 12897 -11
rect 5970 -89 6028 -77
rect 5970 -149 5982 -89
rect 6016 -149 6028 -89
rect 5970 -161 6028 -149
rect 6058 -161 6100 -77
rect 6130 -89 6188 -77
rect 6130 -149 6142 -89
rect 6176 -149 6188 -89
rect 6130 -161 6188 -149
rect 12679 -89 12737 -77
rect 12679 -149 12691 -89
rect 12725 -149 12737 -89
rect 12679 -161 12737 -149
rect 12767 -161 12809 -77
rect 12839 -89 12897 -77
rect 12839 -149 12851 -89
rect 12885 -149 12897 -89
rect 12839 -161 12897 -149
rect 5970 -227 6028 -215
rect 5970 -287 5982 -227
rect 6016 -287 6028 -227
rect 5970 -299 6028 -287
rect 6058 -299 6100 -215
rect 6130 -227 6188 -215
rect 6130 -287 6142 -227
rect 6176 -287 6188 -227
rect 6130 -299 6188 -287
rect 12679 -227 12737 -215
rect 12679 -287 12691 -227
rect 12725 -287 12737 -227
rect 12679 -299 12737 -287
rect 12767 -299 12809 -215
rect 12839 -227 12897 -215
rect 12839 -287 12851 -227
rect 12885 -287 12897 -227
rect 12839 -299 12897 -287
rect 5970 -365 6028 -353
rect 5970 -425 5982 -365
rect 6016 -425 6028 -365
rect 5970 -437 6028 -425
rect 6058 -437 6100 -353
rect 6130 -365 6188 -353
rect 6130 -425 6142 -365
rect 6176 -425 6188 -365
rect 6130 -437 6188 -425
rect 12679 -365 12737 -353
rect 12679 -425 12691 -365
rect 12725 -425 12737 -365
rect 12679 -437 12737 -425
rect 12767 -437 12809 -353
rect 12839 -365 12897 -353
rect 12839 -425 12851 -365
rect 12885 -425 12897 -365
rect 12839 -437 12897 -425
rect 5970 -503 6028 -491
rect 5970 -563 5982 -503
rect 6016 -563 6028 -503
rect 5970 -575 6028 -563
rect 6058 -575 6100 -491
rect 6130 -503 6188 -491
rect 6130 -563 6142 -503
rect 6176 -563 6188 -503
rect 6130 -575 6188 -563
rect 12679 -503 12737 -491
rect 12679 -563 12691 -503
rect 12725 -563 12737 -503
rect 12679 -575 12737 -563
rect 12767 -575 12809 -491
rect 12839 -503 12897 -491
rect 12839 -563 12851 -503
rect 12885 -563 12897 -503
rect 12839 -575 12897 -563
rect 5970 -641 6028 -629
rect 5970 -701 5982 -641
rect 6016 -701 6028 -641
rect 5970 -713 6028 -701
rect 6058 -713 6100 -629
rect 6130 -641 6188 -629
rect 6130 -701 6142 -641
rect 6176 -701 6188 -641
rect 6130 -713 6188 -701
rect 12679 -641 12737 -629
rect 12679 -701 12691 -641
rect 12725 -701 12737 -641
rect 12679 -713 12737 -701
rect 12767 -713 12809 -629
rect 12839 -641 12897 -629
rect 12839 -701 12851 -641
rect 12885 -701 12897 -641
rect 12839 -713 12897 -701
rect 5970 -779 6028 -767
rect 232 -826 290 -814
rect 232 -886 244 -826
rect 278 -886 290 -826
rect 232 -898 290 -886
rect 320 -826 378 -814
rect 320 -886 332 -826
rect 366 -886 378 -826
rect 5970 -839 5982 -779
rect 6016 -839 6028 -779
rect 5970 -851 6028 -839
rect 6058 -851 6100 -767
rect 6130 -779 6188 -767
rect 6130 -839 6142 -779
rect 6176 -839 6188 -779
rect 12679 -779 12737 -767
rect 6130 -851 6188 -839
rect 6941 -826 6999 -814
rect 320 -898 378 -886
rect 6941 -886 6953 -826
rect 6987 -886 6999 -826
rect 6941 -898 6999 -886
rect 7029 -826 7087 -814
rect 7029 -886 7041 -826
rect 7075 -886 7087 -826
rect 12679 -839 12691 -779
rect 12725 -839 12737 -779
rect 12679 -851 12737 -839
rect 12767 -851 12809 -767
rect 12839 -779 12897 -767
rect 12839 -839 12851 -779
rect 12885 -839 12897 -779
rect 12839 -851 12897 -839
rect 7029 -898 7087 -886
rect 40 -964 102 -952
rect 40 -1024 52 -964
rect 86 -1024 102 -964
rect 40 -1036 102 -1024
rect 132 -964 198 -952
rect 132 -1024 148 -964
rect 182 -1024 198 -964
rect 132 -1036 198 -1024
rect 228 -964 290 -952
rect 228 -1024 244 -964
rect 278 -1024 290 -964
rect 228 -1036 290 -1024
rect 320 -964 378 -952
rect 320 -1024 332 -964
rect 366 -1024 378 -964
rect 320 -1036 378 -1024
rect 884 -963 942 -951
rect 884 -1023 896 -963
rect 930 -1023 942 -963
rect 884 -1035 942 -1023
rect 972 -963 1031 -951
rect 972 -1023 985 -963
rect 1019 -1023 1031 -963
rect 972 -1035 1031 -1023
rect 1618 -963 1676 -951
rect 1618 -1023 1630 -963
rect 1664 -1023 1676 -963
rect 1618 -1035 1676 -1023
rect 1706 -963 1798 -951
rect 1706 -1023 1732 -963
rect 1766 -1023 1798 -963
rect 1706 -1035 1798 -1023
rect 1828 -963 1886 -951
rect 1828 -1023 1840 -963
rect 1874 -1023 1886 -963
rect 1828 -1035 1886 -1023
rect 2956 -963 3014 -951
rect 2956 -1023 2968 -963
rect 3002 -1023 3014 -963
rect 2956 -1035 3014 -1023
rect 3044 -963 3136 -951
rect 3044 -1023 3072 -963
rect 3106 -1023 3136 -963
rect 3044 -1035 3136 -1023
rect 3166 -963 3224 -951
rect 3166 -1023 3178 -963
rect 3212 -1023 3224 -963
rect 3166 -1035 3224 -1023
rect 4168 -963 4226 -951
rect 4168 -1023 4180 -963
rect 4214 -1023 4226 -963
rect 4168 -1035 4226 -1023
rect 4256 -963 4348 -951
rect 4256 -1023 4283 -963
rect 4317 -1023 4348 -963
rect 4256 -1035 4348 -1023
rect 4378 -963 4436 -951
rect 4378 -1023 4390 -963
rect 4424 -1023 4436 -963
rect 4378 -1035 4436 -1023
rect 5022 -963 5080 -951
rect 5022 -1023 5032 -963
rect 5066 -1023 5080 -963
rect 5022 -1035 5080 -1023
rect 5110 -963 5168 -951
rect 5110 -1023 5122 -963
rect 5156 -1023 5168 -963
rect 5110 -1035 5168 -1023
rect 6749 -964 6811 -952
rect 6749 -1024 6761 -964
rect 6795 -1024 6811 -964
rect 6749 -1036 6811 -1024
rect 6841 -964 6907 -952
rect 6841 -1024 6857 -964
rect 6891 -1024 6907 -964
rect 6841 -1036 6907 -1024
rect 6937 -964 6999 -952
rect 6937 -1024 6953 -964
rect 6987 -1024 6999 -964
rect 6937 -1036 6999 -1024
rect 7029 -964 7087 -952
rect 7029 -1024 7041 -964
rect 7075 -1024 7087 -964
rect 7029 -1036 7087 -1024
rect 7593 -963 7651 -951
rect 7593 -1023 7605 -963
rect 7639 -1023 7651 -963
rect 7593 -1035 7651 -1023
rect 7681 -963 7740 -951
rect 7681 -1023 7694 -963
rect 7728 -1023 7740 -963
rect 7681 -1035 7740 -1023
rect 8327 -963 8385 -951
rect 8327 -1023 8339 -963
rect 8373 -1023 8385 -963
rect 8327 -1035 8385 -1023
rect 8415 -963 8507 -951
rect 8415 -1023 8441 -963
rect 8475 -1023 8507 -963
rect 8415 -1035 8507 -1023
rect 8537 -963 8595 -951
rect 8537 -1023 8549 -963
rect 8583 -1023 8595 -963
rect 8537 -1035 8595 -1023
rect 9665 -963 9723 -951
rect 9665 -1023 9677 -963
rect 9711 -1023 9723 -963
rect 9665 -1035 9723 -1023
rect 9753 -963 9845 -951
rect 9753 -1023 9781 -963
rect 9815 -1023 9845 -963
rect 9753 -1035 9845 -1023
rect 9875 -963 9933 -951
rect 9875 -1023 9887 -963
rect 9921 -1023 9933 -963
rect 9875 -1035 9933 -1023
rect 10877 -963 10935 -951
rect 10877 -1023 10889 -963
rect 10923 -1023 10935 -963
rect 10877 -1035 10935 -1023
rect 10965 -963 11057 -951
rect 10965 -1023 10992 -963
rect 11026 -1023 11057 -963
rect 10965 -1035 11057 -1023
rect 11087 -963 11145 -951
rect 11087 -1023 11099 -963
rect 11133 -1023 11145 -963
rect 11087 -1035 11145 -1023
rect 11731 -963 11789 -951
rect 11731 -1023 11741 -963
rect 11775 -1023 11789 -963
rect 11731 -1035 11789 -1023
rect 11819 -963 11877 -951
rect 11819 -1023 11831 -963
rect 11865 -1023 11877 -963
rect 11819 -1035 11877 -1023
rect 6301 -1297 6353 -1281
rect 6301 -1331 6309 -1297
rect 6343 -1331 6353 -1297
rect 6301 -1365 6353 -1331
rect 6301 -1399 6309 -1365
rect 6343 -1399 6353 -1365
rect 6301 -1411 6353 -1399
rect 6383 -1297 6435 -1281
rect 6383 -1331 6393 -1297
rect 6427 -1331 6435 -1297
rect 6383 -1365 6435 -1331
rect 6383 -1399 6393 -1365
rect 6427 -1399 6435 -1365
rect 6383 -1411 6435 -1399
rect 6491 -1297 6543 -1281
rect 6491 -1331 6499 -1297
rect 6533 -1331 6543 -1297
rect 6491 -1365 6543 -1331
rect 6491 -1399 6499 -1365
rect 6533 -1399 6543 -1365
rect 6491 -1411 6543 -1399
rect 6573 -1297 6625 -1281
rect 6573 -1331 6583 -1297
rect 6617 -1331 6625 -1297
rect 6573 -1365 6625 -1331
rect 6573 -1399 6583 -1365
rect 6617 -1399 6625 -1365
rect 13010 -1297 13062 -1281
rect 13010 -1331 13018 -1297
rect 13052 -1331 13062 -1297
rect 13010 -1365 13062 -1331
rect 6573 -1411 6625 -1399
rect 13010 -1399 13018 -1365
rect 13052 -1399 13062 -1365
rect 13010 -1411 13062 -1399
rect 13092 -1297 13144 -1281
rect 13092 -1331 13102 -1297
rect 13136 -1331 13144 -1297
rect 13092 -1365 13144 -1331
rect 13092 -1399 13102 -1365
rect 13136 -1399 13144 -1365
rect 13092 -1411 13144 -1399
rect 13200 -1297 13252 -1281
rect 13200 -1331 13208 -1297
rect 13242 -1331 13252 -1297
rect 13200 -1365 13252 -1331
rect 13200 -1399 13208 -1365
rect 13242 -1399 13252 -1365
rect 13200 -1411 13252 -1399
rect 13282 -1297 13334 -1281
rect 13282 -1331 13292 -1297
rect 13326 -1331 13334 -1297
rect 13282 -1365 13334 -1331
rect 13282 -1399 13292 -1365
rect 13326 -1399 13334 -1365
rect 13282 -1411 13334 -1399
<< pdiff >>
rect 592 3687 650 3699
rect 592 3627 604 3687
rect 638 3627 650 3687
rect 592 3615 650 3627
rect 680 3687 738 3699
rect 680 3627 692 3687
rect 726 3627 738 3687
rect 680 3615 738 3627
rect 7301 3687 7359 3699
rect 7301 3627 7313 3687
rect 7347 3627 7359 3687
rect 7301 3615 7359 3627
rect 7389 3687 7447 3699
rect 7389 3627 7401 3687
rect 7435 3627 7447 3687
rect 7389 3615 7447 3627
rect 592 3549 650 3561
rect 592 3489 604 3549
rect 638 3489 650 3549
rect 592 3477 650 3489
rect 680 3549 738 3561
rect 680 3489 692 3549
rect 726 3489 738 3549
rect 680 3477 738 3489
rect 7301 3549 7359 3561
rect 7301 3489 7313 3549
rect 7347 3489 7359 3549
rect 7301 3477 7359 3489
rect 7389 3549 7447 3561
rect 7389 3489 7401 3549
rect 7435 3489 7447 3549
rect 7389 3477 7447 3489
rect 592 3411 650 3423
rect 592 3351 604 3411
rect 638 3351 650 3411
rect 592 3339 650 3351
rect 680 3411 738 3423
rect 680 3351 692 3411
rect 726 3351 738 3411
rect 7301 3411 7359 3423
rect 680 3339 738 3351
rect 7301 3351 7313 3411
rect 7347 3351 7359 3411
rect 7301 3339 7359 3351
rect 7389 3411 7447 3423
rect 7389 3351 7401 3411
rect 7435 3351 7447 3411
rect 7389 3339 7447 3351
rect 592 3273 650 3285
rect 592 3213 604 3273
rect 638 3213 650 3273
rect 592 3201 650 3213
rect 680 3273 738 3285
rect 680 3213 692 3273
rect 726 3213 738 3273
rect 7301 3273 7359 3285
rect 680 3201 738 3213
rect 7301 3213 7313 3273
rect 7347 3213 7359 3273
rect 7301 3201 7359 3213
rect 7389 3273 7447 3285
rect 7389 3213 7401 3273
rect 7435 3213 7447 3273
rect 7389 3201 7447 3213
rect 592 3135 650 3147
rect 592 3075 604 3135
rect 638 3075 650 3135
rect 592 3063 650 3075
rect 680 3135 738 3147
rect 680 3075 692 3135
rect 726 3075 738 3135
rect 7301 3135 7359 3147
rect 680 3063 738 3075
rect 130 3040 182 3052
rect 130 3006 138 3040
rect 172 3006 182 3040
rect 130 2972 182 3006
rect 130 2938 138 2972
rect 172 2938 182 2972
rect 130 2904 182 2938
rect 130 2870 138 2904
rect 172 2870 182 2904
rect 130 2852 182 2870
rect 212 3040 264 3052
rect 212 3006 222 3040
rect 256 3006 264 3040
rect 212 2972 264 3006
rect 212 2938 222 2972
rect 256 2938 264 2972
rect 212 2904 264 2938
rect 212 2870 222 2904
rect 256 2870 264 2904
rect 212 2852 264 2870
rect 320 3040 372 3052
rect 320 3006 328 3040
rect 362 3006 372 3040
rect 320 2972 372 3006
rect 320 2938 328 2972
rect 362 2938 372 2972
rect 320 2904 372 2938
rect 320 2870 328 2904
rect 362 2870 372 2904
rect 320 2852 372 2870
rect 402 3040 454 3052
rect 402 3006 412 3040
rect 446 3006 454 3040
rect 7301 3075 7313 3135
rect 7347 3075 7359 3135
rect 7301 3063 7359 3075
rect 7389 3135 7447 3147
rect 7389 3075 7401 3135
rect 7435 3075 7447 3135
rect 7389 3063 7447 3075
rect 402 2972 454 3006
rect 402 2938 412 2972
rect 446 2938 454 2972
rect 402 2904 454 2938
rect 592 2997 650 3009
rect 592 2937 604 2997
rect 638 2937 650 2997
rect 592 2925 650 2937
rect 680 2997 738 3009
rect 680 2937 692 2997
rect 726 2937 738 2997
rect 6839 3040 6891 3052
rect 6839 3006 6847 3040
rect 6881 3006 6891 3040
rect 680 2925 738 2937
rect 6839 2972 6891 3006
rect 6839 2938 6847 2972
rect 6881 2938 6891 2972
rect 402 2870 412 2904
rect 446 2870 454 2904
rect 6839 2904 6891 2938
rect 402 2852 454 2870
rect 6839 2870 6847 2904
rect 6881 2870 6891 2904
rect 6839 2852 6891 2870
rect 6921 3040 6973 3052
rect 6921 3006 6931 3040
rect 6965 3006 6973 3040
rect 6921 2972 6973 3006
rect 6921 2938 6931 2972
rect 6965 2938 6973 2972
rect 6921 2904 6973 2938
rect 6921 2870 6931 2904
rect 6965 2870 6973 2904
rect 6921 2852 6973 2870
rect 7029 3040 7081 3052
rect 7029 3006 7037 3040
rect 7071 3006 7081 3040
rect 7029 2972 7081 3006
rect 7029 2938 7037 2972
rect 7071 2938 7081 2972
rect 7029 2904 7081 2938
rect 7029 2870 7037 2904
rect 7071 2870 7081 2904
rect 7029 2852 7081 2870
rect 7111 3040 7163 3052
rect 7111 3006 7121 3040
rect 7155 3006 7163 3040
rect 7111 2972 7163 3006
rect 7111 2938 7121 2972
rect 7155 2938 7163 2972
rect 7111 2904 7163 2938
rect 7301 2997 7359 3009
rect 7301 2937 7313 2997
rect 7347 2937 7359 2997
rect 7301 2925 7359 2937
rect 7389 2997 7447 3009
rect 7389 2937 7401 2997
rect 7435 2937 7447 2997
rect 7389 2925 7447 2937
rect 7111 2870 7121 2904
rect 7155 2870 7163 2904
rect 7111 2852 7163 2870
rect 6377 2686 6435 2698
rect 6377 2626 6389 2686
rect 6423 2626 6435 2686
rect 6377 2614 6435 2626
rect 6465 2686 6523 2698
rect 6465 2626 6477 2686
rect 6511 2626 6523 2686
rect 6465 2614 6523 2626
rect 13086 2686 13144 2698
rect 13086 2626 13098 2686
rect 13132 2626 13144 2686
rect 13086 2614 13144 2626
rect 13174 2686 13232 2698
rect 13174 2626 13186 2686
rect 13220 2626 13232 2686
rect 13174 2614 13232 2626
rect 1234 2542 1292 2554
rect 1234 2482 1246 2542
rect 1280 2482 1292 2542
rect 1234 2470 1292 2482
rect 1322 2545 1380 2554
rect 1322 2485 1334 2545
rect 1368 2485 1380 2545
rect 1322 2470 1380 2485
rect 1966 2545 2024 2557
rect 1966 2485 1978 2545
rect 2012 2485 2024 2545
rect 1966 2473 2024 2485
rect 2054 2545 2150 2557
rect 2054 2485 2083 2545
rect 2117 2485 2150 2545
rect 2054 2473 2150 2485
rect 2180 2545 2238 2557
rect 2180 2485 2192 2545
rect 2226 2485 2238 2545
rect 2180 2473 2238 2485
rect 3178 2545 3236 2557
rect 3178 2485 3190 2545
rect 3224 2485 3236 2545
rect 3178 2473 3236 2485
rect 3266 2545 3362 2557
rect 3266 2485 3294 2545
rect 3328 2485 3362 2545
rect 3266 2473 3362 2485
rect 3392 2545 3450 2557
rect 3392 2485 3404 2545
rect 3438 2485 3450 2545
rect 3392 2473 3450 2485
rect 4390 2545 4448 2557
rect 4390 2485 4402 2545
rect 4436 2485 4448 2545
rect 4390 2473 4448 2485
rect 4478 2545 4574 2557
rect 4478 2485 4507 2545
rect 4541 2485 4574 2545
rect 4478 2473 4574 2485
rect 4604 2545 4662 2557
rect 4604 2485 4616 2545
rect 4650 2485 4662 2545
rect 4604 2473 4662 2485
rect 5602 2545 5660 2557
rect 5602 2485 5614 2545
rect 5648 2485 5660 2545
rect 5602 2473 5660 2485
rect 5690 2545 5786 2557
rect 5690 2485 5721 2545
rect 5755 2485 5786 2545
rect 5690 2473 5786 2485
rect 5816 2545 5874 2557
rect 5816 2485 5828 2545
rect 5862 2485 5874 2545
rect 5816 2473 5874 2485
rect 6377 2548 6435 2560
rect 6377 2488 6389 2548
rect 6423 2488 6435 2548
rect 6377 2476 6435 2488
rect 6465 2548 6527 2560
rect 6465 2488 6477 2548
rect 6511 2488 6527 2548
rect 6465 2476 6527 2488
rect 6557 2548 6623 2560
rect 6557 2488 6573 2548
rect 6607 2488 6623 2548
rect 6557 2476 6623 2488
rect 6653 2548 6715 2560
rect 6653 2488 6669 2548
rect 6703 2488 6715 2548
rect 7943 2542 8001 2554
rect 6653 2476 6715 2488
rect 7943 2482 7955 2542
rect 7989 2482 8001 2542
rect 7943 2470 8001 2482
rect 8031 2545 8089 2554
rect 8031 2485 8043 2545
rect 8077 2485 8089 2545
rect 8031 2470 8089 2485
rect 8675 2545 8733 2557
rect 8675 2485 8687 2545
rect 8721 2485 8733 2545
rect 8675 2473 8733 2485
rect 8763 2545 8859 2557
rect 8763 2485 8792 2545
rect 8826 2485 8859 2545
rect 8763 2473 8859 2485
rect 8889 2545 8947 2557
rect 8889 2485 8901 2545
rect 8935 2485 8947 2545
rect 8889 2473 8947 2485
rect 9887 2545 9945 2557
rect 9887 2485 9899 2545
rect 9933 2485 9945 2545
rect 9887 2473 9945 2485
rect 9975 2545 10071 2557
rect 9975 2485 10003 2545
rect 10037 2485 10071 2545
rect 9975 2473 10071 2485
rect 10101 2545 10159 2557
rect 10101 2485 10113 2545
rect 10147 2485 10159 2545
rect 10101 2473 10159 2485
rect 11099 2545 11157 2557
rect 11099 2485 11111 2545
rect 11145 2485 11157 2545
rect 11099 2473 11157 2485
rect 11187 2545 11283 2557
rect 11187 2485 11216 2545
rect 11250 2485 11283 2545
rect 11187 2473 11283 2485
rect 11313 2545 11371 2557
rect 11313 2485 11325 2545
rect 11359 2485 11371 2545
rect 11313 2473 11371 2485
rect 12311 2545 12369 2557
rect 12311 2485 12323 2545
rect 12357 2485 12369 2545
rect 12311 2473 12369 2485
rect 12399 2545 12495 2557
rect 12399 2485 12430 2545
rect 12464 2485 12495 2545
rect 12399 2473 12495 2485
rect 12525 2545 12583 2557
rect 12525 2485 12537 2545
rect 12571 2485 12583 2545
rect 12525 2473 12583 2485
rect 13086 2548 13144 2560
rect 13086 2488 13098 2548
rect 13132 2488 13144 2548
rect 13086 2476 13144 2488
rect 13174 2548 13236 2560
rect 13174 2488 13186 2548
rect 13220 2488 13236 2548
rect 13174 2476 13236 2488
rect 13266 2548 13332 2560
rect 13266 2488 13282 2548
rect 13316 2488 13332 2548
rect 13266 2476 13332 2488
rect 13362 2548 13424 2560
rect 13362 2488 13378 2548
rect 13412 2488 13424 2548
rect 13362 2476 13424 2488
rect 40 -1167 102 -1155
rect 40 -1227 52 -1167
rect 86 -1227 102 -1167
rect 40 -1239 102 -1227
rect 132 -1167 198 -1155
rect 132 -1227 148 -1167
rect 182 -1227 198 -1167
rect 132 -1239 198 -1227
rect 228 -1167 290 -1155
rect 228 -1227 244 -1167
rect 278 -1227 290 -1167
rect 228 -1239 290 -1227
rect 320 -1167 378 -1155
rect 320 -1227 332 -1167
rect 366 -1227 378 -1167
rect 320 -1239 378 -1227
rect 881 -1164 939 -1152
rect 881 -1224 893 -1164
rect 927 -1224 939 -1164
rect 881 -1236 939 -1224
rect 969 -1164 1065 -1152
rect 969 -1224 1000 -1164
rect 1034 -1224 1065 -1164
rect 969 -1236 1065 -1224
rect 1095 -1164 1153 -1152
rect 1095 -1224 1107 -1164
rect 1141 -1224 1153 -1164
rect 1095 -1236 1153 -1224
rect 2093 -1164 2151 -1152
rect 2093 -1224 2105 -1164
rect 2139 -1224 2151 -1164
rect 2093 -1236 2151 -1224
rect 2181 -1164 2277 -1152
rect 2181 -1224 2214 -1164
rect 2248 -1224 2277 -1164
rect 2181 -1236 2277 -1224
rect 2307 -1164 2365 -1152
rect 2307 -1224 2319 -1164
rect 2353 -1224 2365 -1164
rect 2307 -1236 2365 -1224
rect 3305 -1164 3363 -1152
rect 3305 -1224 3317 -1164
rect 3351 -1224 3363 -1164
rect 3305 -1236 3363 -1224
rect 3393 -1164 3489 -1152
rect 3393 -1224 3427 -1164
rect 3461 -1224 3489 -1164
rect 3393 -1236 3489 -1224
rect 3519 -1164 3577 -1152
rect 3519 -1224 3531 -1164
rect 3565 -1224 3577 -1164
rect 3519 -1236 3577 -1224
rect 4517 -1164 4575 -1152
rect 4517 -1224 4529 -1164
rect 4563 -1224 4575 -1164
rect 4517 -1236 4575 -1224
rect 4605 -1164 4701 -1152
rect 4605 -1224 4638 -1164
rect 4672 -1224 4701 -1164
rect 4605 -1236 4701 -1224
rect 4731 -1164 4789 -1152
rect 4731 -1224 4743 -1164
rect 4777 -1224 4789 -1164
rect 4731 -1236 4789 -1224
rect 5375 -1164 5433 -1149
rect 5375 -1224 5387 -1164
rect 5421 -1224 5433 -1164
rect 5375 -1233 5433 -1224
rect 5463 -1161 5521 -1149
rect 5463 -1221 5475 -1161
rect 5509 -1221 5521 -1161
rect 6749 -1167 6811 -1155
rect 5463 -1233 5521 -1221
rect 6749 -1227 6761 -1167
rect 6795 -1227 6811 -1167
rect 6749 -1239 6811 -1227
rect 6841 -1167 6907 -1155
rect 6841 -1227 6857 -1167
rect 6891 -1227 6907 -1167
rect 6841 -1239 6907 -1227
rect 6937 -1167 6999 -1155
rect 6937 -1227 6953 -1167
rect 6987 -1227 6999 -1167
rect 6937 -1239 6999 -1227
rect 7029 -1167 7087 -1155
rect 7029 -1227 7041 -1167
rect 7075 -1227 7087 -1167
rect 7029 -1239 7087 -1227
rect 7590 -1164 7648 -1152
rect 7590 -1224 7602 -1164
rect 7636 -1224 7648 -1164
rect 7590 -1236 7648 -1224
rect 7678 -1164 7774 -1152
rect 7678 -1224 7709 -1164
rect 7743 -1224 7774 -1164
rect 7678 -1236 7774 -1224
rect 7804 -1164 7862 -1152
rect 7804 -1224 7816 -1164
rect 7850 -1224 7862 -1164
rect 7804 -1236 7862 -1224
rect 8802 -1164 8860 -1152
rect 8802 -1224 8814 -1164
rect 8848 -1224 8860 -1164
rect 8802 -1236 8860 -1224
rect 8890 -1164 8986 -1152
rect 8890 -1224 8923 -1164
rect 8957 -1224 8986 -1164
rect 8890 -1236 8986 -1224
rect 9016 -1164 9074 -1152
rect 9016 -1224 9028 -1164
rect 9062 -1224 9074 -1164
rect 9016 -1236 9074 -1224
rect 10014 -1164 10072 -1152
rect 10014 -1224 10026 -1164
rect 10060 -1224 10072 -1164
rect 10014 -1236 10072 -1224
rect 10102 -1164 10198 -1152
rect 10102 -1224 10136 -1164
rect 10170 -1224 10198 -1164
rect 10102 -1236 10198 -1224
rect 10228 -1164 10286 -1152
rect 10228 -1224 10240 -1164
rect 10274 -1224 10286 -1164
rect 10228 -1236 10286 -1224
rect 11226 -1164 11284 -1152
rect 11226 -1224 11238 -1164
rect 11272 -1224 11284 -1164
rect 11226 -1236 11284 -1224
rect 11314 -1164 11410 -1152
rect 11314 -1224 11347 -1164
rect 11381 -1224 11410 -1164
rect 11314 -1236 11410 -1224
rect 11440 -1164 11498 -1152
rect 11440 -1224 11452 -1164
rect 11486 -1224 11498 -1164
rect 11440 -1236 11498 -1224
rect 12084 -1164 12142 -1149
rect 12084 -1224 12096 -1164
rect 12130 -1224 12142 -1164
rect 12084 -1233 12142 -1224
rect 12172 -1161 12230 -1149
rect 12172 -1221 12184 -1161
rect 12218 -1221 12230 -1161
rect 12172 -1233 12230 -1221
rect 232 -1305 290 -1293
rect 232 -1365 244 -1305
rect 278 -1365 290 -1305
rect 232 -1377 290 -1365
rect 320 -1305 378 -1293
rect 320 -1365 332 -1305
rect 366 -1365 378 -1305
rect 320 -1377 378 -1365
rect 6941 -1305 6999 -1293
rect 6941 -1365 6953 -1305
rect 6987 -1365 6999 -1305
rect 6941 -1377 6999 -1365
rect 7029 -1305 7087 -1293
rect 7029 -1365 7041 -1305
rect 7075 -1365 7087 -1305
rect 7029 -1377 7087 -1365
rect 6301 -1549 6353 -1531
rect 6301 -1583 6309 -1549
rect 6343 -1583 6353 -1549
rect 6017 -1616 6075 -1604
rect 6017 -1676 6029 -1616
rect 6063 -1676 6075 -1616
rect 6017 -1688 6075 -1676
rect 6105 -1616 6163 -1604
rect 6105 -1676 6117 -1616
rect 6151 -1676 6163 -1616
rect 6105 -1688 6163 -1676
rect 6301 -1617 6353 -1583
rect 6301 -1651 6309 -1617
rect 6343 -1651 6353 -1617
rect 6301 -1685 6353 -1651
rect 6301 -1719 6309 -1685
rect 6343 -1719 6353 -1685
rect 6301 -1731 6353 -1719
rect 6383 -1549 6435 -1531
rect 6383 -1583 6393 -1549
rect 6427 -1583 6435 -1549
rect 6383 -1617 6435 -1583
rect 6383 -1651 6393 -1617
rect 6427 -1651 6435 -1617
rect 6383 -1685 6435 -1651
rect 6383 -1719 6393 -1685
rect 6427 -1719 6435 -1685
rect 6383 -1731 6435 -1719
rect 6491 -1549 6543 -1531
rect 6491 -1583 6499 -1549
rect 6533 -1583 6543 -1549
rect 6491 -1617 6543 -1583
rect 6491 -1651 6499 -1617
rect 6533 -1651 6543 -1617
rect 6491 -1685 6543 -1651
rect 6491 -1719 6499 -1685
rect 6533 -1719 6543 -1685
rect 6491 -1731 6543 -1719
rect 6573 -1549 6625 -1531
rect 6573 -1583 6583 -1549
rect 6617 -1583 6625 -1549
rect 13010 -1549 13062 -1531
rect 6573 -1617 6625 -1583
rect 13010 -1583 13018 -1549
rect 13052 -1583 13062 -1549
rect 6573 -1651 6583 -1617
rect 6617 -1651 6625 -1617
rect 6573 -1685 6625 -1651
rect 12726 -1616 12784 -1604
rect 6573 -1719 6583 -1685
rect 6617 -1719 6625 -1685
rect 6573 -1731 6625 -1719
rect 12726 -1676 12738 -1616
rect 12772 -1676 12784 -1616
rect 12726 -1688 12784 -1676
rect 12814 -1616 12872 -1604
rect 12814 -1676 12826 -1616
rect 12860 -1676 12872 -1616
rect 12814 -1688 12872 -1676
rect 13010 -1617 13062 -1583
rect 13010 -1651 13018 -1617
rect 13052 -1651 13062 -1617
rect 13010 -1685 13062 -1651
rect 6017 -1754 6075 -1742
rect 6017 -1814 6029 -1754
rect 6063 -1814 6075 -1754
rect 6017 -1826 6075 -1814
rect 6105 -1754 6163 -1742
rect 6105 -1814 6117 -1754
rect 6151 -1814 6163 -1754
rect 13010 -1719 13018 -1685
rect 13052 -1719 13062 -1685
rect 13010 -1731 13062 -1719
rect 13092 -1549 13144 -1531
rect 13092 -1583 13102 -1549
rect 13136 -1583 13144 -1549
rect 13092 -1617 13144 -1583
rect 13092 -1651 13102 -1617
rect 13136 -1651 13144 -1617
rect 13092 -1685 13144 -1651
rect 13092 -1719 13102 -1685
rect 13136 -1719 13144 -1685
rect 13092 -1731 13144 -1719
rect 13200 -1549 13252 -1531
rect 13200 -1583 13208 -1549
rect 13242 -1583 13252 -1549
rect 13200 -1617 13252 -1583
rect 13200 -1651 13208 -1617
rect 13242 -1651 13252 -1617
rect 13200 -1685 13252 -1651
rect 13200 -1719 13208 -1685
rect 13242 -1719 13252 -1685
rect 13200 -1731 13252 -1719
rect 13282 -1549 13334 -1531
rect 13282 -1583 13292 -1549
rect 13326 -1583 13334 -1549
rect 13282 -1617 13334 -1583
rect 13282 -1651 13292 -1617
rect 13326 -1651 13334 -1617
rect 13282 -1685 13334 -1651
rect 13282 -1719 13292 -1685
rect 13326 -1719 13334 -1685
rect 13282 -1731 13334 -1719
rect 12726 -1754 12784 -1742
rect 6105 -1826 6163 -1814
rect 12726 -1814 12738 -1754
rect 12772 -1814 12784 -1754
rect 12726 -1826 12784 -1814
rect 12814 -1754 12872 -1742
rect 12814 -1814 12826 -1754
rect 12860 -1814 12872 -1754
rect 12814 -1826 12872 -1814
rect 6017 -1892 6075 -1880
rect 6017 -1952 6029 -1892
rect 6063 -1952 6075 -1892
rect 6017 -1964 6075 -1952
rect 6105 -1892 6163 -1880
rect 6105 -1952 6117 -1892
rect 6151 -1952 6163 -1892
rect 6105 -1964 6163 -1952
rect 12726 -1892 12784 -1880
rect 12726 -1952 12738 -1892
rect 12772 -1952 12784 -1892
rect 12726 -1964 12784 -1952
rect 12814 -1892 12872 -1880
rect 12814 -1952 12826 -1892
rect 12860 -1952 12872 -1892
rect 12814 -1964 12872 -1952
rect 6017 -2030 6075 -2018
rect 6017 -2090 6029 -2030
rect 6063 -2090 6075 -2030
rect 6017 -2102 6075 -2090
rect 6105 -2030 6163 -2018
rect 6105 -2090 6117 -2030
rect 6151 -2090 6163 -2030
rect 12726 -2030 12784 -2018
rect 6105 -2102 6163 -2090
rect 12726 -2090 12738 -2030
rect 12772 -2090 12784 -2030
rect 12726 -2102 12784 -2090
rect 12814 -2030 12872 -2018
rect 12814 -2090 12826 -2030
rect 12860 -2090 12872 -2030
rect 12814 -2102 12872 -2090
rect 6017 -2168 6075 -2156
rect 6017 -2228 6029 -2168
rect 6063 -2228 6075 -2168
rect 6017 -2240 6075 -2228
rect 6105 -2168 6163 -2156
rect 6105 -2228 6117 -2168
rect 6151 -2228 6163 -2168
rect 6105 -2240 6163 -2228
rect 12726 -2168 12784 -2156
rect 12726 -2228 12738 -2168
rect 12772 -2228 12784 -2168
rect 12726 -2240 12784 -2228
rect 12814 -2168 12872 -2156
rect 12814 -2228 12826 -2168
rect 12860 -2228 12872 -2168
rect 12814 -2240 12872 -2228
rect 6017 -2306 6075 -2294
rect 6017 -2366 6029 -2306
rect 6063 -2366 6075 -2306
rect 6017 -2378 6075 -2366
rect 6105 -2306 6163 -2294
rect 6105 -2366 6117 -2306
rect 6151 -2366 6163 -2306
rect 12726 -2306 12784 -2294
rect 6105 -2378 6163 -2366
rect 12726 -2366 12738 -2306
rect 12772 -2366 12784 -2306
rect 12726 -2378 12784 -2366
rect 12814 -2306 12872 -2294
rect 12814 -2366 12826 -2306
rect 12860 -2366 12872 -2306
rect 12814 -2378 12872 -2366
<< ndiffc >>
rect 138 2686 172 2720
rect 138 2618 172 2652
rect 222 2686 256 2720
rect 222 2618 256 2652
rect 328 2686 362 2720
rect 328 2618 362 2652
rect 412 2686 446 2720
rect 412 2618 446 2652
rect 6847 2686 6881 2720
rect 6847 2618 6881 2652
rect 6931 2686 6965 2720
rect 6931 2618 6965 2652
rect 7037 2686 7071 2720
rect 7037 2618 7071 2652
rect 7121 2686 7155 2720
rect 7121 2618 7155 2652
rect 1599 2284 1633 2344
rect 1689 2284 1723 2344
rect 2331 2284 2365 2344
rect 2438 2284 2472 2344
rect 2541 2284 2575 2344
rect 3543 2284 3577 2344
rect 3649 2284 3683 2344
rect 3753 2284 3787 2344
rect 4881 2284 4915 2344
rect 4989 2284 5023 2344
rect 5091 2284 5125 2344
rect 5736 2284 5770 2344
rect 5825 2284 5859 2344
rect 6389 2285 6423 2345
rect 6477 2285 6511 2345
rect 6573 2285 6607 2345
rect 6669 2285 6703 2345
rect 8308 2284 8342 2344
rect 8398 2284 8432 2344
rect 9040 2284 9074 2344
rect 9147 2284 9181 2344
rect 9250 2284 9284 2344
rect 10252 2284 10286 2344
rect 10358 2284 10392 2344
rect 10462 2284 10496 2344
rect 11590 2284 11624 2344
rect 11698 2284 11732 2344
rect 11800 2284 11834 2344
rect 12445 2284 12479 2344
rect 12534 2284 12568 2344
rect 13098 2285 13132 2345
rect 13186 2285 13220 2345
rect 13282 2285 13316 2345
rect 13378 2285 13412 2345
rect 579 2100 613 2160
rect 739 2100 773 2160
rect 6389 2147 6423 2207
rect 6477 2147 6511 2207
rect 7288 2100 7322 2160
rect 7448 2100 7482 2160
rect 13098 2147 13132 2207
rect 13186 2147 13220 2207
rect 579 1962 613 2022
rect 739 1962 773 2022
rect 7288 1962 7322 2022
rect 7448 1962 7482 2022
rect 579 1824 613 1884
rect 739 1824 773 1884
rect 7288 1824 7322 1884
rect 7448 1824 7482 1884
rect 579 1686 613 1746
rect 739 1686 773 1746
rect 7288 1686 7322 1746
rect 7448 1686 7482 1746
rect 579 1548 613 1608
rect 739 1548 773 1608
rect 7288 1548 7322 1608
rect 7448 1548 7482 1608
rect 579 1410 613 1470
rect 739 1410 773 1470
rect 7288 1410 7322 1470
rect 7448 1410 7482 1470
rect 579 1272 613 1332
rect 739 1272 773 1332
rect 7288 1272 7322 1332
rect 7448 1272 7482 1332
rect 579 1134 613 1194
rect 739 1134 773 1194
rect 7288 1134 7322 1194
rect 7448 1134 7482 1194
rect 5982 127 6016 187
rect 6142 127 6176 187
rect 12691 127 12725 187
rect 12851 127 12885 187
rect 5982 -11 6016 49
rect 6142 -11 6176 49
rect 12691 -11 12725 49
rect 12851 -11 12885 49
rect 5982 -149 6016 -89
rect 6142 -149 6176 -89
rect 12691 -149 12725 -89
rect 12851 -149 12885 -89
rect 5982 -287 6016 -227
rect 6142 -287 6176 -227
rect 12691 -287 12725 -227
rect 12851 -287 12885 -227
rect 5982 -425 6016 -365
rect 6142 -425 6176 -365
rect 12691 -425 12725 -365
rect 12851 -425 12885 -365
rect 5982 -563 6016 -503
rect 6142 -563 6176 -503
rect 12691 -563 12725 -503
rect 12851 -563 12885 -503
rect 5982 -701 6016 -641
rect 6142 -701 6176 -641
rect 12691 -701 12725 -641
rect 12851 -701 12885 -641
rect 244 -886 278 -826
rect 332 -886 366 -826
rect 5982 -839 6016 -779
rect 6142 -839 6176 -779
rect 6953 -886 6987 -826
rect 7041 -886 7075 -826
rect 12691 -839 12725 -779
rect 12851 -839 12885 -779
rect 52 -1024 86 -964
rect 148 -1024 182 -964
rect 244 -1024 278 -964
rect 332 -1024 366 -964
rect 896 -1023 930 -963
rect 985 -1023 1019 -963
rect 1630 -1023 1664 -963
rect 1732 -1023 1766 -963
rect 1840 -1023 1874 -963
rect 2968 -1023 3002 -963
rect 3072 -1023 3106 -963
rect 3178 -1023 3212 -963
rect 4180 -1023 4214 -963
rect 4283 -1023 4317 -963
rect 4390 -1023 4424 -963
rect 5032 -1023 5066 -963
rect 5122 -1023 5156 -963
rect 6761 -1024 6795 -964
rect 6857 -1024 6891 -964
rect 6953 -1024 6987 -964
rect 7041 -1024 7075 -964
rect 7605 -1023 7639 -963
rect 7694 -1023 7728 -963
rect 8339 -1023 8373 -963
rect 8441 -1023 8475 -963
rect 8549 -1023 8583 -963
rect 9677 -1023 9711 -963
rect 9781 -1023 9815 -963
rect 9887 -1023 9921 -963
rect 10889 -1023 10923 -963
rect 10992 -1023 11026 -963
rect 11099 -1023 11133 -963
rect 11741 -1023 11775 -963
rect 11831 -1023 11865 -963
rect 6309 -1331 6343 -1297
rect 6309 -1399 6343 -1365
rect 6393 -1331 6427 -1297
rect 6393 -1399 6427 -1365
rect 6499 -1331 6533 -1297
rect 6499 -1399 6533 -1365
rect 6583 -1331 6617 -1297
rect 6583 -1399 6617 -1365
rect 13018 -1331 13052 -1297
rect 13018 -1399 13052 -1365
rect 13102 -1331 13136 -1297
rect 13102 -1399 13136 -1365
rect 13208 -1331 13242 -1297
rect 13208 -1399 13242 -1365
rect 13292 -1331 13326 -1297
rect 13292 -1399 13326 -1365
<< pdiffc >>
rect 604 3627 638 3687
rect 692 3627 726 3687
rect 7313 3627 7347 3687
rect 7401 3627 7435 3687
rect 604 3489 638 3549
rect 692 3489 726 3549
rect 7313 3489 7347 3549
rect 7401 3489 7435 3549
rect 604 3351 638 3411
rect 692 3351 726 3411
rect 7313 3351 7347 3411
rect 7401 3351 7435 3411
rect 604 3213 638 3273
rect 692 3213 726 3273
rect 7313 3213 7347 3273
rect 7401 3213 7435 3273
rect 604 3075 638 3135
rect 692 3075 726 3135
rect 138 3006 172 3040
rect 138 2938 172 2972
rect 138 2870 172 2904
rect 222 3006 256 3040
rect 222 2938 256 2972
rect 222 2870 256 2904
rect 328 3006 362 3040
rect 328 2938 362 2972
rect 328 2870 362 2904
rect 412 3006 446 3040
rect 7313 3075 7347 3135
rect 7401 3075 7435 3135
rect 412 2938 446 2972
rect 604 2937 638 2997
rect 692 2937 726 2997
rect 6847 3006 6881 3040
rect 6847 2938 6881 2972
rect 412 2870 446 2904
rect 6847 2870 6881 2904
rect 6931 3006 6965 3040
rect 6931 2938 6965 2972
rect 6931 2870 6965 2904
rect 7037 3006 7071 3040
rect 7037 2938 7071 2972
rect 7037 2870 7071 2904
rect 7121 3006 7155 3040
rect 7121 2938 7155 2972
rect 7313 2937 7347 2997
rect 7401 2937 7435 2997
rect 7121 2870 7155 2904
rect 6389 2626 6423 2686
rect 6477 2626 6511 2686
rect 13098 2626 13132 2686
rect 13186 2626 13220 2686
rect 1246 2482 1280 2542
rect 1334 2485 1368 2545
rect 1978 2485 2012 2545
rect 2083 2485 2117 2545
rect 2192 2485 2226 2545
rect 3190 2485 3224 2545
rect 3294 2485 3328 2545
rect 3404 2485 3438 2545
rect 4402 2485 4436 2545
rect 4507 2485 4541 2545
rect 4616 2485 4650 2545
rect 5614 2485 5648 2545
rect 5721 2485 5755 2545
rect 5828 2485 5862 2545
rect 6389 2488 6423 2548
rect 6477 2488 6511 2548
rect 6573 2488 6607 2548
rect 6669 2488 6703 2548
rect 7955 2482 7989 2542
rect 8043 2485 8077 2545
rect 8687 2485 8721 2545
rect 8792 2485 8826 2545
rect 8901 2485 8935 2545
rect 9899 2485 9933 2545
rect 10003 2485 10037 2545
rect 10113 2485 10147 2545
rect 11111 2485 11145 2545
rect 11216 2485 11250 2545
rect 11325 2485 11359 2545
rect 12323 2485 12357 2545
rect 12430 2485 12464 2545
rect 12537 2485 12571 2545
rect 13098 2488 13132 2548
rect 13186 2488 13220 2548
rect 13282 2488 13316 2548
rect 13378 2488 13412 2548
rect 52 -1227 86 -1167
rect 148 -1227 182 -1167
rect 244 -1227 278 -1167
rect 332 -1227 366 -1167
rect 893 -1224 927 -1164
rect 1000 -1224 1034 -1164
rect 1107 -1224 1141 -1164
rect 2105 -1224 2139 -1164
rect 2214 -1224 2248 -1164
rect 2319 -1224 2353 -1164
rect 3317 -1224 3351 -1164
rect 3427 -1224 3461 -1164
rect 3531 -1224 3565 -1164
rect 4529 -1224 4563 -1164
rect 4638 -1224 4672 -1164
rect 4743 -1224 4777 -1164
rect 5387 -1224 5421 -1164
rect 5475 -1221 5509 -1161
rect 6761 -1227 6795 -1167
rect 6857 -1227 6891 -1167
rect 6953 -1227 6987 -1167
rect 7041 -1227 7075 -1167
rect 7602 -1224 7636 -1164
rect 7709 -1224 7743 -1164
rect 7816 -1224 7850 -1164
rect 8814 -1224 8848 -1164
rect 8923 -1224 8957 -1164
rect 9028 -1224 9062 -1164
rect 10026 -1224 10060 -1164
rect 10136 -1224 10170 -1164
rect 10240 -1224 10274 -1164
rect 11238 -1224 11272 -1164
rect 11347 -1224 11381 -1164
rect 11452 -1224 11486 -1164
rect 12096 -1224 12130 -1164
rect 12184 -1221 12218 -1161
rect 244 -1365 278 -1305
rect 332 -1365 366 -1305
rect 6953 -1365 6987 -1305
rect 7041 -1365 7075 -1305
rect 6309 -1583 6343 -1549
rect 6029 -1676 6063 -1616
rect 6117 -1676 6151 -1616
rect 6309 -1651 6343 -1617
rect 6309 -1719 6343 -1685
rect 6393 -1583 6427 -1549
rect 6393 -1651 6427 -1617
rect 6393 -1719 6427 -1685
rect 6499 -1583 6533 -1549
rect 6499 -1651 6533 -1617
rect 6499 -1719 6533 -1685
rect 6583 -1583 6617 -1549
rect 13018 -1583 13052 -1549
rect 6583 -1651 6617 -1617
rect 6583 -1719 6617 -1685
rect 12738 -1676 12772 -1616
rect 12826 -1676 12860 -1616
rect 13018 -1651 13052 -1617
rect 6029 -1814 6063 -1754
rect 6117 -1814 6151 -1754
rect 13018 -1719 13052 -1685
rect 13102 -1583 13136 -1549
rect 13102 -1651 13136 -1617
rect 13102 -1719 13136 -1685
rect 13208 -1583 13242 -1549
rect 13208 -1651 13242 -1617
rect 13208 -1719 13242 -1685
rect 13292 -1583 13326 -1549
rect 13292 -1651 13326 -1617
rect 13292 -1719 13326 -1685
rect 12738 -1814 12772 -1754
rect 12826 -1814 12860 -1754
rect 6029 -1952 6063 -1892
rect 6117 -1952 6151 -1892
rect 12738 -1952 12772 -1892
rect 12826 -1952 12860 -1892
rect 6029 -2090 6063 -2030
rect 6117 -2090 6151 -2030
rect 12738 -2090 12772 -2030
rect 12826 -2090 12860 -2030
rect 6029 -2228 6063 -2168
rect 6117 -2228 6151 -2168
rect 12738 -2228 12772 -2168
rect 12826 -2228 12860 -2168
rect 6029 -2366 6063 -2306
rect 6117 -2366 6151 -2306
rect 12738 -2366 12772 -2306
rect 12826 -2366 12860 -2306
<< psubdiff >>
rect 132 2509 156 2543
rect 190 2509 274 2543
rect 308 2509 418 2543
rect 452 2509 494 2543
rect 132 2507 494 2509
rect 6841 2509 6865 2543
rect 6899 2509 6983 2543
rect 7017 2509 7127 2543
rect 7161 2509 7203 2543
rect 6841 2507 7203 2509
rect 76 1702 194 1722
rect 76 1645 103 1702
rect 169 1645 194 1702
rect 76 1623 194 1645
rect 856 1318 960 1353
rect 856 1284 887 1318
rect 921 1284 960 1318
rect 856 1255 960 1284
rect 7565 1318 7669 1353
rect 7565 1284 7596 1318
rect 7630 1284 7669 1318
rect 7565 1255 7669 1284
rect 1254 1147 1586 1163
rect 1254 1113 1280 1147
rect 1314 1113 1360 1147
rect 1394 1113 1440 1147
rect 1474 1113 1520 1147
rect 1554 1113 1586 1147
rect 1254 1095 1586 1113
rect 1986 1147 2318 1163
rect 1986 1113 2012 1147
rect 2046 1113 2092 1147
rect 2126 1113 2172 1147
rect 2206 1113 2252 1147
rect 2286 1113 2318 1147
rect 1986 1095 2318 1113
rect 2588 1147 2920 1163
rect 2588 1113 2620 1147
rect 2654 1113 2700 1147
rect 2734 1113 2780 1147
rect 2814 1113 2860 1147
rect 2894 1113 2920 1147
rect 2588 1095 2920 1113
rect 3198 1147 3530 1163
rect 3198 1113 3224 1147
rect 3258 1113 3304 1147
rect 3338 1113 3384 1147
rect 3418 1113 3464 1147
rect 3498 1113 3530 1147
rect 3198 1095 3530 1113
rect 3800 1147 4132 1163
rect 3800 1113 3832 1147
rect 3866 1113 3912 1147
rect 3946 1113 3992 1147
rect 4026 1113 4072 1147
rect 4106 1113 4132 1147
rect 3800 1095 4132 1113
rect 4536 1147 4868 1163
rect 4536 1113 4562 1147
rect 4596 1113 4642 1147
rect 4676 1113 4722 1147
rect 4756 1113 4802 1147
rect 4836 1113 4868 1147
rect 4536 1095 4868 1113
rect 5138 1147 5470 1163
rect 5138 1113 5170 1147
rect 5204 1113 5250 1147
rect 5284 1113 5330 1147
rect 5364 1113 5410 1147
rect 5444 1113 5470 1147
rect 5138 1095 5470 1113
rect 5872 1147 6204 1163
rect 5872 1113 5904 1147
rect 5938 1113 5984 1147
rect 6018 1113 6064 1147
rect 6098 1113 6144 1147
rect 6178 1113 6204 1147
rect 7963 1147 8295 1163
rect 5872 1095 6204 1113
rect 7963 1113 7989 1147
rect 8023 1113 8069 1147
rect 8103 1113 8149 1147
rect 8183 1113 8229 1147
rect 8263 1113 8295 1147
rect 7963 1095 8295 1113
rect 8695 1147 9027 1163
rect 8695 1113 8721 1147
rect 8755 1113 8801 1147
rect 8835 1113 8881 1147
rect 8915 1113 8961 1147
rect 8995 1113 9027 1147
rect 8695 1095 9027 1113
rect 9297 1147 9629 1163
rect 9297 1113 9329 1147
rect 9363 1113 9409 1147
rect 9443 1113 9489 1147
rect 9523 1113 9569 1147
rect 9603 1113 9629 1147
rect 9297 1095 9629 1113
rect 9907 1147 10239 1163
rect 9907 1113 9933 1147
rect 9967 1113 10013 1147
rect 10047 1113 10093 1147
rect 10127 1113 10173 1147
rect 10207 1113 10239 1147
rect 9907 1095 10239 1113
rect 10509 1147 10841 1163
rect 10509 1113 10541 1147
rect 10575 1113 10621 1147
rect 10655 1113 10701 1147
rect 10735 1113 10781 1147
rect 10815 1113 10841 1147
rect 10509 1095 10841 1113
rect 11245 1147 11577 1163
rect 11245 1113 11271 1147
rect 11305 1113 11351 1147
rect 11385 1113 11431 1147
rect 11465 1113 11511 1147
rect 11545 1113 11577 1147
rect 11245 1095 11577 1113
rect 11847 1147 12179 1163
rect 11847 1113 11879 1147
rect 11913 1113 11959 1147
rect 11993 1113 12039 1147
rect 12073 1113 12119 1147
rect 12153 1113 12179 1147
rect 11847 1095 12179 1113
rect 12581 1147 12913 1163
rect 12581 1113 12613 1147
rect 12647 1113 12693 1147
rect 12727 1113 12773 1147
rect 12807 1113 12853 1147
rect 12887 1113 12913 1147
rect 12581 1095 12913 1113
rect 551 208 883 226
rect 551 174 577 208
rect 611 174 657 208
rect 691 174 737 208
rect 771 174 817 208
rect 851 174 883 208
rect 551 158 883 174
rect 1285 208 1617 226
rect 1285 174 1311 208
rect 1345 174 1391 208
rect 1425 174 1471 208
rect 1505 174 1551 208
rect 1585 174 1617 208
rect 1285 158 1617 174
rect 1887 208 2219 226
rect 1887 174 1919 208
rect 1953 174 1999 208
rect 2033 174 2079 208
rect 2113 174 2159 208
rect 2193 174 2219 208
rect 1887 158 2219 174
rect 2623 208 2955 226
rect 2623 174 2649 208
rect 2683 174 2729 208
rect 2763 174 2809 208
rect 2843 174 2889 208
rect 2923 174 2955 208
rect 2623 158 2955 174
rect 3225 208 3557 226
rect 3225 174 3257 208
rect 3291 174 3337 208
rect 3371 174 3417 208
rect 3451 174 3497 208
rect 3531 174 3557 208
rect 3225 158 3557 174
rect 3835 208 4167 226
rect 3835 174 3861 208
rect 3895 174 3941 208
rect 3975 174 4021 208
rect 4055 174 4101 208
rect 4135 174 4167 208
rect 3835 158 4167 174
rect 4437 208 4769 226
rect 4437 174 4469 208
rect 4503 174 4549 208
rect 4583 174 4629 208
rect 4663 174 4709 208
rect 4743 174 4769 208
rect 4437 158 4769 174
rect 5169 208 5501 226
rect 5169 174 5201 208
rect 5235 174 5281 208
rect 5315 174 5361 208
rect 5395 174 5441 208
rect 5475 174 5501 208
rect 7260 208 7592 226
rect 5169 158 5501 174
rect 7260 174 7286 208
rect 7320 174 7366 208
rect 7400 174 7446 208
rect 7480 174 7526 208
rect 7560 174 7592 208
rect 7260 158 7592 174
rect 7994 208 8326 226
rect 7994 174 8020 208
rect 8054 174 8100 208
rect 8134 174 8180 208
rect 8214 174 8260 208
rect 8294 174 8326 208
rect 7994 158 8326 174
rect 8596 208 8928 226
rect 8596 174 8628 208
rect 8662 174 8708 208
rect 8742 174 8788 208
rect 8822 174 8868 208
rect 8902 174 8928 208
rect 8596 158 8928 174
rect 9332 208 9664 226
rect 9332 174 9358 208
rect 9392 174 9438 208
rect 9472 174 9518 208
rect 9552 174 9598 208
rect 9632 174 9664 208
rect 9332 158 9664 174
rect 9934 208 10266 226
rect 9934 174 9966 208
rect 10000 174 10046 208
rect 10080 174 10126 208
rect 10160 174 10206 208
rect 10240 174 10266 208
rect 9934 158 10266 174
rect 10544 208 10876 226
rect 10544 174 10570 208
rect 10604 174 10650 208
rect 10684 174 10730 208
rect 10764 174 10810 208
rect 10844 174 10876 208
rect 10544 158 10876 174
rect 11146 208 11478 226
rect 11146 174 11178 208
rect 11212 174 11258 208
rect 11292 174 11338 208
rect 11372 174 11418 208
rect 11452 174 11478 208
rect 11146 158 11478 174
rect 11878 208 12210 226
rect 11878 174 11910 208
rect 11944 174 11990 208
rect 12024 174 12070 208
rect 12104 174 12150 208
rect 12184 174 12210 208
rect 11878 158 12210 174
rect 5795 37 5899 66
rect 5795 3 5834 37
rect 5868 3 5899 37
rect 5795 -32 5899 3
rect 12504 37 12608 66
rect 12504 3 12543 37
rect 12577 3 12608 37
rect 12504 -32 12608 3
rect 6261 -1188 6623 -1186
rect 6261 -1222 6303 -1188
rect 6337 -1222 6447 -1188
rect 6481 -1222 6565 -1188
rect 6599 -1222 6623 -1188
rect 12970 -1188 13332 -1186
rect 12970 -1222 13012 -1188
rect 13046 -1222 13156 -1188
rect 13190 -1222 13274 -1188
rect 13308 -1222 13332 -1188
<< nsubdiff >>
rect 802 3711 1340 3731
rect 802 3677 850 3711
rect 884 3677 930 3711
rect 964 3677 1010 3711
rect 1044 3677 1090 3711
rect 1124 3677 1170 3711
rect 1204 3677 1250 3711
rect 1284 3677 1340 3711
rect 802 3663 1340 3677
rect 1534 3714 2072 3734
rect 1534 3680 1582 3714
rect 1616 3680 1662 3714
rect 1696 3680 1742 3714
rect 1776 3680 1822 3714
rect 1856 3680 1902 3714
rect 1936 3680 1982 3714
rect 2016 3680 2072 3714
rect 1534 3666 2072 3680
rect 2132 3714 2670 3734
rect 2132 3680 2188 3714
rect 2222 3680 2268 3714
rect 2302 3680 2348 3714
rect 2382 3680 2428 3714
rect 2462 3680 2508 3714
rect 2542 3680 2588 3714
rect 2622 3680 2670 3714
rect 2132 3666 2670 3680
rect 2746 3714 3284 3734
rect 2746 3680 2794 3714
rect 2828 3680 2874 3714
rect 2908 3680 2954 3714
rect 2988 3680 3034 3714
rect 3068 3680 3114 3714
rect 3148 3680 3194 3714
rect 3228 3680 3284 3714
rect 2746 3666 3284 3680
rect 3344 3714 3882 3734
rect 3344 3680 3400 3714
rect 3434 3680 3480 3714
rect 3514 3680 3560 3714
rect 3594 3680 3640 3714
rect 3674 3680 3720 3714
rect 3754 3680 3800 3714
rect 3834 3680 3882 3714
rect 3344 3666 3882 3680
rect 3958 3714 4496 3734
rect 3958 3680 4006 3714
rect 4040 3680 4086 3714
rect 4120 3680 4166 3714
rect 4200 3680 4246 3714
rect 4280 3680 4326 3714
rect 4360 3680 4406 3714
rect 4440 3680 4496 3714
rect 3958 3666 4496 3680
rect 4556 3714 5094 3734
rect 4556 3680 4612 3714
rect 4646 3680 4692 3714
rect 4726 3680 4772 3714
rect 4806 3680 4852 3714
rect 4886 3680 4932 3714
rect 4966 3680 5012 3714
rect 5046 3680 5094 3714
rect 4556 3666 5094 3680
rect 5170 3714 5708 3734
rect 5170 3680 5218 3714
rect 5252 3680 5298 3714
rect 5332 3680 5378 3714
rect 5412 3680 5458 3714
rect 5492 3680 5538 3714
rect 5572 3680 5618 3714
rect 5652 3680 5708 3714
rect 5170 3666 5708 3680
rect 5768 3714 6306 3734
rect 5768 3680 5824 3714
rect 5858 3680 5904 3714
rect 5938 3680 5984 3714
rect 6018 3680 6064 3714
rect 6098 3680 6144 3714
rect 6178 3680 6224 3714
rect 6258 3680 6306 3714
rect 7511 3711 8049 3731
rect 5768 3666 6306 3680
rect 6538 3663 6624 3689
rect 6538 3629 6564 3663
rect 6598 3629 6624 3663
rect 6538 3603 6624 3629
rect 7015 3666 7101 3692
rect 7015 3632 7041 3666
rect 7075 3632 7101 3666
rect 7015 3606 7101 3632
rect 7511 3677 7559 3711
rect 7593 3677 7639 3711
rect 7673 3677 7719 3711
rect 7753 3677 7799 3711
rect 7833 3677 7879 3711
rect 7913 3677 7959 3711
rect 7993 3677 8049 3711
rect 7511 3663 8049 3677
rect 8243 3714 8781 3734
rect 8243 3680 8291 3714
rect 8325 3680 8371 3714
rect 8405 3680 8451 3714
rect 8485 3680 8531 3714
rect 8565 3680 8611 3714
rect 8645 3680 8691 3714
rect 8725 3680 8781 3714
rect 8243 3666 8781 3680
rect 8841 3714 9379 3734
rect 8841 3680 8897 3714
rect 8931 3680 8977 3714
rect 9011 3680 9057 3714
rect 9091 3680 9137 3714
rect 9171 3680 9217 3714
rect 9251 3680 9297 3714
rect 9331 3680 9379 3714
rect 8841 3666 9379 3680
rect 9455 3714 9993 3734
rect 9455 3680 9503 3714
rect 9537 3680 9583 3714
rect 9617 3680 9663 3714
rect 9697 3680 9743 3714
rect 9777 3680 9823 3714
rect 9857 3680 9903 3714
rect 9937 3680 9993 3714
rect 9455 3666 9993 3680
rect 10053 3714 10591 3734
rect 10053 3680 10109 3714
rect 10143 3680 10189 3714
rect 10223 3680 10269 3714
rect 10303 3680 10349 3714
rect 10383 3680 10429 3714
rect 10463 3680 10509 3714
rect 10543 3680 10591 3714
rect 10053 3666 10591 3680
rect 10667 3714 11205 3734
rect 10667 3680 10715 3714
rect 10749 3680 10795 3714
rect 10829 3680 10875 3714
rect 10909 3680 10955 3714
rect 10989 3680 11035 3714
rect 11069 3680 11115 3714
rect 11149 3680 11205 3714
rect 10667 3666 11205 3680
rect 11265 3714 11803 3734
rect 11265 3680 11321 3714
rect 11355 3680 11401 3714
rect 11435 3680 11481 3714
rect 11515 3680 11561 3714
rect 11595 3680 11641 3714
rect 11675 3680 11721 3714
rect 11755 3680 11803 3714
rect 11265 3666 11803 3680
rect 11879 3714 12417 3734
rect 11879 3680 11927 3714
rect 11961 3680 12007 3714
rect 12041 3680 12087 3714
rect 12121 3680 12167 3714
rect 12201 3680 12247 3714
rect 12281 3680 12327 3714
rect 12361 3680 12417 3714
rect 11879 3666 12417 3680
rect 12477 3714 13015 3734
rect 12477 3680 12533 3714
rect 12567 3680 12613 3714
rect 12647 3680 12693 3714
rect 12727 3680 12773 3714
rect 12807 3680 12853 3714
rect 12887 3680 12933 3714
rect 12967 3680 13015 3714
rect 12477 3666 13015 3680
rect 13247 3663 13333 3689
rect 13247 3629 13273 3663
rect 13307 3629 13333 3663
rect 13247 3603 13333 3629
rect 792 3533 875 3558
rect 792 3498 817 3533
rect 851 3498 875 3533
rect 792 3474 875 3498
rect 6543 3519 6629 3545
rect 6543 3485 6569 3519
rect 6603 3485 6629 3519
rect 6543 3459 6629 3485
rect 7004 3494 7090 3520
rect 7004 3460 7030 3494
rect 7064 3460 7090 3494
rect 7501 3533 7584 3558
rect 7501 3498 7526 3533
rect 7560 3498 7584 3533
rect 7004 3434 7090 3460
rect 7501 3474 7584 3498
rect 13252 3519 13338 3545
rect 13252 3485 13278 3519
rect 13312 3485 13338 3519
rect 13252 3459 13338 3485
rect 6544 3367 6630 3393
rect 6544 3333 6570 3367
rect 6604 3333 6630 3367
rect 13253 3367 13339 3393
rect 6544 3307 6630 3333
rect 7004 3302 7090 3328
rect 7004 3268 7030 3302
rect 7064 3268 7090 3302
rect 13253 3333 13279 3367
rect 13313 3333 13339 3367
rect 13253 3307 13339 3333
rect 7004 3242 7090 3268
rect 6544 3197 6630 3223
rect 6544 3163 6570 3197
rect 6604 3163 6630 3197
rect 106 3145 522 3147
rect 106 3111 136 3145
rect 170 3111 266 3145
rect 300 3111 412 3145
rect 446 3111 522 3145
rect 106 3107 522 3111
rect 6544 3137 6630 3163
rect 13253 3197 13339 3223
rect 13253 3163 13279 3197
rect 13313 3163 13339 3197
rect 6815 3145 7231 3147
rect 6815 3111 6845 3145
rect 6879 3111 6975 3145
rect 7009 3111 7121 3145
rect 7155 3111 7231 3145
rect 6815 3107 7231 3111
rect 6543 3040 6629 3066
rect 13253 3137 13339 3163
rect 6543 3006 6569 3040
rect 6603 3006 6629 3040
rect 6543 2980 6629 3006
rect 13252 3040 13338 3066
rect 13252 3006 13278 3040
rect 13312 3006 13338 3040
rect 13252 2980 13338 3006
rect 126 -1685 212 -1659
rect 126 -1719 152 -1685
rect 186 -1719 212 -1685
rect 126 -1745 212 -1719
rect 6835 -1685 6921 -1659
rect 6835 -1719 6861 -1685
rect 6895 -1719 6921 -1685
rect 125 -1842 211 -1816
rect 6835 -1745 6921 -1719
rect 6233 -1790 6649 -1786
rect 6233 -1824 6309 -1790
rect 6343 -1824 6455 -1790
rect 6489 -1824 6585 -1790
rect 6619 -1824 6649 -1790
rect 6233 -1826 6649 -1824
rect 125 -1876 151 -1842
rect 185 -1876 211 -1842
rect 125 -1902 211 -1876
rect 6834 -1842 6920 -1816
rect 12942 -1790 13358 -1786
rect 12942 -1824 13018 -1790
rect 13052 -1824 13164 -1790
rect 13198 -1824 13294 -1790
rect 13328 -1824 13358 -1790
rect 12942 -1826 13358 -1824
rect 6834 -1876 6860 -1842
rect 6894 -1876 6920 -1842
rect 6412 -1914 6498 -1888
rect 6834 -1902 6920 -1876
rect 6412 -1948 6438 -1914
rect 6472 -1948 6498 -1914
rect 125 -2012 211 -1986
rect 125 -2046 151 -2012
rect 185 -2046 211 -2012
rect 6412 -1974 6498 -1948
rect 6834 -2012 6920 -1986
rect 125 -2072 211 -2046
rect 6834 -2046 6860 -2012
rect 6894 -2046 6920 -2012
rect 6834 -2072 6920 -2046
rect 126 -2164 212 -2138
rect 126 -2198 152 -2164
rect 186 -2198 212 -2164
rect 126 -2224 212 -2198
rect 5880 -2177 5963 -2153
rect 6412 -2110 6498 -2084
rect 6412 -2144 6438 -2110
rect 6472 -2144 6498 -2110
rect 5880 -2212 5904 -2177
rect 5938 -2212 5963 -2177
rect 5880 -2237 5963 -2212
rect 6412 -2170 6498 -2144
rect 6835 -2164 6921 -2138
rect 6835 -2198 6861 -2164
rect 6895 -2198 6921 -2164
rect 6835 -2224 6921 -2198
rect 12589 -2177 12672 -2153
rect 12589 -2212 12613 -2177
rect 12647 -2212 12672 -2177
rect 12589 -2237 12672 -2212
rect 131 -2308 217 -2282
rect 6412 -2285 6498 -2259
rect 131 -2342 157 -2308
rect 191 -2342 217 -2308
rect 131 -2368 217 -2342
rect 449 -2359 987 -2345
rect 449 -2393 497 -2359
rect 531 -2393 577 -2359
rect 611 -2393 657 -2359
rect 691 -2393 737 -2359
rect 771 -2393 817 -2359
rect 851 -2393 897 -2359
rect 931 -2393 987 -2359
rect 449 -2413 987 -2393
rect 1047 -2359 1585 -2345
rect 1047 -2393 1103 -2359
rect 1137 -2393 1183 -2359
rect 1217 -2393 1263 -2359
rect 1297 -2393 1343 -2359
rect 1377 -2393 1423 -2359
rect 1457 -2393 1503 -2359
rect 1537 -2393 1585 -2359
rect 1047 -2413 1585 -2393
rect 1661 -2359 2199 -2345
rect 1661 -2393 1709 -2359
rect 1743 -2393 1789 -2359
rect 1823 -2393 1869 -2359
rect 1903 -2393 1949 -2359
rect 1983 -2393 2029 -2359
rect 2063 -2393 2109 -2359
rect 2143 -2393 2199 -2359
rect 1661 -2413 2199 -2393
rect 2259 -2359 2797 -2345
rect 2259 -2393 2315 -2359
rect 2349 -2393 2395 -2359
rect 2429 -2393 2475 -2359
rect 2509 -2393 2555 -2359
rect 2589 -2393 2635 -2359
rect 2669 -2393 2715 -2359
rect 2749 -2393 2797 -2359
rect 2259 -2413 2797 -2393
rect 2873 -2359 3411 -2345
rect 2873 -2393 2921 -2359
rect 2955 -2393 3001 -2359
rect 3035 -2393 3081 -2359
rect 3115 -2393 3161 -2359
rect 3195 -2393 3241 -2359
rect 3275 -2393 3321 -2359
rect 3355 -2393 3411 -2359
rect 2873 -2413 3411 -2393
rect 3471 -2359 4009 -2345
rect 3471 -2393 3527 -2359
rect 3561 -2393 3607 -2359
rect 3641 -2393 3687 -2359
rect 3721 -2393 3767 -2359
rect 3801 -2393 3847 -2359
rect 3881 -2393 3927 -2359
rect 3961 -2393 4009 -2359
rect 3471 -2413 4009 -2393
rect 4085 -2359 4623 -2345
rect 4085 -2393 4133 -2359
rect 4167 -2393 4213 -2359
rect 4247 -2393 4293 -2359
rect 4327 -2393 4373 -2359
rect 4407 -2393 4453 -2359
rect 4487 -2393 4533 -2359
rect 4567 -2393 4623 -2359
rect 4085 -2413 4623 -2393
rect 4683 -2359 5221 -2345
rect 4683 -2393 4739 -2359
rect 4773 -2393 4819 -2359
rect 4853 -2393 4899 -2359
rect 4933 -2393 4979 -2359
rect 5013 -2393 5059 -2359
rect 5093 -2393 5139 -2359
rect 5173 -2393 5221 -2359
rect 4683 -2413 5221 -2393
rect 5415 -2356 5953 -2342
rect 5415 -2390 5471 -2356
rect 5505 -2390 5551 -2356
rect 5585 -2390 5631 -2356
rect 5665 -2390 5711 -2356
rect 5745 -2390 5791 -2356
rect 5825 -2390 5871 -2356
rect 5905 -2390 5953 -2356
rect 6412 -2319 6438 -2285
rect 6472 -2319 6498 -2285
rect 6412 -2345 6498 -2319
rect 6840 -2308 6926 -2282
rect 6840 -2342 6866 -2308
rect 6900 -2342 6926 -2308
rect 6840 -2368 6926 -2342
rect 7158 -2359 7696 -2345
rect 5415 -2410 5953 -2390
rect 7158 -2393 7206 -2359
rect 7240 -2393 7286 -2359
rect 7320 -2393 7366 -2359
rect 7400 -2393 7446 -2359
rect 7480 -2393 7526 -2359
rect 7560 -2393 7606 -2359
rect 7640 -2393 7696 -2359
rect 7158 -2413 7696 -2393
rect 7756 -2359 8294 -2345
rect 7756 -2393 7812 -2359
rect 7846 -2393 7892 -2359
rect 7926 -2393 7972 -2359
rect 8006 -2393 8052 -2359
rect 8086 -2393 8132 -2359
rect 8166 -2393 8212 -2359
rect 8246 -2393 8294 -2359
rect 7756 -2413 8294 -2393
rect 8370 -2359 8908 -2345
rect 8370 -2393 8418 -2359
rect 8452 -2393 8498 -2359
rect 8532 -2393 8578 -2359
rect 8612 -2393 8658 -2359
rect 8692 -2393 8738 -2359
rect 8772 -2393 8818 -2359
rect 8852 -2393 8908 -2359
rect 8370 -2413 8908 -2393
rect 8968 -2359 9506 -2345
rect 8968 -2393 9024 -2359
rect 9058 -2393 9104 -2359
rect 9138 -2393 9184 -2359
rect 9218 -2393 9264 -2359
rect 9298 -2393 9344 -2359
rect 9378 -2393 9424 -2359
rect 9458 -2393 9506 -2359
rect 8968 -2413 9506 -2393
rect 9582 -2359 10120 -2345
rect 9582 -2393 9630 -2359
rect 9664 -2393 9710 -2359
rect 9744 -2393 9790 -2359
rect 9824 -2393 9870 -2359
rect 9904 -2393 9950 -2359
rect 9984 -2393 10030 -2359
rect 10064 -2393 10120 -2359
rect 9582 -2413 10120 -2393
rect 10180 -2359 10718 -2345
rect 10180 -2393 10236 -2359
rect 10270 -2393 10316 -2359
rect 10350 -2393 10396 -2359
rect 10430 -2393 10476 -2359
rect 10510 -2393 10556 -2359
rect 10590 -2393 10636 -2359
rect 10670 -2393 10718 -2359
rect 10180 -2413 10718 -2393
rect 10794 -2359 11332 -2345
rect 10794 -2393 10842 -2359
rect 10876 -2393 10922 -2359
rect 10956 -2393 11002 -2359
rect 11036 -2393 11082 -2359
rect 11116 -2393 11162 -2359
rect 11196 -2393 11242 -2359
rect 11276 -2393 11332 -2359
rect 10794 -2413 11332 -2393
rect 11392 -2359 11930 -2345
rect 11392 -2393 11448 -2359
rect 11482 -2393 11528 -2359
rect 11562 -2393 11608 -2359
rect 11642 -2393 11688 -2359
rect 11722 -2393 11768 -2359
rect 11802 -2393 11848 -2359
rect 11882 -2393 11930 -2359
rect 11392 -2413 11930 -2393
rect 12124 -2356 12662 -2342
rect 12124 -2390 12180 -2356
rect 12214 -2390 12260 -2356
rect 12294 -2390 12340 -2356
rect 12374 -2390 12420 -2356
rect 12454 -2390 12500 -2356
rect 12534 -2390 12580 -2356
rect 12614 -2390 12662 -2356
rect 12124 -2410 12662 -2390
<< psubdiffcont >>
rect 156 2509 190 2543
rect 274 2509 308 2543
rect 418 2509 452 2543
rect 6865 2509 6899 2543
rect 6983 2509 7017 2543
rect 7127 2509 7161 2543
rect 103 1645 169 1702
rect 887 1284 921 1318
rect 7596 1284 7630 1318
rect 1280 1113 1314 1147
rect 1360 1113 1394 1147
rect 1440 1113 1474 1147
rect 1520 1113 1554 1147
rect 2012 1113 2046 1147
rect 2092 1113 2126 1147
rect 2172 1113 2206 1147
rect 2252 1113 2286 1147
rect 2620 1113 2654 1147
rect 2700 1113 2734 1147
rect 2780 1113 2814 1147
rect 2860 1113 2894 1147
rect 3224 1113 3258 1147
rect 3304 1113 3338 1147
rect 3384 1113 3418 1147
rect 3464 1113 3498 1147
rect 3832 1113 3866 1147
rect 3912 1113 3946 1147
rect 3992 1113 4026 1147
rect 4072 1113 4106 1147
rect 4562 1113 4596 1147
rect 4642 1113 4676 1147
rect 4722 1113 4756 1147
rect 4802 1113 4836 1147
rect 5170 1113 5204 1147
rect 5250 1113 5284 1147
rect 5330 1113 5364 1147
rect 5410 1113 5444 1147
rect 5904 1113 5938 1147
rect 5984 1113 6018 1147
rect 6064 1113 6098 1147
rect 6144 1113 6178 1147
rect 7989 1113 8023 1147
rect 8069 1113 8103 1147
rect 8149 1113 8183 1147
rect 8229 1113 8263 1147
rect 8721 1113 8755 1147
rect 8801 1113 8835 1147
rect 8881 1113 8915 1147
rect 8961 1113 8995 1147
rect 9329 1113 9363 1147
rect 9409 1113 9443 1147
rect 9489 1113 9523 1147
rect 9569 1113 9603 1147
rect 9933 1113 9967 1147
rect 10013 1113 10047 1147
rect 10093 1113 10127 1147
rect 10173 1113 10207 1147
rect 10541 1113 10575 1147
rect 10621 1113 10655 1147
rect 10701 1113 10735 1147
rect 10781 1113 10815 1147
rect 11271 1113 11305 1147
rect 11351 1113 11385 1147
rect 11431 1113 11465 1147
rect 11511 1113 11545 1147
rect 11879 1113 11913 1147
rect 11959 1113 11993 1147
rect 12039 1113 12073 1147
rect 12119 1113 12153 1147
rect 12613 1113 12647 1147
rect 12693 1113 12727 1147
rect 12773 1113 12807 1147
rect 12853 1113 12887 1147
rect 577 174 611 208
rect 657 174 691 208
rect 737 174 771 208
rect 817 174 851 208
rect 1311 174 1345 208
rect 1391 174 1425 208
rect 1471 174 1505 208
rect 1551 174 1585 208
rect 1919 174 1953 208
rect 1999 174 2033 208
rect 2079 174 2113 208
rect 2159 174 2193 208
rect 2649 174 2683 208
rect 2729 174 2763 208
rect 2809 174 2843 208
rect 2889 174 2923 208
rect 3257 174 3291 208
rect 3337 174 3371 208
rect 3417 174 3451 208
rect 3497 174 3531 208
rect 3861 174 3895 208
rect 3941 174 3975 208
rect 4021 174 4055 208
rect 4101 174 4135 208
rect 4469 174 4503 208
rect 4549 174 4583 208
rect 4629 174 4663 208
rect 4709 174 4743 208
rect 5201 174 5235 208
rect 5281 174 5315 208
rect 5361 174 5395 208
rect 5441 174 5475 208
rect 7286 174 7320 208
rect 7366 174 7400 208
rect 7446 174 7480 208
rect 7526 174 7560 208
rect 8020 174 8054 208
rect 8100 174 8134 208
rect 8180 174 8214 208
rect 8260 174 8294 208
rect 8628 174 8662 208
rect 8708 174 8742 208
rect 8788 174 8822 208
rect 8868 174 8902 208
rect 9358 174 9392 208
rect 9438 174 9472 208
rect 9518 174 9552 208
rect 9598 174 9632 208
rect 9966 174 10000 208
rect 10046 174 10080 208
rect 10126 174 10160 208
rect 10206 174 10240 208
rect 10570 174 10604 208
rect 10650 174 10684 208
rect 10730 174 10764 208
rect 10810 174 10844 208
rect 11178 174 11212 208
rect 11258 174 11292 208
rect 11338 174 11372 208
rect 11418 174 11452 208
rect 11910 174 11944 208
rect 11990 174 12024 208
rect 12070 174 12104 208
rect 12150 174 12184 208
rect 5834 3 5868 37
rect 12543 3 12577 37
rect 6303 -1222 6337 -1188
rect 6447 -1222 6481 -1188
rect 6565 -1222 6599 -1188
rect 13012 -1222 13046 -1188
rect 13156 -1222 13190 -1188
rect 13274 -1222 13308 -1188
<< nsubdiffcont >>
rect 850 3677 884 3711
rect 930 3677 964 3711
rect 1010 3677 1044 3711
rect 1090 3677 1124 3711
rect 1170 3677 1204 3711
rect 1250 3677 1284 3711
rect 1582 3680 1616 3714
rect 1662 3680 1696 3714
rect 1742 3680 1776 3714
rect 1822 3680 1856 3714
rect 1902 3680 1936 3714
rect 1982 3680 2016 3714
rect 2188 3680 2222 3714
rect 2268 3680 2302 3714
rect 2348 3680 2382 3714
rect 2428 3680 2462 3714
rect 2508 3680 2542 3714
rect 2588 3680 2622 3714
rect 2794 3680 2828 3714
rect 2874 3680 2908 3714
rect 2954 3680 2988 3714
rect 3034 3680 3068 3714
rect 3114 3680 3148 3714
rect 3194 3680 3228 3714
rect 3400 3680 3434 3714
rect 3480 3680 3514 3714
rect 3560 3680 3594 3714
rect 3640 3680 3674 3714
rect 3720 3680 3754 3714
rect 3800 3680 3834 3714
rect 4006 3680 4040 3714
rect 4086 3680 4120 3714
rect 4166 3680 4200 3714
rect 4246 3680 4280 3714
rect 4326 3680 4360 3714
rect 4406 3680 4440 3714
rect 4612 3680 4646 3714
rect 4692 3680 4726 3714
rect 4772 3680 4806 3714
rect 4852 3680 4886 3714
rect 4932 3680 4966 3714
rect 5012 3680 5046 3714
rect 5218 3680 5252 3714
rect 5298 3680 5332 3714
rect 5378 3680 5412 3714
rect 5458 3680 5492 3714
rect 5538 3680 5572 3714
rect 5618 3680 5652 3714
rect 5824 3680 5858 3714
rect 5904 3680 5938 3714
rect 5984 3680 6018 3714
rect 6064 3680 6098 3714
rect 6144 3680 6178 3714
rect 6224 3680 6258 3714
rect 6564 3629 6598 3663
rect 7041 3632 7075 3666
rect 7559 3677 7593 3711
rect 7639 3677 7673 3711
rect 7719 3677 7753 3711
rect 7799 3677 7833 3711
rect 7879 3677 7913 3711
rect 7959 3677 7993 3711
rect 8291 3680 8325 3714
rect 8371 3680 8405 3714
rect 8451 3680 8485 3714
rect 8531 3680 8565 3714
rect 8611 3680 8645 3714
rect 8691 3680 8725 3714
rect 8897 3680 8931 3714
rect 8977 3680 9011 3714
rect 9057 3680 9091 3714
rect 9137 3680 9171 3714
rect 9217 3680 9251 3714
rect 9297 3680 9331 3714
rect 9503 3680 9537 3714
rect 9583 3680 9617 3714
rect 9663 3680 9697 3714
rect 9743 3680 9777 3714
rect 9823 3680 9857 3714
rect 9903 3680 9937 3714
rect 10109 3680 10143 3714
rect 10189 3680 10223 3714
rect 10269 3680 10303 3714
rect 10349 3680 10383 3714
rect 10429 3680 10463 3714
rect 10509 3680 10543 3714
rect 10715 3680 10749 3714
rect 10795 3680 10829 3714
rect 10875 3680 10909 3714
rect 10955 3680 10989 3714
rect 11035 3680 11069 3714
rect 11115 3680 11149 3714
rect 11321 3680 11355 3714
rect 11401 3680 11435 3714
rect 11481 3680 11515 3714
rect 11561 3680 11595 3714
rect 11641 3680 11675 3714
rect 11721 3680 11755 3714
rect 11927 3680 11961 3714
rect 12007 3680 12041 3714
rect 12087 3680 12121 3714
rect 12167 3680 12201 3714
rect 12247 3680 12281 3714
rect 12327 3680 12361 3714
rect 12533 3680 12567 3714
rect 12613 3680 12647 3714
rect 12693 3680 12727 3714
rect 12773 3680 12807 3714
rect 12853 3680 12887 3714
rect 12933 3680 12967 3714
rect 13273 3629 13307 3663
rect 817 3498 851 3533
rect 6569 3485 6603 3519
rect 7030 3460 7064 3494
rect 7526 3498 7560 3533
rect 13278 3485 13312 3519
rect 6570 3333 6604 3367
rect 7030 3268 7064 3302
rect 13279 3333 13313 3367
rect 6570 3163 6604 3197
rect 136 3111 170 3145
rect 266 3111 300 3145
rect 412 3111 446 3145
rect 13279 3163 13313 3197
rect 6845 3111 6879 3145
rect 6975 3111 7009 3145
rect 7121 3111 7155 3145
rect 6569 3006 6603 3040
rect 13278 3006 13312 3040
rect 152 -1719 186 -1685
rect 6861 -1719 6895 -1685
rect 6309 -1824 6343 -1790
rect 6455 -1824 6489 -1790
rect 6585 -1824 6619 -1790
rect 151 -1876 185 -1842
rect 13018 -1824 13052 -1790
rect 13164 -1824 13198 -1790
rect 13294 -1824 13328 -1790
rect 6860 -1876 6894 -1842
rect 6438 -1948 6472 -1914
rect 151 -2046 185 -2012
rect 6860 -2046 6894 -2012
rect 152 -2198 186 -2164
rect 6438 -2144 6472 -2110
rect 5904 -2212 5938 -2177
rect 6861 -2198 6895 -2164
rect 12613 -2212 12647 -2177
rect 157 -2342 191 -2308
rect 497 -2393 531 -2359
rect 577 -2393 611 -2359
rect 657 -2393 691 -2359
rect 737 -2393 771 -2359
rect 817 -2393 851 -2359
rect 897 -2393 931 -2359
rect 1103 -2393 1137 -2359
rect 1183 -2393 1217 -2359
rect 1263 -2393 1297 -2359
rect 1343 -2393 1377 -2359
rect 1423 -2393 1457 -2359
rect 1503 -2393 1537 -2359
rect 1709 -2393 1743 -2359
rect 1789 -2393 1823 -2359
rect 1869 -2393 1903 -2359
rect 1949 -2393 1983 -2359
rect 2029 -2393 2063 -2359
rect 2109 -2393 2143 -2359
rect 2315 -2393 2349 -2359
rect 2395 -2393 2429 -2359
rect 2475 -2393 2509 -2359
rect 2555 -2393 2589 -2359
rect 2635 -2393 2669 -2359
rect 2715 -2393 2749 -2359
rect 2921 -2393 2955 -2359
rect 3001 -2393 3035 -2359
rect 3081 -2393 3115 -2359
rect 3161 -2393 3195 -2359
rect 3241 -2393 3275 -2359
rect 3321 -2393 3355 -2359
rect 3527 -2393 3561 -2359
rect 3607 -2393 3641 -2359
rect 3687 -2393 3721 -2359
rect 3767 -2393 3801 -2359
rect 3847 -2393 3881 -2359
rect 3927 -2393 3961 -2359
rect 4133 -2393 4167 -2359
rect 4213 -2393 4247 -2359
rect 4293 -2393 4327 -2359
rect 4373 -2393 4407 -2359
rect 4453 -2393 4487 -2359
rect 4533 -2393 4567 -2359
rect 4739 -2393 4773 -2359
rect 4819 -2393 4853 -2359
rect 4899 -2393 4933 -2359
rect 4979 -2393 5013 -2359
rect 5059 -2393 5093 -2359
rect 5139 -2393 5173 -2359
rect 5471 -2390 5505 -2356
rect 5551 -2390 5585 -2356
rect 5631 -2390 5665 -2356
rect 5711 -2390 5745 -2356
rect 5791 -2390 5825 -2356
rect 5871 -2390 5905 -2356
rect 6438 -2319 6472 -2285
rect 6866 -2342 6900 -2308
rect 7206 -2393 7240 -2359
rect 7286 -2393 7320 -2359
rect 7366 -2393 7400 -2359
rect 7446 -2393 7480 -2359
rect 7526 -2393 7560 -2359
rect 7606 -2393 7640 -2359
rect 7812 -2393 7846 -2359
rect 7892 -2393 7926 -2359
rect 7972 -2393 8006 -2359
rect 8052 -2393 8086 -2359
rect 8132 -2393 8166 -2359
rect 8212 -2393 8246 -2359
rect 8418 -2393 8452 -2359
rect 8498 -2393 8532 -2359
rect 8578 -2393 8612 -2359
rect 8658 -2393 8692 -2359
rect 8738 -2393 8772 -2359
rect 8818 -2393 8852 -2359
rect 9024 -2393 9058 -2359
rect 9104 -2393 9138 -2359
rect 9184 -2393 9218 -2359
rect 9264 -2393 9298 -2359
rect 9344 -2393 9378 -2359
rect 9424 -2393 9458 -2359
rect 9630 -2393 9664 -2359
rect 9710 -2393 9744 -2359
rect 9790 -2393 9824 -2359
rect 9870 -2393 9904 -2359
rect 9950 -2393 9984 -2359
rect 10030 -2393 10064 -2359
rect 10236 -2393 10270 -2359
rect 10316 -2393 10350 -2359
rect 10396 -2393 10430 -2359
rect 10476 -2393 10510 -2359
rect 10556 -2393 10590 -2359
rect 10636 -2393 10670 -2359
rect 10842 -2393 10876 -2359
rect 10922 -2393 10956 -2359
rect 11002 -2393 11036 -2359
rect 11082 -2393 11116 -2359
rect 11162 -2393 11196 -2359
rect 11242 -2393 11276 -2359
rect 11448 -2393 11482 -2359
rect 11528 -2393 11562 -2359
rect 11608 -2393 11642 -2359
rect 11688 -2393 11722 -2359
rect 11768 -2393 11802 -2359
rect 11848 -2393 11882 -2359
rect 12180 -2390 12214 -2356
rect 12260 -2390 12294 -2356
rect 12340 -2390 12374 -2356
rect 12420 -2390 12454 -2356
rect 12500 -2390 12534 -2356
rect 12580 -2390 12614 -2356
<< poly >>
rect 650 3699 680 3729
rect 7359 3699 7389 3729
rect 650 3561 680 3615
rect 7359 3561 7389 3615
rect 650 3423 680 3477
rect 7359 3423 7389 3477
rect 650 3285 680 3339
rect 7359 3285 7389 3339
rect 650 3147 680 3201
rect 182 3052 212 3078
rect 372 3052 402 3078
rect 7359 3147 7389 3201
rect 650 3009 680 3063
rect 6891 3052 6921 3078
rect 7081 3052 7111 3078
rect 650 2894 680 2925
rect 632 2878 698 2894
rect 182 2820 212 2852
rect 126 2804 212 2820
rect 126 2770 142 2804
rect 176 2770 212 2804
rect 126 2754 212 2770
rect 182 2732 212 2754
rect 372 2820 402 2852
rect 632 2844 648 2878
rect 682 2844 698 2878
rect 7359 3009 7389 3063
rect 7359 2894 7389 2925
rect 7341 2878 7407 2894
rect 632 2828 698 2844
rect 6891 2820 6921 2852
rect 372 2804 458 2820
rect 372 2770 408 2804
rect 442 2770 458 2804
rect 372 2754 458 2770
rect 6835 2804 6921 2820
rect 6835 2770 6851 2804
rect 6885 2770 6921 2804
rect 6835 2754 6921 2770
rect 372 2732 402 2754
rect 6891 2732 6921 2754
rect 7081 2820 7111 2852
rect 7341 2844 7357 2878
rect 7391 2844 7407 2878
rect 7341 2828 7407 2844
rect 7081 2804 7167 2820
rect 7081 2770 7117 2804
rect 7151 2770 7167 2804
rect 7081 2754 7167 2770
rect 7081 2732 7111 2754
rect 6435 2698 6465 2729
rect 1274 2635 1340 2651
rect 182 2576 212 2602
rect 372 2576 402 2602
rect 1274 2601 1290 2635
rect 1324 2601 1340 2635
rect 1274 2585 1340 2601
rect 2006 2638 2072 2654
rect 2006 2604 2022 2638
rect 2056 2604 2072 2638
rect 2006 2588 2072 2604
rect 2132 2638 2198 2654
rect 2132 2604 2148 2638
rect 2182 2604 2198 2638
rect 2132 2588 2198 2604
rect 3218 2638 3284 2654
rect 3218 2604 3234 2638
rect 3268 2604 3284 2638
rect 3218 2588 3284 2604
rect 3344 2638 3410 2654
rect 3344 2604 3360 2638
rect 3394 2604 3410 2638
rect 3344 2588 3410 2604
rect 4430 2638 4496 2654
rect 4430 2604 4446 2638
rect 4480 2604 4496 2638
rect 4430 2588 4496 2604
rect 4556 2638 4622 2654
rect 4556 2604 4572 2638
rect 4606 2604 4622 2638
rect 4556 2588 4622 2604
rect 5642 2638 5708 2654
rect 5642 2604 5658 2638
rect 5692 2604 5708 2638
rect 5642 2588 5708 2604
rect 5768 2638 5834 2654
rect 5768 2604 5784 2638
rect 5818 2604 5834 2638
rect 5768 2588 5834 2604
rect 1292 2554 1322 2585
rect 2024 2557 2054 2588
rect 2150 2557 2180 2588
rect 3236 2557 3266 2588
rect 3362 2557 3392 2588
rect 4448 2557 4478 2588
rect 4574 2557 4604 2588
rect 5660 2557 5690 2588
rect 5786 2557 5816 2588
rect 6435 2560 6465 2614
rect 13144 2698 13174 2729
rect 7983 2635 8049 2651
rect 6527 2560 6557 2586
rect 6623 2560 6653 2591
rect 6891 2576 6921 2602
rect 7081 2576 7111 2602
rect 7983 2601 7999 2635
rect 8033 2601 8049 2635
rect 7983 2585 8049 2601
rect 8715 2638 8781 2654
rect 8715 2604 8731 2638
rect 8765 2604 8781 2638
rect 8715 2588 8781 2604
rect 8841 2638 8907 2654
rect 8841 2604 8857 2638
rect 8891 2604 8907 2638
rect 8841 2588 8907 2604
rect 9927 2638 9993 2654
rect 9927 2604 9943 2638
rect 9977 2604 9993 2638
rect 9927 2588 9993 2604
rect 10053 2638 10119 2654
rect 10053 2604 10069 2638
rect 10103 2604 10119 2638
rect 10053 2588 10119 2604
rect 11139 2638 11205 2654
rect 11139 2604 11155 2638
rect 11189 2604 11205 2638
rect 11139 2588 11205 2604
rect 11265 2638 11331 2654
rect 11265 2604 11281 2638
rect 11315 2604 11331 2638
rect 11265 2588 11331 2604
rect 12351 2638 12417 2654
rect 12351 2604 12367 2638
rect 12401 2604 12417 2638
rect 12351 2588 12417 2604
rect 12477 2638 12543 2654
rect 12477 2604 12493 2638
rect 12527 2604 12543 2638
rect 12477 2588 12543 2604
rect 8001 2554 8031 2585
rect 8733 2557 8763 2588
rect 8859 2557 8889 2588
rect 9945 2557 9975 2588
rect 10071 2557 10101 2588
rect 11157 2557 11187 2588
rect 11283 2557 11313 2588
rect 12369 2557 12399 2588
rect 12495 2557 12525 2588
rect 13144 2560 13174 2614
rect 13236 2560 13266 2586
rect 13332 2560 13362 2591
rect 1292 2442 1322 2470
rect 2024 2445 2054 2473
rect 2150 2445 2180 2473
rect 3236 2445 3266 2473
rect 3362 2445 3392 2473
rect 4448 2445 4478 2473
rect 4574 2445 4604 2473
rect 5660 2445 5690 2473
rect 5786 2445 5816 2473
rect 6435 2451 6465 2476
rect 6306 2431 6465 2451
rect 6527 2451 6557 2476
rect 6623 2451 6653 2476
rect 6527 2445 6653 2451
rect 6306 2397 6318 2431
rect 6352 2397 6465 2431
rect 1645 2356 1675 2382
rect 2377 2356 2407 2382
rect 2499 2356 2529 2382
rect 3589 2356 3619 2382
rect 3711 2356 3741 2382
rect 4927 2356 4957 2382
rect 5049 2356 5079 2382
rect 5783 2356 5813 2382
rect 6306 2378 6465 2397
rect 6509 2429 6653 2445
rect 8001 2442 8031 2470
rect 8733 2445 8763 2473
rect 8859 2445 8889 2473
rect 9945 2445 9975 2473
rect 10071 2445 10101 2473
rect 11157 2445 11187 2473
rect 11283 2445 11313 2473
rect 12369 2445 12399 2473
rect 12495 2445 12525 2473
rect 13144 2451 13174 2476
rect 6509 2395 6525 2429
rect 6559 2395 6653 2429
rect 6509 2379 6653 2395
rect 13015 2431 13174 2451
rect 13236 2451 13266 2476
rect 13332 2451 13362 2476
rect 13236 2445 13362 2451
rect 13015 2397 13027 2431
rect 13061 2397 13174 2431
rect 6435 2357 6465 2378
rect 6527 2372 6653 2379
rect 6527 2357 6557 2372
rect 6623 2357 6653 2372
rect 8354 2356 8384 2382
rect 9086 2356 9116 2382
rect 9208 2356 9238 2382
rect 10298 2356 10328 2382
rect 10420 2356 10450 2382
rect 11636 2356 11666 2382
rect 11758 2356 11788 2382
rect 12492 2356 12522 2382
rect 13015 2378 13174 2397
rect 13218 2429 13362 2445
rect 13218 2395 13234 2429
rect 13268 2395 13362 2429
rect 13218 2379 13362 2395
rect 13144 2357 13174 2378
rect 13236 2372 13362 2379
rect 13236 2357 13266 2372
rect 13332 2357 13362 2372
rect 643 2244 709 2260
rect 1645 2250 1675 2272
rect 2377 2250 2407 2272
rect 2499 2250 2529 2272
rect 3589 2250 3619 2272
rect 3711 2250 3741 2272
rect 4927 2250 4957 2272
rect 5049 2250 5079 2272
rect 5783 2250 5813 2272
rect 643 2217 659 2244
rect 625 2210 659 2217
rect 693 2217 709 2244
rect 1627 2234 1693 2250
rect 693 2210 727 2217
rect 625 2187 727 2210
rect 625 2172 655 2187
rect 697 2172 727 2187
rect 1627 2200 1643 2234
rect 1677 2200 1693 2234
rect 1627 2184 1693 2200
rect 2359 2234 2425 2250
rect 2359 2200 2375 2234
rect 2409 2200 2425 2234
rect 2359 2184 2425 2200
rect 2481 2234 2547 2250
rect 2481 2200 2497 2234
rect 2531 2200 2547 2234
rect 2481 2184 2547 2200
rect 3571 2234 3637 2250
rect 3571 2200 3587 2234
rect 3621 2200 3637 2234
rect 3571 2184 3637 2200
rect 3693 2234 3759 2250
rect 3693 2200 3709 2234
rect 3743 2200 3759 2234
rect 3693 2184 3759 2200
rect 4909 2234 4975 2250
rect 4909 2200 4925 2234
rect 4959 2200 4975 2234
rect 4909 2184 4975 2200
rect 5031 2234 5097 2250
rect 5031 2200 5047 2234
rect 5081 2200 5097 2234
rect 5031 2184 5097 2200
rect 5765 2234 5831 2250
rect 5765 2200 5781 2234
rect 5815 2200 5831 2234
rect 6435 2219 6465 2273
rect 6527 2247 6557 2273
rect 6623 2247 6653 2273
rect 7352 2244 7418 2260
rect 8354 2250 8384 2272
rect 9086 2250 9116 2272
rect 9208 2250 9238 2272
rect 10298 2250 10328 2272
rect 10420 2250 10450 2272
rect 11636 2250 11666 2272
rect 11758 2250 11788 2272
rect 12492 2250 12522 2272
rect 5765 2184 5831 2200
rect 7352 2217 7368 2244
rect 7334 2210 7368 2217
rect 7402 2217 7418 2244
rect 8336 2234 8402 2250
rect 7402 2210 7436 2217
rect 7334 2187 7436 2210
rect 7334 2172 7364 2187
rect 7406 2172 7436 2187
rect 8336 2200 8352 2234
rect 8386 2200 8402 2234
rect 8336 2184 8402 2200
rect 9068 2234 9134 2250
rect 9068 2200 9084 2234
rect 9118 2200 9134 2234
rect 9068 2184 9134 2200
rect 9190 2234 9256 2250
rect 9190 2200 9206 2234
rect 9240 2200 9256 2234
rect 9190 2184 9256 2200
rect 10280 2234 10346 2250
rect 10280 2200 10296 2234
rect 10330 2200 10346 2234
rect 10280 2184 10346 2200
rect 10402 2234 10468 2250
rect 10402 2200 10418 2234
rect 10452 2200 10468 2234
rect 10402 2184 10468 2200
rect 11618 2234 11684 2250
rect 11618 2200 11634 2234
rect 11668 2200 11684 2234
rect 11618 2184 11684 2200
rect 11740 2234 11806 2250
rect 11740 2200 11756 2234
rect 11790 2200 11806 2234
rect 11740 2184 11806 2200
rect 12474 2234 12540 2250
rect 12474 2200 12490 2234
rect 12524 2200 12540 2234
rect 13144 2219 13174 2273
rect 13236 2247 13266 2273
rect 13332 2247 13362 2273
rect 12474 2184 12540 2200
rect 6435 2108 6465 2135
rect 13144 2108 13174 2135
rect 625 2034 655 2088
rect 697 2034 727 2088
rect 7334 2034 7364 2088
rect 7406 2034 7436 2088
rect 625 1896 655 1950
rect 697 1896 727 1950
rect 7334 1896 7364 1950
rect 7406 1896 7436 1950
rect 625 1758 655 1812
rect 697 1758 727 1812
rect 7334 1758 7364 1812
rect 7406 1758 7436 1812
rect 625 1620 655 1674
rect 697 1620 727 1674
rect 7334 1620 7364 1674
rect 7406 1620 7436 1674
rect 625 1482 655 1536
rect 697 1482 727 1536
rect 7334 1482 7364 1536
rect 7406 1482 7436 1536
rect 625 1344 655 1398
rect 697 1344 727 1398
rect 7334 1344 7364 1398
rect 7406 1344 7436 1398
rect 625 1206 655 1260
rect 697 1206 727 1260
rect 7334 1206 7364 1260
rect 7406 1206 7436 1260
rect 625 1096 655 1122
rect 697 1096 727 1122
rect 7334 1096 7364 1122
rect 7406 1096 7436 1122
rect 6028 199 6058 225
rect 6100 199 6130 225
rect 12737 199 12767 225
rect 12809 199 12839 225
rect 6028 61 6058 115
rect 6100 61 6130 115
rect 12737 61 12767 115
rect 12809 61 12839 115
rect 6028 -77 6058 -23
rect 6100 -77 6130 -23
rect 12737 -77 12767 -23
rect 12809 -77 12839 -23
rect 6028 -215 6058 -161
rect 6100 -215 6130 -161
rect 12737 -215 12767 -161
rect 12809 -215 12839 -161
rect 6028 -353 6058 -299
rect 6100 -353 6130 -299
rect 12737 -353 12767 -299
rect 12809 -353 12839 -299
rect 6028 -491 6058 -437
rect 6100 -491 6130 -437
rect 12737 -491 12767 -437
rect 12809 -491 12839 -437
rect 6028 -629 6058 -575
rect 6100 -629 6130 -575
rect 12737 -629 12767 -575
rect 12809 -629 12839 -575
rect 6028 -767 6058 -713
rect 6100 -767 6130 -713
rect 12737 -767 12767 -713
rect 12809 -767 12839 -713
rect 290 -814 320 -787
rect 6999 -814 7029 -787
rect 924 -879 990 -863
rect 102 -952 132 -926
rect 198 -952 228 -926
rect 290 -952 320 -898
rect 924 -913 940 -879
rect 974 -913 990 -879
rect 924 -929 990 -913
rect 1658 -879 1724 -863
rect 1658 -913 1674 -879
rect 1708 -913 1724 -879
rect 1658 -929 1724 -913
rect 1780 -879 1846 -863
rect 1780 -913 1796 -879
rect 1830 -913 1846 -879
rect 1780 -929 1846 -913
rect 2996 -879 3062 -863
rect 2996 -913 3012 -879
rect 3046 -913 3062 -879
rect 2996 -929 3062 -913
rect 3118 -879 3184 -863
rect 3118 -913 3134 -879
rect 3168 -913 3184 -879
rect 3118 -929 3184 -913
rect 4208 -879 4274 -863
rect 4208 -913 4224 -879
rect 4258 -913 4274 -879
rect 4208 -929 4274 -913
rect 4330 -879 4396 -863
rect 4330 -913 4346 -879
rect 4380 -913 4396 -879
rect 4330 -929 4396 -913
rect 5062 -879 5128 -863
rect 5062 -913 5078 -879
rect 5112 -913 5128 -879
rect 6028 -866 6058 -851
rect 6100 -866 6130 -851
rect 6028 -889 6130 -866
rect 6028 -896 6062 -889
rect 5062 -929 5128 -913
rect 6046 -923 6062 -896
rect 6096 -896 6130 -889
rect 6096 -923 6112 -896
rect 7633 -879 7699 -863
rect 942 -951 972 -929
rect 1676 -951 1706 -929
rect 1798 -951 1828 -929
rect 3014 -951 3044 -929
rect 3136 -951 3166 -929
rect 4226 -951 4256 -929
rect 4348 -951 4378 -929
rect 5080 -951 5110 -929
rect 6046 -939 6112 -923
rect 6811 -952 6841 -926
rect 6907 -952 6937 -926
rect 6999 -952 7029 -898
rect 7633 -913 7649 -879
rect 7683 -913 7699 -879
rect 7633 -929 7699 -913
rect 8367 -879 8433 -863
rect 8367 -913 8383 -879
rect 8417 -913 8433 -879
rect 8367 -929 8433 -913
rect 8489 -879 8555 -863
rect 8489 -913 8505 -879
rect 8539 -913 8555 -879
rect 8489 -929 8555 -913
rect 9705 -879 9771 -863
rect 9705 -913 9721 -879
rect 9755 -913 9771 -879
rect 9705 -929 9771 -913
rect 9827 -879 9893 -863
rect 9827 -913 9843 -879
rect 9877 -913 9893 -879
rect 9827 -929 9893 -913
rect 10917 -879 10983 -863
rect 10917 -913 10933 -879
rect 10967 -913 10983 -879
rect 10917 -929 10983 -913
rect 11039 -879 11105 -863
rect 11039 -913 11055 -879
rect 11089 -913 11105 -879
rect 11039 -929 11105 -913
rect 11771 -879 11837 -863
rect 11771 -913 11787 -879
rect 11821 -913 11837 -879
rect 12737 -866 12767 -851
rect 12809 -866 12839 -851
rect 12737 -889 12839 -866
rect 12737 -896 12771 -889
rect 11771 -929 11837 -913
rect 12755 -923 12771 -896
rect 12805 -896 12839 -889
rect 12805 -923 12821 -896
rect 7651 -951 7681 -929
rect 8385 -951 8415 -929
rect 8507 -951 8537 -929
rect 9723 -951 9753 -929
rect 9845 -951 9875 -929
rect 10935 -951 10965 -929
rect 11057 -951 11087 -929
rect 11789 -951 11819 -929
rect 12755 -939 12821 -923
rect 102 -1051 132 -1036
rect 198 -1051 228 -1036
rect 102 -1058 228 -1051
rect 290 -1057 320 -1036
rect 102 -1074 246 -1058
rect 102 -1108 196 -1074
rect 230 -1108 246 -1074
rect 102 -1124 246 -1108
rect 290 -1076 449 -1057
rect 942 -1061 972 -1035
rect 1676 -1061 1706 -1035
rect 1798 -1061 1828 -1035
rect 3014 -1061 3044 -1035
rect 3136 -1061 3166 -1035
rect 4226 -1061 4256 -1035
rect 4348 -1061 4378 -1035
rect 5080 -1061 5110 -1035
rect 6811 -1051 6841 -1036
rect 6907 -1051 6937 -1036
rect 6811 -1058 6937 -1051
rect 6999 -1057 7029 -1036
rect 290 -1110 403 -1076
rect 437 -1110 449 -1076
rect 102 -1130 228 -1124
rect 102 -1155 132 -1130
rect 198 -1155 228 -1130
rect 290 -1130 449 -1110
rect 6811 -1074 6955 -1058
rect 6811 -1108 6905 -1074
rect 6939 -1108 6955 -1074
rect 290 -1155 320 -1130
rect 939 -1152 969 -1124
rect 1065 -1152 1095 -1124
rect 2151 -1152 2181 -1124
rect 2277 -1152 2307 -1124
rect 3363 -1152 3393 -1124
rect 3489 -1152 3519 -1124
rect 4575 -1152 4605 -1124
rect 4701 -1152 4731 -1124
rect 5433 -1149 5463 -1121
rect 6811 -1124 6955 -1108
rect 6999 -1076 7158 -1057
rect 7651 -1061 7681 -1035
rect 8385 -1061 8415 -1035
rect 8507 -1061 8537 -1035
rect 9723 -1061 9753 -1035
rect 9845 -1061 9875 -1035
rect 10935 -1061 10965 -1035
rect 11057 -1061 11087 -1035
rect 11789 -1061 11819 -1035
rect 6999 -1110 7112 -1076
rect 7146 -1110 7158 -1076
rect 6811 -1130 6937 -1124
rect 6811 -1155 6841 -1130
rect 6907 -1155 6937 -1130
rect 6999 -1130 7158 -1110
rect 6999 -1155 7029 -1130
rect 7648 -1152 7678 -1124
rect 7774 -1152 7804 -1124
rect 8860 -1152 8890 -1124
rect 8986 -1152 9016 -1124
rect 10072 -1152 10102 -1124
rect 10198 -1152 10228 -1124
rect 11284 -1152 11314 -1124
rect 11410 -1152 11440 -1124
rect 12142 -1149 12172 -1121
rect 102 -1270 132 -1239
rect 198 -1265 228 -1239
rect 290 -1293 320 -1239
rect 939 -1267 969 -1236
rect 1065 -1267 1095 -1236
rect 2151 -1267 2181 -1236
rect 2277 -1267 2307 -1236
rect 3363 -1267 3393 -1236
rect 3489 -1267 3519 -1236
rect 4575 -1267 4605 -1236
rect 4701 -1267 4731 -1236
rect 5433 -1264 5463 -1233
rect 921 -1283 987 -1267
rect 921 -1317 937 -1283
rect 971 -1317 987 -1283
rect 921 -1333 987 -1317
rect 1047 -1283 1113 -1267
rect 1047 -1317 1063 -1283
rect 1097 -1317 1113 -1283
rect 1047 -1333 1113 -1317
rect 2133 -1283 2199 -1267
rect 2133 -1317 2149 -1283
rect 2183 -1317 2199 -1283
rect 2133 -1333 2199 -1317
rect 2259 -1283 2325 -1267
rect 2259 -1317 2275 -1283
rect 2309 -1317 2325 -1283
rect 2259 -1333 2325 -1317
rect 3345 -1283 3411 -1267
rect 3345 -1317 3361 -1283
rect 3395 -1317 3411 -1283
rect 3345 -1333 3411 -1317
rect 3471 -1283 3537 -1267
rect 3471 -1317 3487 -1283
rect 3521 -1317 3537 -1283
rect 3471 -1333 3537 -1317
rect 4557 -1283 4623 -1267
rect 4557 -1317 4573 -1283
rect 4607 -1317 4623 -1283
rect 4557 -1333 4623 -1317
rect 4683 -1283 4749 -1267
rect 4683 -1317 4699 -1283
rect 4733 -1317 4749 -1283
rect 4683 -1333 4749 -1317
rect 5415 -1280 5481 -1264
rect 5415 -1314 5431 -1280
rect 5465 -1314 5481 -1280
rect 6353 -1281 6383 -1255
rect 6543 -1281 6573 -1255
rect 6811 -1270 6841 -1239
rect 6907 -1265 6937 -1239
rect 5415 -1330 5481 -1314
rect 290 -1408 320 -1377
rect 6999 -1293 7029 -1239
rect 7648 -1267 7678 -1236
rect 7774 -1267 7804 -1236
rect 8860 -1267 8890 -1236
rect 8986 -1267 9016 -1236
rect 10072 -1267 10102 -1236
rect 10198 -1267 10228 -1236
rect 11284 -1267 11314 -1236
rect 11410 -1267 11440 -1236
rect 12142 -1264 12172 -1233
rect 7630 -1283 7696 -1267
rect 7630 -1317 7646 -1283
rect 7680 -1317 7696 -1283
rect 7630 -1333 7696 -1317
rect 7756 -1283 7822 -1267
rect 7756 -1317 7772 -1283
rect 7806 -1317 7822 -1283
rect 7756 -1333 7822 -1317
rect 8842 -1283 8908 -1267
rect 8842 -1317 8858 -1283
rect 8892 -1317 8908 -1283
rect 8842 -1333 8908 -1317
rect 8968 -1283 9034 -1267
rect 8968 -1317 8984 -1283
rect 9018 -1317 9034 -1283
rect 8968 -1333 9034 -1317
rect 10054 -1283 10120 -1267
rect 10054 -1317 10070 -1283
rect 10104 -1317 10120 -1283
rect 10054 -1333 10120 -1317
rect 10180 -1283 10246 -1267
rect 10180 -1317 10196 -1283
rect 10230 -1317 10246 -1283
rect 10180 -1333 10246 -1317
rect 11266 -1283 11332 -1267
rect 11266 -1317 11282 -1283
rect 11316 -1317 11332 -1283
rect 11266 -1333 11332 -1317
rect 11392 -1283 11458 -1267
rect 11392 -1317 11408 -1283
rect 11442 -1317 11458 -1283
rect 11392 -1333 11458 -1317
rect 12124 -1280 12190 -1264
rect 12124 -1314 12140 -1280
rect 12174 -1314 12190 -1280
rect 13062 -1281 13092 -1255
rect 13252 -1281 13282 -1255
rect 12124 -1330 12190 -1314
rect 6999 -1408 7029 -1377
rect 6353 -1433 6383 -1411
rect 6297 -1449 6383 -1433
rect 6297 -1483 6313 -1449
rect 6347 -1483 6383 -1449
rect 6297 -1499 6383 -1483
rect 6057 -1523 6123 -1507
rect 6057 -1557 6073 -1523
rect 6107 -1557 6123 -1523
rect 6353 -1531 6383 -1499
rect 6543 -1433 6573 -1411
rect 13062 -1433 13092 -1411
rect 6543 -1449 6629 -1433
rect 6543 -1483 6579 -1449
rect 6613 -1483 6629 -1449
rect 6543 -1499 6629 -1483
rect 13006 -1449 13092 -1433
rect 13006 -1483 13022 -1449
rect 13056 -1483 13092 -1449
rect 13006 -1499 13092 -1483
rect 6543 -1531 6573 -1499
rect 12766 -1523 12832 -1507
rect 6057 -1573 6123 -1557
rect 6075 -1604 6105 -1573
rect 6075 -1742 6105 -1688
rect 12766 -1557 12782 -1523
rect 12816 -1557 12832 -1523
rect 13062 -1531 13092 -1499
rect 13252 -1433 13282 -1411
rect 13252 -1449 13338 -1433
rect 13252 -1483 13288 -1449
rect 13322 -1483 13338 -1449
rect 13252 -1499 13338 -1483
rect 13252 -1531 13282 -1499
rect 12766 -1573 12832 -1557
rect 12784 -1604 12814 -1573
rect 6353 -1757 6383 -1731
rect 6543 -1757 6573 -1731
rect 12784 -1742 12814 -1688
rect 6075 -1880 6105 -1826
rect 13062 -1757 13092 -1731
rect 13252 -1757 13282 -1731
rect 12784 -1880 12814 -1826
rect 6075 -2018 6105 -1964
rect 12784 -2018 12814 -1964
rect 6075 -2156 6105 -2102
rect 12784 -2156 12814 -2102
rect 6075 -2294 6105 -2240
rect 12784 -2294 12814 -2240
rect 6075 -2408 6105 -2378
rect 12784 -2408 12814 -2378
<< polycont >>
rect 142 2770 176 2804
rect 648 2844 682 2878
rect 408 2770 442 2804
rect 6851 2770 6885 2804
rect 7357 2844 7391 2878
rect 7117 2770 7151 2804
rect 1290 2601 1324 2635
rect 2022 2604 2056 2638
rect 2148 2604 2182 2638
rect 3234 2604 3268 2638
rect 3360 2604 3394 2638
rect 4446 2604 4480 2638
rect 4572 2604 4606 2638
rect 5658 2604 5692 2638
rect 5784 2604 5818 2638
rect 7999 2601 8033 2635
rect 8731 2604 8765 2638
rect 8857 2604 8891 2638
rect 9943 2604 9977 2638
rect 10069 2604 10103 2638
rect 11155 2604 11189 2638
rect 11281 2604 11315 2638
rect 12367 2604 12401 2638
rect 12493 2604 12527 2638
rect 6318 2397 6352 2431
rect 6525 2395 6559 2429
rect 13027 2397 13061 2431
rect 13234 2395 13268 2429
rect 659 2210 693 2244
rect 1643 2200 1677 2234
rect 2375 2200 2409 2234
rect 2497 2200 2531 2234
rect 3587 2200 3621 2234
rect 3709 2200 3743 2234
rect 4925 2200 4959 2234
rect 5047 2200 5081 2234
rect 5781 2200 5815 2234
rect 7368 2210 7402 2244
rect 8352 2200 8386 2234
rect 9084 2200 9118 2234
rect 9206 2200 9240 2234
rect 10296 2200 10330 2234
rect 10418 2200 10452 2234
rect 11634 2200 11668 2234
rect 11756 2200 11790 2234
rect 12490 2200 12524 2234
rect 940 -913 974 -879
rect 1674 -913 1708 -879
rect 1796 -913 1830 -879
rect 3012 -913 3046 -879
rect 3134 -913 3168 -879
rect 4224 -913 4258 -879
rect 4346 -913 4380 -879
rect 5078 -913 5112 -879
rect 6062 -923 6096 -889
rect 7649 -913 7683 -879
rect 8383 -913 8417 -879
rect 8505 -913 8539 -879
rect 9721 -913 9755 -879
rect 9843 -913 9877 -879
rect 10933 -913 10967 -879
rect 11055 -913 11089 -879
rect 11787 -913 11821 -879
rect 12771 -923 12805 -889
rect 196 -1108 230 -1074
rect 403 -1110 437 -1076
rect 6905 -1108 6939 -1074
rect 7112 -1110 7146 -1076
rect 937 -1317 971 -1283
rect 1063 -1317 1097 -1283
rect 2149 -1317 2183 -1283
rect 2275 -1317 2309 -1283
rect 3361 -1317 3395 -1283
rect 3487 -1317 3521 -1283
rect 4573 -1317 4607 -1283
rect 4699 -1317 4733 -1283
rect 5431 -1314 5465 -1280
rect 7646 -1317 7680 -1283
rect 7772 -1317 7806 -1283
rect 8858 -1317 8892 -1283
rect 8984 -1317 9018 -1283
rect 10070 -1317 10104 -1283
rect 10196 -1317 10230 -1283
rect 11282 -1317 11316 -1283
rect 11408 -1317 11442 -1283
rect 12140 -1314 12174 -1280
rect 6313 -1483 6347 -1449
rect 6073 -1557 6107 -1523
rect 6579 -1483 6613 -1449
rect 13022 -1483 13056 -1449
rect 12782 -1557 12816 -1523
rect 13288 -1483 13322 -1449
<< locali >>
rect 734 3711 1404 3729
rect 734 3703 850 3711
rect 604 3687 638 3703
rect 604 3611 638 3627
rect 692 3687 850 3703
rect 726 3677 850 3687
rect 886 3677 930 3711
rect 966 3677 1010 3711
rect 1046 3677 1090 3711
rect 1126 3677 1170 3711
rect 1206 3677 1250 3711
rect 1286 3677 1404 3711
rect 726 3663 1404 3677
rect 1466 3714 6374 3732
rect 1466 3680 1582 3714
rect 1618 3680 1662 3714
rect 1698 3680 1742 3714
rect 1778 3680 1822 3714
rect 1858 3680 1902 3714
rect 1938 3680 1982 3714
rect 2018 3680 2186 3714
rect 2222 3680 2266 3714
rect 2302 3680 2346 3714
rect 2382 3680 2426 3714
rect 2462 3680 2506 3714
rect 2542 3680 2586 3714
rect 2622 3680 2794 3714
rect 2830 3680 2874 3714
rect 2910 3680 2954 3714
rect 2990 3680 3034 3714
rect 3070 3680 3114 3714
rect 3150 3680 3194 3714
rect 3230 3680 3398 3714
rect 3434 3680 3478 3714
rect 3514 3680 3558 3714
rect 3594 3680 3638 3714
rect 3674 3680 3718 3714
rect 3754 3680 3798 3714
rect 3834 3680 4006 3714
rect 4042 3680 4086 3714
rect 4122 3680 4166 3714
rect 4202 3680 4246 3714
rect 4282 3680 4326 3714
rect 4362 3680 4406 3714
rect 4442 3680 4610 3714
rect 4646 3680 4690 3714
rect 4726 3680 4770 3714
rect 4806 3680 4850 3714
rect 4886 3680 4930 3714
rect 4966 3680 5010 3714
rect 5046 3680 5218 3714
rect 5254 3680 5298 3714
rect 5334 3680 5378 3714
rect 5414 3680 5458 3714
rect 5494 3680 5538 3714
rect 5574 3680 5618 3714
rect 5654 3680 5822 3714
rect 5858 3680 5902 3714
rect 5938 3680 5982 3714
rect 6018 3680 6062 3714
rect 6098 3680 6142 3714
rect 6178 3680 6222 3714
rect 6258 3680 6374 3714
rect 7443 3711 8113 3729
rect 7443 3703 7559 3711
rect 1466 3666 6374 3680
rect 6538 3663 6624 3689
rect 726 3627 862 3663
rect 692 3622 862 3627
rect 692 3611 726 3622
rect 604 3549 638 3565
rect 604 3473 638 3489
rect 692 3549 726 3565
rect 805 3558 862 3622
rect 6538 3629 6564 3663
rect 6598 3629 6624 3663
rect 6538 3603 6624 3629
rect 7015 3666 7101 3692
rect 7015 3632 7041 3666
rect 7075 3632 7101 3666
rect 7015 3606 7101 3632
rect 7313 3687 7347 3703
rect 7313 3611 7347 3627
rect 7401 3687 7559 3703
rect 7435 3677 7559 3687
rect 7595 3677 7639 3711
rect 7675 3677 7719 3711
rect 7755 3677 7799 3711
rect 7835 3677 7879 3711
rect 7915 3677 7959 3711
rect 7995 3677 8113 3711
rect 7435 3663 8113 3677
rect 8175 3714 13083 3732
rect 8175 3680 8291 3714
rect 8327 3680 8371 3714
rect 8407 3680 8451 3714
rect 8487 3680 8531 3714
rect 8567 3680 8611 3714
rect 8647 3680 8691 3714
rect 8727 3680 8895 3714
rect 8931 3680 8975 3714
rect 9011 3680 9055 3714
rect 9091 3680 9135 3714
rect 9171 3680 9215 3714
rect 9251 3680 9295 3714
rect 9331 3680 9503 3714
rect 9539 3680 9583 3714
rect 9619 3680 9663 3714
rect 9699 3680 9743 3714
rect 9779 3680 9823 3714
rect 9859 3680 9903 3714
rect 9939 3680 10107 3714
rect 10143 3680 10187 3714
rect 10223 3680 10267 3714
rect 10303 3680 10347 3714
rect 10383 3680 10427 3714
rect 10463 3680 10507 3714
rect 10543 3680 10715 3714
rect 10751 3680 10795 3714
rect 10831 3680 10875 3714
rect 10911 3680 10955 3714
rect 10991 3680 11035 3714
rect 11071 3680 11115 3714
rect 11151 3680 11319 3714
rect 11355 3680 11399 3714
rect 11435 3680 11479 3714
rect 11515 3680 11559 3714
rect 11595 3680 11639 3714
rect 11675 3680 11719 3714
rect 11755 3680 11927 3714
rect 11963 3680 12007 3714
rect 12043 3680 12087 3714
rect 12123 3680 12167 3714
rect 12203 3680 12247 3714
rect 12283 3680 12327 3714
rect 12363 3680 12531 3714
rect 12567 3680 12611 3714
rect 12647 3680 12691 3714
rect 12727 3680 12771 3714
rect 12807 3680 12851 3714
rect 12887 3680 12931 3714
rect 12967 3680 13083 3714
rect 8175 3666 13083 3680
rect 13247 3663 13333 3689
rect 7435 3627 7571 3663
rect 7401 3622 7571 3627
rect 7401 3611 7435 3622
rect 692 3473 726 3489
rect 792 3533 875 3558
rect 7313 3549 7347 3565
rect 792 3498 817 3533
rect 851 3498 875 3533
rect 792 3474 875 3498
rect 6543 3519 6629 3545
rect 6543 3485 6569 3519
rect 6603 3485 6629 3519
rect 6543 3459 6629 3485
rect 7004 3494 7090 3520
rect 7004 3460 7030 3494
rect 7064 3460 7090 3494
rect 7313 3473 7347 3489
rect 7401 3549 7435 3565
rect 7514 3558 7571 3622
rect 13247 3629 13273 3663
rect 13307 3629 13333 3663
rect 13247 3603 13333 3629
rect 7401 3473 7435 3489
rect 7501 3533 7584 3558
rect 7501 3498 7526 3533
rect 7560 3498 7584 3533
rect 7501 3474 7584 3498
rect 13252 3519 13338 3545
rect 13252 3485 13278 3519
rect 13312 3485 13338 3519
rect 7004 3434 7090 3460
rect 13252 3459 13338 3485
rect 604 3411 638 3427
rect 604 3335 638 3351
rect 692 3411 726 3427
rect 7313 3411 7347 3427
rect 692 3335 726 3351
rect 6544 3367 6630 3393
rect 6544 3333 6570 3367
rect 6604 3333 6630 3367
rect 7313 3335 7347 3351
rect 7401 3411 7435 3427
rect 7401 3335 7435 3351
rect 13253 3367 13339 3393
rect 6544 3307 6630 3333
rect 13253 3333 13279 3367
rect 13313 3333 13339 3367
rect 7004 3302 7090 3328
rect 13253 3307 13339 3333
rect 604 3273 638 3289
rect 604 3197 638 3213
rect 692 3273 726 3289
rect 7004 3268 7030 3302
rect 7064 3268 7090 3302
rect 7004 3242 7090 3268
rect 7313 3273 7347 3289
rect 692 3197 726 3213
rect 6544 3197 6630 3223
rect 7313 3197 7347 3213
rect 7401 3273 7435 3289
rect 7401 3197 7435 3213
rect 13253 3197 13339 3223
rect 6544 3163 6570 3197
rect 6604 3163 6630 3197
rect 120 3116 136 3145
rect 62 3082 91 3116
rect 125 3111 136 3116
rect 170 3116 186 3145
rect 250 3116 266 3145
rect 300 3116 320 3145
rect 396 3116 412 3145
rect 170 3111 183 3116
rect 125 3082 183 3111
rect 217 3111 266 3116
rect 217 3082 275 3111
rect 309 3082 367 3116
rect 401 3111 412 3116
rect 446 3116 466 3145
rect 604 3135 638 3151
rect 446 3111 459 3116
rect 401 3082 459 3111
rect 493 3082 522 3116
rect 130 3040 172 3082
rect 130 3006 138 3040
rect 130 2972 172 3006
rect 130 2938 138 2972
rect 130 2904 172 2938
rect 130 2870 138 2904
rect 130 2854 172 2870
rect 206 3040 272 3048
rect 206 3006 222 3040
rect 256 3006 272 3040
rect 206 2973 272 3006
rect 206 2939 219 2973
rect 253 2972 272 2973
rect 206 2938 222 2939
rect 256 2938 272 2972
rect 206 2904 272 2938
rect 206 2870 222 2904
rect 256 2870 272 2904
rect 206 2852 272 2870
rect 126 2808 192 2818
rect 126 2774 138 2808
rect 172 2804 192 2808
rect 126 2770 142 2774
rect 176 2770 192 2804
rect 126 2720 172 2736
rect 226 2732 272 2852
rect 126 2686 138 2720
rect 126 2652 172 2686
rect 126 2618 138 2652
rect 126 2572 172 2618
rect 206 2720 272 2732
rect 206 2686 222 2720
rect 256 2686 272 2720
rect 206 2652 272 2686
rect 206 2618 222 2652
rect 256 2618 272 2652
rect 206 2606 272 2618
rect 312 3040 378 3048
rect 312 3006 328 3040
rect 362 3006 378 3040
rect 312 2972 378 3006
rect 312 2938 328 2972
rect 362 2938 378 2972
rect 312 2918 378 2938
rect 312 2870 328 2918
rect 362 2870 378 2918
rect 312 2852 378 2870
rect 412 3040 454 3082
rect 604 3059 638 3075
rect 692 3135 726 3151
rect 6544 3137 6630 3163
rect 13253 3163 13279 3197
rect 13313 3163 13339 3197
rect 6829 3116 6845 3145
rect 6771 3082 6800 3116
rect 6834 3111 6845 3116
rect 6879 3116 6895 3145
rect 6959 3116 6975 3145
rect 7009 3116 7029 3145
rect 7105 3116 7121 3145
rect 6879 3111 6892 3116
rect 6834 3082 6892 3111
rect 6926 3111 6975 3116
rect 6926 3082 6984 3111
rect 7018 3082 7076 3116
rect 7110 3111 7121 3116
rect 7155 3116 7175 3145
rect 7313 3135 7347 3151
rect 7155 3111 7168 3116
rect 7110 3082 7168 3111
rect 7202 3082 7231 3116
rect 692 3059 726 3075
rect 446 3006 454 3040
rect 6543 3040 6629 3066
rect 412 2972 454 3006
rect 446 2938 454 2972
rect 412 2904 454 2938
rect 604 2997 638 3013
rect 604 2921 638 2937
rect 692 2997 726 3013
rect 6543 3006 6569 3040
rect 6603 3006 6629 3040
rect 6543 2980 6629 3006
rect 6839 3040 6881 3082
rect 6839 3006 6847 3040
rect 692 2921 726 2937
rect 6839 2972 6881 3006
rect 6839 2938 6847 2972
rect 446 2870 454 2904
rect 6839 2904 6881 2938
rect 412 2854 454 2870
rect 312 2732 358 2852
rect 632 2844 648 2878
rect 682 2844 698 2878
rect 6839 2870 6847 2904
rect 6839 2854 6881 2870
rect 6915 3040 6981 3048
rect 6915 3006 6931 3040
rect 6965 3006 6981 3040
rect 6915 2973 6981 3006
rect 6915 2939 6928 2973
rect 6962 2972 6981 2973
rect 6915 2938 6931 2939
rect 6965 2938 6981 2972
rect 6915 2904 6981 2938
rect 6915 2870 6931 2904
rect 6965 2870 6981 2904
rect 6915 2852 6981 2870
rect 392 2807 458 2818
rect 392 2804 412 2807
rect 392 2770 408 2804
rect 446 2773 458 2807
rect 442 2770 458 2773
rect 542 2808 591 2820
rect 542 2774 551 2808
rect 585 2803 591 2808
rect 6835 2808 6901 2818
rect 585 2774 874 2803
rect 542 2768 874 2774
rect 6835 2774 6847 2808
rect 6881 2804 6901 2808
rect 6835 2770 6851 2774
rect 6885 2770 6901 2804
rect 542 2761 591 2768
rect 839 2745 874 2768
rect 312 2720 378 2732
rect 312 2686 328 2720
rect 362 2686 378 2720
rect 312 2652 378 2686
rect 312 2618 328 2652
rect 362 2618 378 2652
rect 312 2606 378 2618
rect 412 2720 458 2736
rect 839 2733 888 2745
rect 446 2686 458 2720
rect 412 2652 458 2686
rect 580 2715 629 2727
rect 580 2681 589 2715
rect 623 2681 790 2715
rect 839 2699 848 2733
rect 882 2699 888 2733
rect 6835 2720 6881 2736
rect 6935 2732 6981 2852
rect 839 2686 888 2699
rect 6389 2686 6423 2702
rect 580 2668 629 2681
rect 446 2618 458 2652
rect 412 2572 458 2618
rect 749 2639 790 2681
rect 840 2640 889 2652
rect 840 2639 849 2640
rect 749 2606 849 2639
rect 883 2606 889 2640
rect 749 2605 889 2606
rect 840 2593 889 2605
rect 1274 2601 1290 2635
rect 1324 2601 1340 2635
rect 2006 2604 2022 2638
rect 2056 2604 2072 2638
rect 2132 2604 2148 2638
rect 2182 2604 2198 2638
rect 3218 2604 3234 2638
rect 3268 2604 3284 2638
rect 3344 2604 3360 2638
rect 3394 2604 3410 2638
rect 4430 2604 4446 2638
rect 4480 2604 4496 2638
rect 4556 2604 4572 2638
rect 4606 2604 4622 2638
rect 5642 2604 5658 2638
rect 5692 2604 5708 2638
rect 5768 2604 5784 2638
rect 5818 2604 5834 2638
rect 6389 2610 6423 2626
rect 6477 2686 6511 2702
rect 6477 2610 6511 2626
rect 6835 2686 6847 2720
rect 6835 2652 6881 2686
rect 6835 2618 6847 2652
rect 6835 2572 6881 2618
rect 6915 2720 6981 2732
rect 6915 2686 6931 2720
rect 6965 2686 6981 2720
rect 6915 2652 6981 2686
rect 6915 2618 6931 2652
rect 6965 2618 6981 2652
rect 6915 2606 6981 2618
rect 7021 3040 7087 3048
rect 7021 3006 7037 3040
rect 7071 3006 7087 3040
rect 7021 2972 7087 3006
rect 7021 2938 7037 2972
rect 7071 2938 7087 2972
rect 7021 2918 7087 2938
rect 7021 2870 7037 2918
rect 7071 2870 7087 2918
rect 7021 2852 7087 2870
rect 7121 3040 7163 3082
rect 7313 3059 7347 3075
rect 7401 3135 7435 3151
rect 13253 3137 13339 3163
rect 7401 3059 7435 3075
rect 7155 3006 7163 3040
rect 13252 3040 13338 3066
rect 7121 2972 7163 3006
rect 7155 2938 7163 2972
rect 7121 2904 7163 2938
rect 7313 2997 7347 3013
rect 7313 2921 7347 2937
rect 7401 2997 7435 3013
rect 13252 3006 13278 3040
rect 13312 3006 13338 3040
rect 13252 2980 13338 3006
rect 7401 2921 7435 2937
rect 7155 2870 7163 2904
rect 7121 2854 7163 2870
rect 7021 2732 7067 2852
rect 7341 2844 7357 2878
rect 7391 2844 7407 2878
rect 7101 2807 7167 2818
rect 7101 2804 7121 2807
rect 7101 2770 7117 2804
rect 7155 2773 7167 2807
rect 7151 2770 7167 2773
rect 7251 2808 7300 2820
rect 7251 2774 7260 2808
rect 7294 2803 7300 2808
rect 7294 2774 7583 2803
rect 7251 2768 7583 2774
rect 7251 2761 7300 2768
rect 7548 2745 7583 2768
rect 7021 2720 7087 2732
rect 7021 2686 7037 2720
rect 7071 2686 7087 2720
rect 7021 2652 7087 2686
rect 7021 2618 7037 2652
rect 7071 2618 7087 2652
rect 7021 2606 7087 2618
rect 7121 2720 7167 2736
rect 7548 2733 7597 2745
rect 7155 2686 7167 2720
rect 7121 2652 7167 2686
rect 7289 2715 7338 2727
rect 7289 2681 7298 2715
rect 7332 2681 7499 2715
rect 7548 2699 7557 2733
rect 7591 2699 7597 2733
rect 7548 2686 7597 2699
rect 13098 2686 13132 2702
rect 7289 2668 7338 2681
rect 7155 2618 7167 2652
rect 7121 2572 7167 2618
rect 7458 2639 7499 2681
rect 7549 2640 7598 2652
rect 7549 2639 7558 2640
rect 7458 2606 7558 2639
rect 7592 2606 7598 2640
rect 7458 2605 7598 2606
rect 7549 2593 7598 2605
rect 7983 2601 7999 2635
rect 8033 2601 8049 2635
rect 8715 2604 8731 2638
rect 8765 2604 8781 2638
rect 8841 2604 8857 2638
rect 8891 2604 8907 2638
rect 9927 2604 9943 2638
rect 9977 2604 9993 2638
rect 10053 2604 10069 2638
rect 10103 2604 10119 2638
rect 11139 2604 11155 2638
rect 11189 2604 11205 2638
rect 11265 2604 11281 2638
rect 11315 2604 11331 2638
rect 12351 2604 12367 2638
rect 12401 2604 12417 2638
rect 12477 2604 12493 2638
rect 12527 2604 12543 2638
rect 13098 2610 13132 2626
rect 13186 2686 13220 2702
rect 13186 2610 13220 2626
rect 62 2538 91 2572
rect 125 2543 183 2572
rect 217 2543 275 2572
rect 125 2538 156 2543
rect 217 2538 274 2543
rect 309 2538 367 2572
rect 401 2543 459 2572
rect 401 2538 418 2543
rect 140 2509 156 2538
rect 190 2509 216 2538
rect 258 2509 274 2538
rect 308 2509 334 2538
rect 400 2509 418 2538
rect 452 2538 459 2543
rect 493 2538 522 2572
rect 1246 2542 1280 2558
rect 452 2509 468 2538
rect 1246 2466 1280 2482
rect 1334 2545 1368 2561
rect 1334 2469 1368 2485
rect 1978 2545 2012 2561
rect 1978 2469 2012 2485
rect 2083 2545 2117 2561
rect 2083 2469 2117 2485
rect 2192 2545 2226 2561
rect 2192 2469 2226 2485
rect 3190 2545 3224 2561
rect 3190 2469 3224 2485
rect 3294 2545 3328 2561
rect 3294 2469 3328 2485
rect 3404 2545 3438 2561
rect 3404 2469 3438 2485
rect 4402 2545 4436 2561
rect 4402 2469 4436 2485
rect 4507 2545 4541 2561
rect 4507 2469 4541 2485
rect 4616 2545 4650 2561
rect 4616 2469 4650 2485
rect 5614 2545 5648 2561
rect 5614 2469 5648 2485
rect 5721 2545 5755 2561
rect 5721 2469 5755 2485
rect 5828 2545 5862 2561
rect 5828 2469 5862 2485
rect 6389 2548 6423 2564
rect 6389 2472 6423 2488
rect 6477 2548 6511 2564
rect 6477 2472 6511 2488
rect 6573 2548 6607 2564
rect 6573 2472 6607 2488
rect 6669 2548 6703 2564
rect 6771 2538 6800 2572
rect 6834 2543 6892 2572
rect 6926 2543 6984 2572
rect 6834 2538 6865 2543
rect 6926 2538 6983 2543
rect 7018 2538 7076 2572
rect 7110 2543 7168 2572
rect 7110 2538 7127 2543
rect 6849 2509 6865 2538
rect 6899 2509 6925 2538
rect 6967 2509 6983 2538
rect 7017 2509 7043 2538
rect 7109 2509 7127 2538
rect 7161 2538 7168 2543
rect 7202 2538 7231 2572
rect 7955 2542 7989 2558
rect 7161 2509 7177 2538
rect 6669 2472 6703 2488
rect 7955 2466 7989 2482
rect 8043 2545 8077 2561
rect 8043 2469 8077 2485
rect 8687 2545 8721 2561
rect 8687 2469 8721 2485
rect 8792 2545 8826 2561
rect 8792 2469 8826 2485
rect 8901 2545 8935 2561
rect 8901 2469 8935 2485
rect 9899 2545 9933 2561
rect 9899 2469 9933 2485
rect 10003 2545 10037 2561
rect 10003 2469 10037 2485
rect 10113 2545 10147 2561
rect 10113 2469 10147 2485
rect 11111 2545 11145 2561
rect 11111 2469 11145 2485
rect 11216 2545 11250 2561
rect 11216 2469 11250 2485
rect 11325 2545 11359 2561
rect 11325 2469 11359 2485
rect 12323 2545 12357 2561
rect 12323 2469 12357 2485
rect 12430 2545 12464 2561
rect 12430 2469 12464 2485
rect 12537 2545 12571 2561
rect 12537 2469 12571 2485
rect 13098 2548 13132 2564
rect 13098 2472 13132 2488
rect 13186 2548 13220 2564
rect 13186 2472 13220 2488
rect 13282 2548 13316 2564
rect 13282 2472 13316 2488
rect 13378 2548 13412 2564
rect 13378 2472 13412 2488
rect 6302 2397 6318 2431
rect 6352 2397 6368 2431
rect 6509 2395 6525 2429
rect 6559 2395 6575 2429
rect 13011 2397 13027 2431
rect 13061 2397 13077 2431
rect 13218 2395 13234 2429
rect 13268 2395 13284 2429
rect 1599 2344 1633 2360
rect 1599 2268 1633 2284
rect 1689 2344 1723 2360
rect 1689 2268 1723 2284
rect 2331 2344 2365 2360
rect 2331 2268 2365 2284
rect 2438 2344 2472 2360
rect 2438 2268 2472 2284
rect 2541 2344 2575 2360
rect 2541 2268 2575 2284
rect 3543 2344 3577 2360
rect 3543 2268 3577 2284
rect 3649 2344 3683 2360
rect 3649 2268 3683 2284
rect 3753 2344 3787 2360
rect 3753 2268 3787 2284
rect 4881 2344 4915 2360
rect 4881 2268 4915 2284
rect 4989 2344 5023 2360
rect 4989 2268 5023 2284
rect 5091 2344 5125 2360
rect 5091 2268 5125 2284
rect 5736 2344 5770 2360
rect 5736 2268 5770 2284
rect 5825 2344 5859 2360
rect 5825 2268 5859 2284
rect 6389 2345 6423 2361
rect 6389 2269 6423 2285
rect 6477 2345 6511 2361
rect 6477 2269 6511 2285
rect 6573 2345 6607 2361
rect 6573 2269 6607 2285
rect 6669 2345 6703 2361
rect 6669 2269 6703 2285
rect 8308 2344 8342 2360
rect 8308 2268 8342 2284
rect 8398 2344 8432 2360
rect 8398 2268 8432 2284
rect 9040 2344 9074 2360
rect 9040 2268 9074 2284
rect 9147 2344 9181 2360
rect 9147 2268 9181 2284
rect 9250 2344 9284 2360
rect 9250 2268 9284 2284
rect 10252 2344 10286 2360
rect 10252 2268 10286 2284
rect 10358 2344 10392 2360
rect 10358 2268 10392 2284
rect 10462 2344 10496 2360
rect 10462 2268 10496 2284
rect 11590 2344 11624 2360
rect 11590 2268 11624 2284
rect 11698 2344 11732 2360
rect 11698 2268 11732 2284
rect 11800 2344 11834 2360
rect 11800 2268 11834 2284
rect 12445 2344 12479 2360
rect 12445 2268 12479 2284
rect 12534 2344 12568 2360
rect 12534 2268 12568 2284
rect 13098 2345 13132 2361
rect 13098 2269 13132 2285
rect 13186 2345 13220 2361
rect 13186 2269 13220 2285
rect 13282 2345 13316 2361
rect 13282 2269 13316 2285
rect 13378 2345 13412 2361
rect 13378 2269 13412 2285
rect 643 2210 659 2244
rect 693 2210 709 2244
rect 1627 2200 1643 2234
rect 1677 2200 1693 2234
rect 2359 2200 2375 2234
rect 2409 2200 2425 2234
rect 2481 2200 2497 2234
rect 2531 2200 2547 2234
rect 3571 2200 3587 2234
rect 3621 2200 3637 2234
rect 3693 2200 3709 2234
rect 3743 2200 3759 2234
rect 4909 2200 4925 2234
rect 4959 2200 4975 2234
rect 5031 2200 5047 2234
rect 5081 2200 5097 2234
rect 5765 2200 5781 2234
rect 5815 2200 5831 2234
rect 6389 2207 6423 2223
rect 579 2160 613 2176
rect 579 2084 613 2100
rect 739 2160 773 2176
rect 6389 2131 6423 2147
rect 6477 2207 6511 2223
rect 7352 2210 7368 2244
rect 7402 2210 7418 2244
rect 8336 2200 8352 2234
rect 8386 2200 8402 2234
rect 9068 2200 9084 2234
rect 9118 2200 9134 2234
rect 9190 2200 9206 2234
rect 9240 2200 9256 2234
rect 10280 2200 10296 2234
rect 10330 2200 10346 2234
rect 10402 2200 10418 2234
rect 10452 2200 10468 2234
rect 11618 2200 11634 2234
rect 11668 2200 11684 2234
rect 11740 2200 11756 2234
rect 11790 2200 11806 2234
rect 12474 2200 12490 2234
rect 12524 2200 12540 2234
rect 13098 2207 13132 2223
rect 6477 2131 6511 2147
rect 7288 2160 7322 2176
rect 739 2084 773 2100
rect 7288 2084 7322 2100
rect 7448 2160 7482 2176
rect 13098 2131 13132 2147
rect 13186 2207 13220 2223
rect 13186 2131 13220 2147
rect 7448 2084 7482 2100
rect 579 2022 613 2038
rect 579 1946 613 1962
rect 739 2022 773 2038
rect 739 1946 773 1962
rect 7288 2022 7322 2038
rect 7288 1946 7322 1962
rect 7448 2022 7482 2038
rect 7448 1946 7482 1962
rect 579 1884 613 1900
rect 579 1808 613 1824
rect 739 1884 773 1900
rect 739 1808 773 1824
rect 7288 1884 7322 1900
rect 7288 1808 7322 1824
rect 7448 1884 7482 1900
rect 7448 1808 7482 1824
rect 579 1746 613 1762
rect 77 1702 195 1721
rect 77 1645 103 1702
rect 169 1645 195 1702
rect 579 1670 613 1686
rect 739 1746 773 1762
rect 739 1670 773 1686
rect 7288 1746 7322 1762
rect 7288 1670 7322 1686
rect 7448 1746 7482 1762
rect 7448 1670 7482 1686
rect 77 1622 195 1645
rect 579 1608 613 1624
rect 579 1532 613 1548
rect 739 1608 773 1624
rect 739 1532 773 1548
rect 7288 1608 7322 1624
rect 7288 1532 7322 1548
rect 7448 1608 7482 1624
rect 7448 1532 7482 1548
rect 579 1470 613 1486
rect 579 1394 613 1410
rect 739 1470 773 1486
rect 739 1394 773 1410
rect 7288 1470 7322 1486
rect 7288 1394 7322 1410
rect 7448 1470 7482 1486
rect 7448 1394 7482 1410
rect 579 1332 613 1348
rect 579 1256 613 1272
rect 739 1332 773 1348
rect 739 1256 773 1272
rect 855 1318 960 1353
rect 855 1284 887 1318
rect 921 1284 960 1318
rect 855 1255 960 1284
rect 7288 1332 7322 1348
rect 7288 1256 7322 1272
rect 7448 1332 7482 1348
rect 7448 1256 7482 1272
rect 7564 1318 7669 1353
rect 7564 1284 7596 1318
rect 7630 1284 7669 1318
rect 7564 1255 7669 1284
rect 579 1194 613 1210
rect 579 1118 613 1134
rect 739 1200 773 1210
rect 869 1200 946 1255
rect 739 1194 946 1200
rect 773 1134 946 1194
rect 7288 1194 7322 1210
rect 739 1131 946 1134
rect 1254 1147 1586 1163
rect 739 1118 773 1131
rect 1254 1113 1280 1147
rect 1314 1113 1360 1147
rect 1394 1113 1440 1147
rect 1474 1113 1520 1147
rect 1554 1113 1586 1147
rect 1254 1095 1586 1113
rect 1986 1147 2318 1163
rect 1986 1113 2012 1147
rect 2046 1113 2092 1147
rect 2126 1113 2172 1147
rect 2206 1113 2252 1147
rect 2286 1113 2318 1147
rect 1986 1095 2318 1113
rect 2588 1147 2920 1163
rect 2588 1113 2620 1147
rect 2654 1113 2700 1147
rect 2734 1113 2780 1147
rect 2814 1113 2860 1147
rect 2894 1113 2920 1147
rect 2588 1095 2920 1113
rect 3198 1147 3530 1163
rect 3198 1113 3224 1147
rect 3258 1113 3304 1147
rect 3338 1113 3384 1147
rect 3418 1113 3464 1147
rect 3498 1113 3530 1147
rect 3198 1095 3530 1113
rect 3800 1147 4132 1163
rect 3800 1113 3832 1147
rect 3866 1113 3912 1147
rect 3946 1113 3992 1147
rect 4026 1113 4072 1147
rect 4106 1113 4132 1147
rect 3800 1095 4132 1113
rect 4536 1147 4868 1163
rect 4536 1113 4562 1147
rect 4596 1113 4642 1147
rect 4676 1113 4722 1147
rect 4756 1113 4802 1147
rect 4836 1113 4868 1147
rect 4536 1095 4868 1113
rect 5138 1147 5470 1163
rect 5138 1113 5170 1147
rect 5204 1113 5250 1147
rect 5284 1113 5330 1147
rect 5364 1113 5410 1147
rect 5444 1113 5470 1147
rect 5138 1095 5470 1113
rect 5872 1147 6204 1163
rect 5872 1113 5904 1147
rect 5938 1113 5984 1147
rect 6018 1113 6064 1147
rect 6098 1113 6144 1147
rect 6178 1113 6204 1147
rect 7288 1118 7322 1134
rect 7448 1200 7482 1210
rect 7578 1200 7655 1255
rect 7448 1194 7655 1200
rect 7482 1134 7655 1194
rect 7448 1131 7655 1134
rect 7963 1147 8295 1163
rect 7448 1118 7482 1131
rect 5872 1095 6204 1113
rect 7963 1113 7989 1147
rect 8023 1113 8069 1147
rect 8103 1113 8149 1147
rect 8183 1113 8229 1147
rect 8263 1113 8295 1147
rect 7963 1095 8295 1113
rect 8695 1147 9027 1163
rect 8695 1113 8721 1147
rect 8755 1113 8801 1147
rect 8835 1113 8881 1147
rect 8915 1113 8961 1147
rect 8995 1113 9027 1147
rect 8695 1095 9027 1113
rect 9297 1147 9629 1163
rect 9297 1113 9329 1147
rect 9363 1113 9409 1147
rect 9443 1113 9489 1147
rect 9523 1113 9569 1147
rect 9603 1113 9629 1147
rect 9297 1095 9629 1113
rect 9907 1147 10239 1163
rect 9907 1113 9933 1147
rect 9967 1113 10013 1147
rect 10047 1113 10093 1147
rect 10127 1113 10173 1147
rect 10207 1113 10239 1147
rect 9907 1095 10239 1113
rect 10509 1147 10841 1163
rect 10509 1113 10541 1147
rect 10575 1113 10621 1147
rect 10655 1113 10701 1147
rect 10735 1113 10781 1147
rect 10815 1113 10841 1147
rect 10509 1095 10841 1113
rect 11245 1147 11577 1163
rect 11245 1113 11271 1147
rect 11305 1113 11351 1147
rect 11385 1113 11431 1147
rect 11465 1113 11511 1147
rect 11545 1113 11577 1147
rect 11245 1095 11577 1113
rect 11847 1147 12179 1163
rect 11847 1113 11879 1147
rect 11913 1113 11959 1147
rect 11993 1113 12039 1147
rect 12073 1113 12119 1147
rect 12153 1113 12179 1147
rect 11847 1095 12179 1113
rect 12581 1147 12913 1163
rect 12581 1113 12613 1147
rect 12647 1113 12693 1147
rect 12727 1113 12773 1147
rect 12807 1113 12853 1147
rect 12887 1113 12913 1147
rect 12581 1095 12913 1113
rect 551 208 883 226
rect 551 174 577 208
rect 611 174 657 208
rect 691 174 737 208
rect 771 174 817 208
rect 851 174 883 208
rect 551 158 883 174
rect 1285 208 1617 226
rect 1285 174 1311 208
rect 1345 174 1391 208
rect 1425 174 1471 208
rect 1505 174 1551 208
rect 1585 174 1617 208
rect 1285 158 1617 174
rect 1887 208 2219 226
rect 1887 174 1919 208
rect 1953 174 1999 208
rect 2033 174 2079 208
rect 2113 174 2159 208
rect 2193 174 2219 208
rect 1887 158 2219 174
rect 2623 208 2955 226
rect 2623 174 2649 208
rect 2683 174 2729 208
rect 2763 174 2809 208
rect 2843 174 2889 208
rect 2923 174 2955 208
rect 2623 158 2955 174
rect 3225 208 3557 226
rect 3225 174 3257 208
rect 3291 174 3337 208
rect 3371 174 3417 208
rect 3451 174 3497 208
rect 3531 174 3557 208
rect 3225 158 3557 174
rect 3835 208 4167 226
rect 3835 174 3861 208
rect 3895 174 3941 208
rect 3975 174 4021 208
rect 4055 174 4101 208
rect 4135 174 4167 208
rect 3835 158 4167 174
rect 4437 208 4769 226
rect 4437 174 4469 208
rect 4503 174 4549 208
rect 4583 174 4629 208
rect 4663 174 4709 208
rect 4743 174 4769 208
rect 4437 158 4769 174
rect 5169 208 5501 226
rect 5169 174 5201 208
rect 5235 174 5281 208
rect 5315 174 5361 208
rect 5395 174 5441 208
rect 5475 174 5501 208
rect 7260 208 7592 226
rect 5982 190 6016 203
rect 5169 158 5501 174
rect 5809 187 6016 190
rect 5809 127 5982 187
rect 5809 121 6016 127
rect 5809 66 5886 121
rect 5982 111 6016 121
rect 6142 187 6176 203
rect 7260 174 7286 208
rect 7320 174 7366 208
rect 7400 174 7446 208
rect 7480 174 7526 208
rect 7560 174 7592 208
rect 7260 158 7592 174
rect 7994 208 8326 226
rect 7994 174 8020 208
rect 8054 174 8100 208
rect 8134 174 8180 208
rect 8214 174 8260 208
rect 8294 174 8326 208
rect 7994 158 8326 174
rect 8596 208 8928 226
rect 8596 174 8628 208
rect 8662 174 8708 208
rect 8742 174 8788 208
rect 8822 174 8868 208
rect 8902 174 8928 208
rect 8596 158 8928 174
rect 9332 208 9664 226
rect 9332 174 9358 208
rect 9392 174 9438 208
rect 9472 174 9518 208
rect 9552 174 9598 208
rect 9632 174 9664 208
rect 9332 158 9664 174
rect 9934 208 10266 226
rect 9934 174 9966 208
rect 10000 174 10046 208
rect 10080 174 10126 208
rect 10160 174 10206 208
rect 10240 174 10266 208
rect 9934 158 10266 174
rect 10544 208 10876 226
rect 10544 174 10570 208
rect 10604 174 10650 208
rect 10684 174 10730 208
rect 10764 174 10810 208
rect 10844 174 10876 208
rect 10544 158 10876 174
rect 11146 208 11478 226
rect 11146 174 11178 208
rect 11212 174 11258 208
rect 11292 174 11338 208
rect 11372 174 11418 208
rect 11452 174 11478 208
rect 11146 158 11478 174
rect 11878 208 12210 226
rect 11878 174 11910 208
rect 11944 174 11990 208
rect 12024 174 12070 208
rect 12104 174 12150 208
rect 12184 174 12210 208
rect 12691 190 12725 203
rect 11878 158 12210 174
rect 12518 187 12725 190
rect 6142 111 6176 127
rect 12518 127 12691 187
rect 12518 121 12725 127
rect 12518 66 12595 121
rect 12691 111 12725 121
rect 12851 187 12885 203
rect 12851 111 12885 127
rect 5795 37 5900 66
rect 5795 3 5834 37
rect 5868 3 5900 37
rect 5795 -32 5900 3
rect 5982 49 6016 65
rect 5982 -27 6016 -11
rect 6142 49 6176 65
rect 6142 -27 6176 -11
rect 12504 37 12609 66
rect 12504 3 12543 37
rect 12577 3 12609 37
rect 12504 -32 12609 3
rect 12691 49 12725 65
rect 12691 -27 12725 -11
rect 12851 49 12885 65
rect 12851 -27 12885 -11
rect 5982 -89 6016 -73
rect 5982 -165 6016 -149
rect 6142 -89 6176 -73
rect 6142 -165 6176 -149
rect 12691 -89 12725 -73
rect 12691 -165 12725 -149
rect 12851 -89 12885 -73
rect 12851 -165 12885 -149
rect 5982 -227 6016 -211
rect 5982 -303 6016 -287
rect 6142 -227 6176 -211
rect 6142 -303 6176 -287
rect 12691 -227 12725 -211
rect 12691 -303 12725 -287
rect 12851 -227 12885 -211
rect 12851 -303 12885 -287
rect 5982 -365 6016 -349
rect 5982 -441 6016 -425
rect 6142 -365 6176 -349
rect 6142 -441 6176 -425
rect 12691 -365 12725 -349
rect 12691 -441 12725 -425
rect 12851 -365 12885 -349
rect 12851 -441 12885 -425
rect 5982 -503 6016 -487
rect 5982 -579 6016 -563
rect 6142 -503 6176 -487
rect 6142 -579 6176 -563
rect 12691 -503 12725 -487
rect 12691 -579 12725 -563
rect 12851 -503 12885 -487
rect 12851 -579 12885 -563
rect 5982 -641 6016 -625
rect 5982 -717 6016 -701
rect 6142 -641 6176 -625
rect 6142 -717 6176 -701
rect 12691 -641 12725 -625
rect 12691 -717 12725 -701
rect 12851 -641 12885 -625
rect 12851 -717 12885 -701
rect 5982 -779 6016 -763
rect 244 -826 278 -810
rect 244 -902 278 -886
rect 332 -826 366 -810
rect 5982 -855 6016 -839
rect 6142 -779 6176 -763
rect 12691 -779 12725 -763
rect 6142 -855 6176 -839
rect 6953 -826 6987 -810
rect 332 -902 366 -886
rect 924 -913 940 -879
rect 974 -913 990 -879
rect 1658 -913 1674 -879
rect 1708 -913 1724 -879
rect 1780 -913 1796 -879
rect 1830 -913 1846 -879
rect 2996 -913 3012 -879
rect 3046 -913 3062 -879
rect 3118 -913 3134 -879
rect 3168 -913 3184 -879
rect 4208 -913 4224 -879
rect 4258 -913 4274 -879
rect 4330 -913 4346 -879
rect 4380 -913 4396 -879
rect 5062 -913 5078 -879
rect 5112 -913 5128 -879
rect 6046 -923 6062 -889
rect 6096 -923 6112 -889
rect 6953 -902 6987 -886
rect 7041 -826 7075 -810
rect 12691 -855 12725 -839
rect 12851 -779 12885 -763
rect 12851 -855 12885 -839
rect 7041 -902 7075 -886
rect 7633 -913 7649 -879
rect 7683 -913 7699 -879
rect 8367 -913 8383 -879
rect 8417 -913 8433 -879
rect 8489 -913 8505 -879
rect 8539 -913 8555 -879
rect 9705 -913 9721 -879
rect 9755 -913 9771 -879
rect 9827 -913 9843 -879
rect 9877 -913 9893 -879
rect 10917 -913 10933 -879
rect 10967 -913 10983 -879
rect 11039 -913 11055 -879
rect 11089 -913 11105 -879
rect 11771 -913 11787 -879
rect 11821 -913 11837 -879
rect 12755 -923 12771 -889
rect 12805 -923 12821 -889
rect 52 -964 86 -948
rect 52 -1040 86 -1024
rect 148 -964 182 -948
rect 148 -1040 182 -1024
rect 244 -964 278 -948
rect 244 -1040 278 -1024
rect 332 -964 366 -948
rect 332 -1040 366 -1024
rect 896 -963 930 -947
rect 896 -1039 930 -1023
rect 985 -963 1019 -947
rect 985 -1039 1019 -1023
rect 1630 -963 1664 -947
rect 1630 -1039 1664 -1023
rect 1732 -963 1766 -947
rect 1732 -1039 1766 -1023
rect 1840 -963 1874 -947
rect 1840 -1039 1874 -1023
rect 2968 -963 3002 -947
rect 2968 -1039 3002 -1023
rect 3072 -963 3106 -947
rect 3072 -1039 3106 -1023
rect 3178 -963 3212 -947
rect 3178 -1039 3212 -1023
rect 4180 -963 4214 -947
rect 4180 -1039 4214 -1023
rect 4283 -963 4317 -947
rect 4283 -1039 4317 -1023
rect 4390 -963 4424 -947
rect 4390 -1039 4424 -1023
rect 5032 -963 5066 -947
rect 5032 -1039 5066 -1023
rect 5122 -963 5156 -947
rect 5122 -1039 5156 -1023
rect 6761 -964 6795 -948
rect 6761 -1040 6795 -1024
rect 6857 -964 6891 -948
rect 6857 -1040 6891 -1024
rect 6953 -964 6987 -948
rect 6953 -1040 6987 -1024
rect 7041 -964 7075 -948
rect 7041 -1040 7075 -1024
rect 7605 -963 7639 -947
rect 7605 -1039 7639 -1023
rect 7694 -963 7728 -947
rect 7694 -1039 7728 -1023
rect 8339 -963 8373 -947
rect 8339 -1039 8373 -1023
rect 8441 -963 8475 -947
rect 8441 -1039 8475 -1023
rect 8549 -963 8583 -947
rect 8549 -1039 8583 -1023
rect 9677 -963 9711 -947
rect 9677 -1039 9711 -1023
rect 9781 -963 9815 -947
rect 9781 -1039 9815 -1023
rect 9887 -963 9921 -947
rect 9887 -1039 9921 -1023
rect 10889 -963 10923 -947
rect 10889 -1039 10923 -1023
rect 10992 -963 11026 -947
rect 10992 -1039 11026 -1023
rect 11099 -963 11133 -947
rect 11099 -1039 11133 -1023
rect 11741 -963 11775 -947
rect 11741 -1039 11775 -1023
rect 11831 -963 11865 -947
rect 11831 -1039 11865 -1023
rect 180 -1108 196 -1074
rect 230 -1108 246 -1074
rect 387 -1110 403 -1076
rect 437 -1110 453 -1076
rect 6889 -1108 6905 -1074
rect 6939 -1108 6955 -1074
rect 7096 -1110 7112 -1076
rect 7146 -1110 7162 -1076
rect 52 -1167 86 -1151
rect 52 -1243 86 -1227
rect 148 -1167 182 -1151
rect 148 -1243 182 -1227
rect 244 -1167 278 -1151
rect 244 -1243 278 -1227
rect 332 -1167 366 -1151
rect 332 -1243 366 -1227
rect 893 -1164 927 -1148
rect 893 -1240 927 -1224
rect 1000 -1164 1034 -1148
rect 1000 -1240 1034 -1224
rect 1107 -1164 1141 -1148
rect 1107 -1240 1141 -1224
rect 2105 -1164 2139 -1148
rect 2105 -1240 2139 -1224
rect 2214 -1164 2248 -1148
rect 2214 -1240 2248 -1224
rect 2319 -1164 2353 -1148
rect 2319 -1240 2353 -1224
rect 3317 -1164 3351 -1148
rect 3317 -1240 3351 -1224
rect 3427 -1164 3461 -1148
rect 3427 -1240 3461 -1224
rect 3531 -1164 3565 -1148
rect 3531 -1240 3565 -1224
rect 4529 -1164 4563 -1148
rect 4529 -1240 4563 -1224
rect 4638 -1164 4672 -1148
rect 4638 -1240 4672 -1224
rect 4743 -1164 4777 -1148
rect 4743 -1240 4777 -1224
rect 5387 -1164 5421 -1148
rect 5387 -1240 5421 -1224
rect 5475 -1161 5509 -1145
rect 6761 -1167 6795 -1151
rect 6287 -1217 6303 -1188
rect 5475 -1237 5509 -1221
rect 6233 -1251 6262 -1217
rect 6296 -1222 6303 -1217
rect 6337 -1217 6355 -1188
rect 6421 -1217 6447 -1188
rect 6481 -1217 6497 -1188
rect 6539 -1217 6565 -1188
rect 6599 -1217 6615 -1188
rect 6337 -1222 6354 -1217
rect 6296 -1251 6354 -1222
rect 6388 -1251 6446 -1217
rect 6481 -1222 6538 -1217
rect 6599 -1222 6630 -1217
rect 6480 -1251 6538 -1222
rect 6572 -1251 6630 -1222
rect 6664 -1251 6693 -1217
rect 6761 -1243 6795 -1227
rect 6857 -1167 6891 -1151
rect 6857 -1243 6891 -1227
rect 6953 -1167 6987 -1151
rect 6953 -1243 6987 -1227
rect 7041 -1167 7075 -1151
rect 7041 -1243 7075 -1227
rect 7602 -1164 7636 -1148
rect 7602 -1240 7636 -1224
rect 7709 -1164 7743 -1148
rect 7709 -1240 7743 -1224
rect 7816 -1164 7850 -1148
rect 7816 -1240 7850 -1224
rect 8814 -1164 8848 -1148
rect 8814 -1240 8848 -1224
rect 8923 -1164 8957 -1148
rect 8923 -1240 8957 -1224
rect 9028 -1164 9062 -1148
rect 9028 -1240 9062 -1224
rect 10026 -1164 10060 -1148
rect 10026 -1240 10060 -1224
rect 10136 -1164 10170 -1148
rect 10136 -1240 10170 -1224
rect 10240 -1164 10274 -1148
rect 10240 -1240 10274 -1224
rect 11238 -1164 11272 -1148
rect 11238 -1240 11272 -1224
rect 11347 -1164 11381 -1148
rect 11347 -1240 11381 -1224
rect 11452 -1164 11486 -1148
rect 11452 -1240 11486 -1224
rect 12096 -1164 12130 -1148
rect 12096 -1240 12130 -1224
rect 12184 -1161 12218 -1145
rect 12996 -1217 13012 -1188
rect 12184 -1237 12218 -1221
rect 12942 -1251 12971 -1217
rect 13005 -1222 13012 -1217
rect 13046 -1217 13064 -1188
rect 13130 -1217 13156 -1188
rect 13190 -1217 13206 -1188
rect 13248 -1217 13274 -1188
rect 13308 -1217 13324 -1188
rect 13046 -1222 13063 -1217
rect 13005 -1251 13063 -1222
rect 13097 -1251 13155 -1217
rect 13190 -1222 13247 -1217
rect 13308 -1222 13339 -1217
rect 13189 -1251 13247 -1222
rect 13281 -1251 13339 -1222
rect 13373 -1251 13402 -1217
rect 244 -1305 278 -1289
rect 244 -1381 278 -1365
rect 332 -1305 366 -1289
rect 921 -1317 937 -1283
rect 971 -1317 987 -1283
rect 1047 -1317 1063 -1283
rect 1097 -1317 1113 -1283
rect 2133 -1317 2149 -1283
rect 2183 -1317 2199 -1283
rect 2259 -1317 2275 -1283
rect 2309 -1317 2325 -1283
rect 3345 -1317 3361 -1283
rect 3395 -1317 3411 -1283
rect 3471 -1317 3487 -1283
rect 3521 -1317 3537 -1283
rect 4557 -1317 4573 -1283
rect 4607 -1317 4623 -1283
rect 4683 -1317 4699 -1283
rect 4733 -1317 4749 -1283
rect 5415 -1314 5431 -1280
rect 5465 -1314 5481 -1280
rect 5866 -1284 5915 -1272
rect 5866 -1285 6006 -1284
rect 5866 -1319 5872 -1285
rect 5906 -1318 6006 -1285
rect 5906 -1319 5915 -1318
rect 5866 -1331 5915 -1319
rect 5965 -1360 6006 -1318
rect 6297 -1297 6343 -1251
rect 6297 -1331 6309 -1297
rect 6126 -1360 6175 -1347
rect 332 -1381 366 -1365
rect 5867 -1378 5916 -1365
rect 5867 -1412 5873 -1378
rect 5907 -1412 5916 -1378
rect 5965 -1394 6132 -1360
rect 6166 -1394 6175 -1360
rect 6126 -1406 6175 -1394
rect 6297 -1365 6343 -1331
rect 6297 -1399 6309 -1365
rect 5867 -1424 5916 -1412
rect 6297 -1415 6343 -1399
rect 6377 -1297 6443 -1285
rect 6377 -1331 6393 -1297
rect 6427 -1331 6443 -1297
rect 6377 -1365 6443 -1331
rect 6377 -1399 6393 -1365
rect 6427 -1399 6443 -1365
rect 6377 -1411 6443 -1399
rect 5881 -1447 5916 -1424
rect 6164 -1447 6213 -1440
rect 5881 -1453 6213 -1447
rect 5881 -1482 6170 -1453
rect 6164 -1487 6170 -1482
rect 6204 -1487 6213 -1453
rect 6164 -1499 6213 -1487
rect 6297 -1452 6313 -1449
rect 6297 -1486 6309 -1452
rect 6347 -1483 6363 -1449
rect 6343 -1486 6363 -1483
rect 6297 -1497 6363 -1486
rect 6057 -1557 6073 -1523
rect 6107 -1557 6123 -1523
rect 6397 -1531 6443 -1411
rect 6301 -1549 6343 -1533
rect 6301 -1583 6309 -1549
rect 6029 -1616 6063 -1600
rect 126 -1685 212 -1659
rect 126 -1719 152 -1685
rect 186 -1719 212 -1685
rect 6029 -1692 6063 -1676
rect 6117 -1616 6151 -1600
rect 6117 -1692 6151 -1676
rect 6301 -1617 6343 -1583
rect 6301 -1651 6309 -1617
rect 6301 -1685 6343 -1651
rect 126 -1745 212 -1719
rect 6301 -1719 6309 -1685
rect 6029 -1754 6063 -1738
rect 125 -1842 211 -1816
rect 6029 -1830 6063 -1814
rect 6117 -1754 6151 -1738
rect 6301 -1761 6343 -1719
rect 6377 -1549 6443 -1531
rect 6377 -1597 6393 -1549
rect 6427 -1597 6443 -1549
rect 6377 -1617 6443 -1597
rect 6377 -1651 6393 -1617
rect 6427 -1651 6443 -1617
rect 6377 -1685 6443 -1651
rect 6377 -1719 6393 -1685
rect 6427 -1719 6443 -1685
rect 6377 -1727 6443 -1719
rect 6483 -1297 6549 -1285
rect 6483 -1331 6499 -1297
rect 6533 -1331 6549 -1297
rect 6483 -1365 6549 -1331
rect 6483 -1399 6499 -1365
rect 6533 -1399 6549 -1365
rect 6483 -1411 6549 -1399
rect 6583 -1297 6629 -1251
rect 6617 -1331 6629 -1297
rect 6583 -1365 6629 -1331
rect 6617 -1399 6629 -1365
rect 6953 -1305 6987 -1289
rect 6953 -1381 6987 -1365
rect 7041 -1305 7075 -1289
rect 7630 -1317 7646 -1283
rect 7680 -1317 7696 -1283
rect 7756 -1317 7772 -1283
rect 7806 -1317 7822 -1283
rect 8842 -1317 8858 -1283
rect 8892 -1317 8908 -1283
rect 8968 -1317 8984 -1283
rect 9018 -1317 9034 -1283
rect 10054 -1317 10070 -1283
rect 10104 -1317 10120 -1283
rect 10180 -1317 10196 -1283
rect 10230 -1317 10246 -1283
rect 11266 -1317 11282 -1283
rect 11316 -1317 11332 -1283
rect 11392 -1317 11408 -1283
rect 11442 -1317 11458 -1283
rect 12124 -1314 12140 -1280
rect 12174 -1314 12190 -1280
rect 12575 -1284 12624 -1272
rect 12575 -1285 12715 -1284
rect 12575 -1319 12581 -1285
rect 12615 -1318 12715 -1285
rect 12615 -1319 12624 -1318
rect 12575 -1331 12624 -1319
rect 12674 -1360 12715 -1318
rect 13006 -1297 13052 -1251
rect 13006 -1331 13018 -1297
rect 12835 -1360 12884 -1347
rect 7041 -1381 7075 -1365
rect 12576 -1378 12625 -1365
rect 6483 -1531 6529 -1411
rect 6583 -1415 6629 -1399
rect 12576 -1412 12582 -1378
rect 12616 -1412 12625 -1378
rect 12674 -1394 12841 -1360
rect 12875 -1394 12884 -1360
rect 12835 -1406 12884 -1394
rect 13006 -1365 13052 -1331
rect 13006 -1399 13018 -1365
rect 12576 -1424 12625 -1412
rect 13006 -1415 13052 -1399
rect 13086 -1297 13152 -1285
rect 13086 -1331 13102 -1297
rect 13136 -1331 13152 -1297
rect 13086 -1365 13152 -1331
rect 13086 -1399 13102 -1365
rect 13136 -1399 13152 -1365
rect 13086 -1411 13152 -1399
rect 12590 -1447 12625 -1424
rect 12873 -1447 12922 -1440
rect 6563 -1483 6579 -1449
rect 6613 -1453 6629 -1449
rect 6563 -1487 6583 -1483
rect 6617 -1487 6629 -1453
rect 12590 -1453 12922 -1447
rect 12590 -1482 12879 -1453
rect 6563 -1497 6629 -1487
rect 12873 -1487 12879 -1482
rect 12913 -1487 12922 -1453
rect 12873 -1499 12922 -1487
rect 13006 -1452 13022 -1449
rect 13006 -1486 13018 -1452
rect 13056 -1483 13072 -1449
rect 13052 -1486 13072 -1483
rect 13006 -1497 13072 -1486
rect 6483 -1549 6549 -1531
rect 6483 -1583 6499 -1549
rect 6533 -1583 6549 -1549
rect 6483 -1617 6549 -1583
rect 6483 -1651 6499 -1617
rect 6533 -1618 6549 -1617
rect 6483 -1652 6502 -1651
rect 6536 -1652 6549 -1618
rect 6483 -1685 6549 -1652
rect 6483 -1719 6499 -1685
rect 6533 -1719 6549 -1685
rect 6483 -1727 6549 -1719
rect 6583 -1549 6625 -1533
rect 6617 -1583 6625 -1549
rect 12766 -1557 12782 -1523
rect 12816 -1557 12832 -1523
rect 13106 -1531 13152 -1411
rect 13010 -1549 13052 -1533
rect 6583 -1617 6625 -1583
rect 13010 -1583 13018 -1549
rect 6617 -1651 6625 -1617
rect 6583 -1685 6625 -1651
rect 12738 -1616 12772 -1600
rect 6617 -1719 6625 -1685
rect 6583 -1761 6625 -1719
rect 6835 -1685 6921 -1659
rect 6835 -1719 6861 -1685
rect 6895 -1719 6921 -1685
rect 12738 -1692 12772 -1676
rect 12826 -1616 12860 -1600
rect 12826 -1692 12860 -1676
rect 13010 -1617 13052 -1583
rect 13010 -1651 13018 -1617
rect 13010 -1685 13052 -1651
rect 6835 -1745 6921 -1719
rect 13010 -1719 13018 -1685
rect 12738 -1754 12772 -1738
rect 6233 -1795 6262 -1761
rect 6296 -1790 6354 -1761
rect 6296 -1795 6309 -1790
rect 6117 -1830 6151 -1814
rect 6289 -1824 6309 -1795
rect 6343 -1795 6354 -1790
rect 6388 -1795 6446 -1761
rect 6480 -1790 6538 -1761
rect 6489 -1795 6538 -1790
rect 6572 -1790 6630 -1761
rect 6572 -1795 6585 -1790
rect 6343 -1824 6359 -1795
rect 6435 -1824 6455 -1795
rect 6489 -1824 6505 -1795
rect 6569 -1824 6585 -1795
rect 6619 -1795 6630 -1790
rect 6664 -1795 6693 -1761
rect 6619 -1824 6635 -1795
rect 125 -1876 151 -1842
rect 185 -1876 211 -1842
rect 6834 -1842 6920 -1816
rect 12738 -1830 12772 -1814
rect 12826 -1754 12860 -1738
rect 13010 -1761 13052 -1719
rect 13086 -1549 13152 -1531
rect 13086 -1597 13102 -1549
rect 13136 -1597 13152 -1549
rect 13086 -1617 13152 -1597
rect 13086 -1651 13102 -1617
rect 13136 -1651 13152 -1617
rect 13086 -1685 13152 -1651
rect 13086 -1719 13102 -1685
rect 13136 -1719 13152 -1685
rect 13086 -1727 13152 -1719
rect 13192 -1297 13258 -1285
rect 13192 -1331 13208 -1297
rect 13242 -1331 13258 -1297
rect 13192 -1365 13258 -1331
rect 13192 -1399 13208 -1365
rect 13242 -1399 13258 -1365
rect 13192 -1411 13258 -1399
rect 13292 -1297 13338 -1251
rect 13326 -1331 13338 -1297
rect 13292 -1365 13338 -1331
rect 13326 -1399 13338 -1365
rect 13192 -1531 13238 -1411
rect 13292 -1415 13338 -1399
rect 13272 -1483 13288 -1449
rect 13322 -1453 13338 -1449
rect 13272 -1487 13292 -1483
rect 13326 -1487 13338 -1453
rect 13272 -1497 13338 -1487
rect 13192 -1549 13258 -1531
rect 13192 -1583 13208 -1549
rect 13242 -1583 13258 -1549
rect 13192 -1617 13258 -1583
rect 13192 -1651 13208 -1617
rect 13242 -1618 13258 -1617
rect 13192 -1652 13211 -1651
rect 13245 -1652 13258 -1618
rect 13192 -1685 13258 -1652
rect 13192 -1719 13208 -1685
rect 13242 -1719 13258 -1685
rect 13192 -1727 13258 -1719
rect 13292 -1549 13334 -1533
rect 13326 -1583 13334 -1549
rect 13292 -1617 13334 -1583
rect 13326 -1651 13334 -1617
rect 13292 -1685 13334 -1651
rect 13326 -1719 13334 -1685
rect 13292 -1761 13334 -1719
rect 12942 -1795 12971 -1761
rect 13005 -1790 13063 -1761
rect 13005 -1795 13018 -1790
rect 12826 -1830 12860 -1814
rect 12998 -1824 13018 -1795
rect 13052 -1795 13063 -1790
rect 13097 -1795 13155 -1761
rect 13189 -1790 13247 -1761
rect 13198 -1795 13247 -1790
rect 13281 -1790 13339 -1761
rect 13281 -1795 13294 -1790
rect 13052 -1824 13068 -1795
rect 13144 -1824 13164 -1795
rect 13198 -1824 13214 -1795
rect 13278 -1824 13294 -1795
rect 13328 -1795 13339 -1790
rect 13373 -1795 13402 -1761
rect 13328 -1824 13344 -1795
rect 6834 -1876 6860 -1842
rect 6894 -1876 6920 -1842
rect 125 -1902 211 -1876
rect 6029 -1892 6063 -1876
rect 6029 -1968 6063 -1952
rect 6117 -1892 6151 -1876
rect 6117 -1968 6151 -1952
rect 6412 -1914 6498 -1888
rect 6834 -1902 6920 -1876
rect 12738 -1892 12772 -1876
rect 6412 -1948 6438 -1914
rect 6472 -1948 6498 -1914
rect 6412 -1974 6498 -1948
rect 12738 -1968 12772 -1952
rect 12826 -1892 12860 -1876
rect 12826 -1968 12860 -1952
rect 125 -2012 211 -1986
rect 125 -2046 151 -2012
rect 185 -2046 211 -2012
rect 6834 -2012 6920 -1986
rect 125 -2072 211 -2046
rect 6029 -2030 6063 -2014
rect 6029 -2106 6063 -2090
rect 6117 -2030 6151 -2014
rect 6834 -2046 6860 -2012
rect 6894 -2046 6920 -2012
rect 6834 -2072 6920 -2046
rect 12738 -2030 12772 -2014
rect 6117 -2106 6151 -2090
rect 6412 -2110 6498 -2084
rect 12738 -2106 12772 -2090
rect 12826 -2030 12860 -2014
rect 12826 -2106 12860 -2090
rect 126 -2164 212 -2138
rect 6412 -2144 6438 -2110
rect 6472 -2144 6498 -2110
rect 126 -2198 152 -2164
rect 186 -2198 212 -2164
rect 126 -2224 212 -2198
rect 5880 -2177 5963 -2153
rect 5880 -2212 5904 -2177
rect 5938 -2212 5963 -2177
rect 5880 -2237 5963 -2212
rect 6029 -2168 6063 -2152
rect 131 -2308 217 -2282
rect 131 -2342 157 -2308
rect 191 -2342 217 -2308
rect 5893 -2301 5950 -2237
rect 6029 -2244 6063 -2228
rect 6117 -2168 6151 -2152
rect 6412 -2170 6498 -2144
rect 6835 -2164 6921 -2138
rect 6835 -2198 6861 -2164
rect 6895 -2198 6921 -2164
rect 6835 -2224 6921 -2198
rect 12589 -2177 12672 -2153
rect 12589 -2212 12613 -2177
rect 12647 -2212 12672 -2177
rect 6117 -2244 6151 -2228
rect 12589 -2237 12672 -2212
rect 12738 -2168 12772 -2152
rect 6412 -2285 6498 -2259
rect 6029 -2301 6063 -2290
rect 5893 -2306 6063 -2301
rect 5893 -2342 6029 -2306
rect 131 -2368 217 -2342
rect 381 -2359 5289 -2345
rect 381 -2393 497 -2359
rect 533 -2393 577 -2359
rect 613 -2393 657 -2359
rect 693 -2393 737 -2359
rect 773 -2393 817 -2359
rect 853 -2393 897 -2359
rect 933 -2393 1101 -2359
rect 1137 -2393 1181 -2359
rect 1217 -2393 1261 -2359
rect 1297 -2393 1341 -2359
rect 1377 -2393 1421 -2359
rect 1457 -2393 1501 -2359
rect 1537 -2393 1709 -2359
rect 1745 -2393 1789 -2359
rect 1825 -2393 1869 -2359
rect 1905 -2393 1949 -2359
rect 1985 -2393 2029 -2359
rect 2065 -2393 2109 -2359
rect 2145 -2393 2313 -2359
rect 2349 -2393 2393 -2359
rect 2429 -2393 2473 -2359
rect 2509 -2393 2553 -2359
rect 2589 -2393 2633 -2359
rect 2669 -2393 2713 -2359
rect 2749 -2393 2921 -2359
rect 2957 -2393 3001 -2359
rect 3037 -2393 3081 -2359
rect 3117 -2393 3161 -2359
rect 3197 -2393 3241 -2359
rect 3277 -2393 3321 -2359
rect 3357 -2393 3525 -2359
rect 3561 -2393 3605 -2359
rect 3641 -2393 3685 -2359
rect 3721 -2393 3765 -2359
rect 3801 -2393 3845 -2359
rect 3881 -2393 3925 -2359
rect 3961 -2393 4133 -2359
rect 4169 -2393 4213 -2359
rect 4249 -2393 4293 -2359
rect 4329 -2393 4373 -2359
rect 4409 -2393 4453 -2359
rect 4489 -2393 4533 -2359
rect 4569 -2393 4737 -2359
rect 4773 -2393 4817 -2359
rect 4853 -2393 4897 -2359
rect 4933 -2393 4977 -2359
rect 5013 -2393 5057 -2359
rect 5093 -2393 5137 -2359
rect 5173 -2393 5289 -2359
rect 381 -2411 5289 -2393
rect 5351 -2356 6029 -2342
rect 5351 -2390 5469 -2356
rect 5505 -2390 5549 -2356
rect 5585 -2390 5629 -2356
rect 5665 -2390 5709 -2356
rect 5745 -2390 5789 -2356
rect 5825 -2390 5869 -2356
rect 5905 -2366 6029 -2356
rect 5905 -2382 6063 -2366
rect 6117 -2306 6151 -2290
rect 6412 -2319 6438 -2285
rect 6472 -2319 6498 -2285
rect 6412 -2345 6498 -2319
rect 6840 -2308 6926 -2282
rect 6840 -2342 6866 -2308
rect 6900 -2342 6926 -2308
rect 12602 -2301 12659 -2237
rect 12738 -2244 12772 -2228
rect 12826 -2168 12860 -2152
rect 12826 -2244 12860 -2228
rect 12738 -2301 12772 -2290
rect 12602 -2306 12772 -2301
rect 12602 -2342 12738 -2306
rect 6117 -2382 6151 -2366
rect 6840 -2368 6926 -2342
rect 7090 -2359 11998 -2345
rect 5905 -2390 6021 -2382
rect 5351 -2408 6021 -2390
rect 7090 -2393 7206 -2359
rect 7242 -2393 7286 -2359
rect 7322 -2393 7366 -2359
rect 7402 -2393 7446 -2359
rect 7482 -2393 7526 -2359
rect 7562 -2393 7606 -2359
rect 7642 -2393 7810 -2359
rect 7846 -2393 7890 -2359
rect 7926 -2393 7970 -2359
rect 8006 -2393 8050 -2359
rect 8086 -2393 8130 -2359
rect 8166 -2393 8210 -2359
rect 8246 -2393 8418 -2359
rect 8454 -2393 8498 -2359
rect 8534 -2393 8578 -2359
rect 8614 -2393 8658 -2359
rect 8694 -2393 8738 -2359
rect 8774 -2393 8818 -2359
rect 8854 -2393 9022 -2359
rect 9058 -2393 9102 -2359
rect 9138 -2393 9182 -2359
rect 9218 -2393 9262 -2359
rect 9298 -2393 9342 -2359
rect 9378 -2393 9422 -2359
rect 9458 -2393 9630 -2359
rect 9666 -2393 9710 -2359
rect 9746 -2393 9790 -2359
rect 9826 -2393 9870 -2359
rect 9906 -2393 9950 -2359
rect 9986 -2393 10030 -2359
rect 10066 -2393 10234 -2359
rect 10270 -2393 10314 -2359
rect 10350 -2393 10394 -2359
rect 10430 -2393 10474 -2359
rect 10510 -2393 10554 -2359
rect 10590 -2393 10634 -2359
rect 10670 -2393 10842 -2359
rect 10878 -2393 10922 -2359
rect 10958 -2393 11002 -2359
rect 11038 -2393 11082 -2359
rect 11118 -2393 11162 -2359
rect 11198 -2393 11242 -2359
rect 11278 -2393 11446 -2359
rect 11482 -2393 11526 -2359
rect 11562 -2393 11606 -2359
rect 11642 -2393 11686 -2359
rect 11722 -2393 11766 -2359
rect 11802 -2393 11846 -2359
rect 11882 -2393 11998 -2359
rect 7090 -2411 11998 -2393
rect 12060 -2356 12738 -2342
rect 12060 -2390 12178 -2356
rect 12214 -2390 12258 -2356
rect 12294 -2390 12338 -2356
rect 12374 -2390 12418 -2356
rect 12454 -2390 12498 -2356
rect 12534 -2390 12578 -2356
rect 12614 -2366 12738 -2356
rect 12614 -2382 12772 -2366
rect 12826 -2306 12860 -2290
rect 12826 -2382 12860 -2366
rect 12614 -2390 12730 -2382
rect 12060 -2408 12730 -2390
<< viali >>
rect 604 3627 638 3687
rect 692 3627 726 3687
rect 852 3677 884 3711
rect 884 3677 886 3711
rect 932 3677 964 3711
rect 964 3677 966 3711
rect 1012 3677 1044 3711
rect 1044 3677 1046 3711
rect 1092 3677 1124 3711
rect 1124 3677 1126 3711
rect 1172 3677 1204 3711
rect 1204 3677 1206 3711
rect 1252 3677 1284 3711
rect 1284 3677 1286 3711
rect 1584 3680 1616 3714
rect 1616 3680 1618 3714
rect 1664 3680 1696 3714
rect 1696 3680 1698 3714
rect 1744 3680 1776 3714
rect 1776 3680 1778 3714
rect 1824 3680 1856 3714
rect 1856 3680 1858 3714
rect 1904 3680 1936 3714
rect 1936 3680 1938 3714
rect 1984 3680 2016 3714
rect 2016 3680 2018 3714
rect 2186 3680 2188 3714
rect 2188 3680 2220 3714
rect 2266 3680 2268 3714
rect 2268 3680 2300 3714
rect 2346 3680 2348 3714
rect 2348 3680 2380 3714
rect 2426 3680 2428 3714
rect 2428 3680 2460 3714
rect 2506 3680 2508 3714
rect 2508 3680 2540 3714
rect 2586 3680 2588 3714
rect 2588 3680 2620 3714
rect 2796 3680 2828 3714
rect 2828 3680 2830 3714
rect 2876 3680 2908 3714
rect 2908 3680 2910 3714
rect 2956 3680 2988 3714
rect 2988 3680 2990 3714
rect 3036 3680 3068 3714
rect 3068 3680 3070 3714
rect 3116 3680 3148 3714
rect 3148 3680 3150 3714
rect 3196 3680 3228 3714
rect 3228 3680 3230 3714
rect 3398 3680 3400 3714
rect 3400 3680 3432 3714
rect 3478 3680 3480 3714
rect 3480 3680 3512 3714
rect 3558 3680 3560 3714
rect 3560 3680 3592 3714
rect 3638 3680 3640 3714
rect 3640 3680 3672 3714
rect 3718 3680 3720 3714
rect 3720 3680 3752 3714
rect 3798 3680 3800 3714
rect 3800 3680 3832 3714
rect 4008 3680 4040 3714
rect 4040 3680 4042 3714
rect 4088 3680 4120 3714
rect 4120 3680 4122 3714
rect 4168 3680 4200 3714
rect 4200 3680 4202 3714
rect 4248 3680 4280 3714
rect 4280 3680 4282 3714
rect 4328 3680 4360 3714
rect 4360 3680 4362 3714
rect 4408 3680 4440 3714
rect 4440 3680 4442 3714
rect 4610 3680 4612 3714
rect 4612 3680 4644 3714
rect 4690 3680 4692 3714
rect 4692 3680 4724 3714
rect 4770 3680 4772 3714
rect 4772 3680 4804 3714
rect 4850 3680 4852 3714
rect 4852 3680 4884 3714
rect 4930 3680 4932 3714
rect 4932 3680 4964 3714
rect 5010 3680 5012 3714
rect 5012 3680 5044 3714
rect 5220 3680 5252 3714
rect 5252 3680 5254 3714
rect 5300 3680 5332 3714
rect 5332 3680 5334 3714
rect 5380 3680 5412 3714
rect 5412 3680 5414 3714
rect 5460 3680 5492 3714
rect 5492 3680 5494 3714
rect 5540 3680 5572 3714
rect 5572 3680 5574 3714
rect 5620 3680 5652 3714
rect 5652 3680 5654 3714
rect 5822 3680 5824 3714
rect 5824 3680 5856 3714
rect 5902 3680 5904 3714
rect 5904 3680 5936 3714
rect 5982 3680 5984 3714
rect 5984 3680 6016 3714
rect 6062 3680 6064 3714
rect 6064 3680 6096 3714
rect 6142 3680 6144 3714
rect 6144 3680 6176 3714
rect 6222 3680 6224 3714
rect 6224 3680 6256 3714
rect 604 3489 638 3549
rect 6564 3629 6598 3663
rect 7041 3632 7075 3666
rect 7313 3627 7347 3687
rect 7401 3627 7435 3687
rect 7561 3677 7593 3711
rect 7593 3677 7595 3711
rect 7641 3677 7673 3711
rect 7673 3677 7675 3711
rect 7721 3677 7753 3711
rect 7753 3677 7755 3711
rect 7801 3677 7833 3711
rect 7833 3677 7835 3711
rect 7881 3677 7913 3711
rect 7913 3677 7915 3711
rect 7961 3677 7993 3711
rect 7993 3677 7995 3711
rect 8293 3680 8325 3714
rect 8325 3680 8327 3714
rect 8373 3680 8405 3714
rect 8405 3680 8407 3714
rect 8453 3680 8485 3714
rect 8485 3680 8487 3714
rect 8533 3680 8565 3714
rect 8565 3680 8567 3714
rect 8613 3680 8645 3714
rect 8645 3680 8647 3714
rect 8693 3680 8725 3714
rect 8725 3680 8727 3714
rect 8895 3680 8897 3714
rect 8897 3680 8929 3714
rect 8975 3680 8977 3714
rect 8977 3680 9009 3714
rect 9055 3680 9057 3714
rect 9057 3680 9089 3714
rect 9135 3680 9137 3714
rect 9137 3680 9169 3714
rect 9215 3680 9217 3714
rect 9217 3680 9249 3714
rect 9295 3680 9297 3714
rect 9297 3680 9329 3714
rect 9505 3680 9537 3714
rect 9537 3680 9539 3714
rect 9585 3680 9617 3714
rect 9617 3680 9619 3714
rect 9665 3680 9697 3714
rect 9697 3680 9699 3714
rect 9745 3680 9777 3714
rect 9777 3680 9779 3714
rect 9825 3680 9857 3714
rect 9857 3680 9859 3714
rect 9905 3680 9937 3714
rect 9937 3680 9939 3714
rect 10107 3680 10109 3714
rect 10109 3680 10141 3714
rect 10187 3680 10189 3714
rect 10189 3680 10221 3714
rect 10267 3680 10269 3714
rect 10269 3680 10301 3714
rect 10347 3680 10349 3714
rect 10349 3680 10381 3714
rect 10427 3680 10429 3714
rect 10429 3680 10461 3714
rect 10507 3680 10509 3714
rect 10509 3680 10541 3714
rect 10717 3680 10749 3714
rect 10749 3680 10751 3714
rect 10797 3680 10829 3714
rect 10829 3680 10831 3714
rect 10877 3680 10909 3714
rect 10909 3680 10911 3714
rect 10957 3680 10989 3714
rect 10989 3680 10991 3714
rect 11037 3680 11069 3714
rect 11069 3680 11071 3714
rect 11117 3680 11149 3714
rect 11149 3680 11151 3714
rect 11319 3680 11321 3714
rect 11321 3680 11353 3714
rect 11399 3680 11401 3714
rect 11401 3680 11433 3714
rect 11479 3680 11481 3714
rect 11481 3680 11513 3714
rect 11559 3680 11561 3714
rect 11561 3680 11593 3714
rect 11639 3680 11641 3714
rect 11641 3680 11673 3714
rect 11719 3680 11721 3714
rect 11721 3680 11753 3714
rect 11929 3680 11961 3714
rect 11961 3680 11963 3714
rect 12009 3680 12041 3714
rect 12041 3680 12043 3714
rect 12089 3680 12121 3714
rect 12121 3680 12123 3714
rect 12169 3680 12201 3714
rect 12201 3680 12203 3714
rect 12249 3680 12281 3714
rect 12281 3680 12283 3714
rect 12329 3680 12361 3714
rect 12361 3680 12363 3714
rect 12531 3680 12533 3714
rect 12533 3680 12565 3714
rect 12611 3680 12613 3714
rect 12613 3680 12645 3714
rect 12691 3680 12693 3714
rect 12693 3680 12725 3714
rect 12771 3680 12773 3714
rect 12773 3680 12805 3714
rect 12851 3680 12853 3714
rect 12853 3680 12885 3714
rect 12931 3680 12933 3714
rect 12933 3680 12965 3714
rect 692 3489 726 3549
rect 6569 3485 6603 3519
rect 7030 3460 7064 3494
rect 7313 3489 7347 3549
rect 13273 3629 13307 3663
rect 7401 3489 7435 3549
rect 13278 3485 13312 3519
rect 604 3351 638 3411
rect 692 3351 726 3411
rect 6570 3333 6604 3367
rect 7313 3351 7347 3411
rect 7401 3351 7435 3411
rect 13279 3333 13313 3367
rect 604 3213 638 3273
rect 692 3213 726 3273
rect 7030 3268 7064 3302
rect 7313 3213 7347 3273
rect 7401 3213 7435 3273
rect 6570 3163 6604 3197
rect 91 3082 125 3116
rect 183 3082 217 3116
rect 275 3111 300 3116
rect 300 3111 309 3116
rect 275 3082 309 3111
rect 367 3082 401 3116
rect 459 3082 493 3116
rect 219 2972 253 2973
rect 219 2939 222 2972
rect 222 2939 253 2972
rect 138 2804 172 2808
rect 138 2774 142 2804
rect 142 2774 172 2804
rect 328 2904 362 2918
rect 328 2884 362 2904
rect 604 3075 638 3135
rect 13279 3163 13313 3197
rect 692 3075 726 3135
rect 6800 3082 6834 3116
rect 6892 3082 6926 3116
rect 6984 3111 7009 3116
rect 7009 3111 7018 3116
rect 6984 3082 7018 3111
rect 7076 3082 7110 3116
rect 7168 3082 7202 3116
rect 604 2937 638 2997
rect 692 2937 726 2997
rect 6569 3006 6603 3040
rect 648 2844 682 2878
rect 6928 2972 6962 2973
rect 6928 2939 6931 2972
rect 6931 2939 6962 2972
rect 412 2804 446 2807
rect 412 2773 442 2804
rect 442 2773 446 2804
rect 551 2774 585 2808
rect 6847 2804 6881 2808
rect 6847 2774 6851 2804
rect 6851 2774 6881 2804
rect 589 2681 623 2715
rect 848 2699 882 2733
rect 849 2606 883 2640
rect 1290 2601 1324 2635
rect 2022 2604 2056 2638
rect 2148 2604 2182 2638
rect 3234 2604 3268 2638
rect 3360 2604 3394 2638
rect 4446 2604 4480 2638
rect 4572 2604 4606 2638
rect 5658 2604 5692 2638
rect 5784 2604 5818 2638
rect 6389 2626 6423 2686
rect 6477 2626 6511 2686
rect 7037 2904 7071 2918
rect 7037 2884 7071 2904
rect 7313 3075 7347 3135
rect 7401 3075 7435 3135
rect 7313 2937 7347 2997
rect 7401 2937 7435 2997
rect 13278 3006 13312 3040
rect 7357 2844 7391 2878
rect 7121 2804 7155 2807
rect 7121 2773 7151 2804
rect 7151 2773 7155 2804
rect 7260 2774 7294 2808
rect 7298 2681 7332 2715
rect 7557 2699 7591 2733
rect 7558 2606 7592 2640
rect 7999 2601 8033 2635
rect 8731 2604 8765 2638
rect 8857 2604 8891 2638
rect 9943 2604 9977 2638
rect 10069 2604 10103 2638
rect 11155 2604 11189 2638
rect 11281 2604 11315 2638
rect 12367 2604 12401 2638
rect 12493 2604 12527 2638
rect 13098 2626 13132 2686
rect 13186 2626 13220 2686
rect 91 2538 125 2572
rect 183 2543 217 2572
rect 275 2543 309 2572
rect 183 2538 190 2543
rect 190 2538 217 2543
rect 275 2538 308 2543
rect 308 2538 309 2543
rect 367 2538 401 2572
rect 459 2538 493 2572
rect 1246 2482 1280 2542
rect 1334 2485 1368 2545
rect 1978 2485 2012 2545
rect 2083 2485 2117 2545
rect 2192 2485 2226 2545
rect 3190 2485 3224 2545
rect 3294 2485 3328 2545
rect 3404 2485 3438 2545
rect 4402 2485 4436 2545
rect 4507 2485 4541 2545
rect 4616 2485 4650 2545
rect 5614 2485 5648 2545
rect 5721 2485 5755 2545
rect 5828 2485 5862 2545
rect 6389 2488 6423 2548
rect 6477 2488 6511 2548
rect 6573 2488 6607 2548
rect 6669 2488 6703 2548
rect 6800 2538 6834 2572
rect 6892 2543 6926 2572
rect 6984 2543 7018 2572
rect 6892 2538 6899 2543
rect 6899 2538 6926 2543
rect 6984 2538 7017 2543
rect 7017 2538 7018 2543
rect 7076 2538 7110 2572
rect 7168 2538 7202 2572
rect 7955 2482 7989 2542
rect 8043 2485 8077 2545
rect 8687 2485 8721 2545
rect 8792 2485 8826 2545
rect 8901 2485 8935 2545
rect 9899 2485 9933 2545
rect 10003 2485 10037 2545
rect 10113 2485 10147 2545
rect 11111 2485 11145 2545
rect 11216 2485 11250 2545
rect 11325 2485 11359 2545
rect 12323 2485 12357 2545
rect 12430 2485 12464 2545
rect 12537 2485 12571 2545
rect 13098 2488 13132 2548
rect 13186 2488 13220 2548
rect 13282 2488 13316 2548
rect 13378 2488 13412 2548
rect 6318 2397 6352 2431
rect 6525 2395 6559 2429
rect 13027 2397 13061 2431
rect 13234 2395 13268 2429
rect 1599 2284 1633 2344
rect 1689 2284 1723 2344
rect 2331 2284 2365 2344
rect 2438 2284 2472 2344
rect 2541 2284 2575 2344
rect 3543 2284 3577 2344
rect 3649 2284 3683 2344
rect 3753 2284 3787 2344
rect 4881 2284 4915 2344
rect 4989 2284 5023 2344
rect 5091 2284 5125 2344
rect 5736 2284 5770 2344
rect 5825 2284 5859 2344
rect 6389 2285 6423 2345
rect 6477 2285 6511 2345
rect 6573 2285 6607 2345
rect 6669 2285 6703 2345
rect 8308 2284 8342 2344
rect 8398 2284 8432 2344
rect 9040 2284 9074 2344
rect 9147 2284 9181 2344
rect 9250 2284 9284 2344
rect 10252 2284 10286 2344
rect 10358 2284 10392 2344
rect 10462 2284 10496 2344
rect 11590 2284 11624 2344
rect 11698 2284 11732 2344
rect 11800 2284 11834 2344
rect 12445 2284 12479 2344
rect 12534 2284 12568 2344
rect 13098 2285 13132 2345
rect 13186 2285 13220 2345
rect 13282 2285 13316 2345
rect 13378 2285 13412 2345
rect 659 2210 693 2244
rect 1643 2200 1677 2234
rect 2375 2200 2409 2234
rect 2497 2200 2531 2234
rect 3587 2200 3621 2234
rect 3709 2200 3743 2234
rect 4925 2200 4959 2234
rect 5047 2200 5081 2234
rect 5781 2200 5815 2234
rect 579 2100 613 2160
rect 739 2100 773 2160
rect 6389 2147 6423 2207
rect 7368 2210 7402 2244
rect 6477 2147 6511 2207
rect 8352 2200 8386 2234
rect 9084 2200 9118 2234
rect 9206 2200 9240 2234
rect 10296 2200 10330 2234
rect 10418 2200 10452 2234
rect 11634 2200 11668 2234
rect 11756 2200 11790 2234
rect 12490 2200 12524 2234
rect 7288 2100 7322 2160
rect 7448 2100 7482 2160
rect 13098 2147 13132 2207
rect 13186 2147 13220 2207
rect 579 1962 613 2022
rect 739 1962 773 2022
rect 7288 1962 7322 2022
rect 7448 1962 7482 2022
rect 579 1824 613 1884
rect 739 1824 773 1884
rect 7288 1824 7322 1884
rect 7448 1824 7482 1884
rect 105 1649 163 1700
rect 579 1686 613 1746
rect 739 1686 773 1746
rect 7288 1686 7322 1746
rect 7448 1686 7482 1746
rect 579 1548 613 1608
rect 739 1548 773 1608
rect 7288 1548 7322 1608
rect 7448 1548 7482 1608
rect 579 1410 613 1470
rect 739 1410 773 1470
rect 7288 1410 7322 1470
rect 7448 1410 7482 1470
rect 579 1272 613 1332
rect 739 1272 773 1332
rect 7288 1272 7322 1332
rect 7448 1272 7482 1332
rect 579 1134 613 1194
rect 739 1134 773 1194
rect 1280 1113 1314 1147
rect 1360 1113 1394 1147
rect 1440 1113 1474 1147
rect 1520 1113 1554 1147
rect 2012 1113 2046 1147
rect 2092 1113 2126 1147
rect 2172 1113 2206 1147
rect 2252 1113 2286 1147
rect 2620 1113 2654 1147
rect 2700 1113 2734 1147
rect 2780 1113 2814 1147
rect 2860 1113 2894 1147
rect 3224 1113 3258 1147
rect 3304 1113 3338 1147
rect 3384 1113 3418 1147
rect 3464 1113 3498 1147
rect 3832 1113 3866 1147
rect 3912 1113 3946 1147
rect 3992 1113 4026 1147
rect 4072 1113 4106 1147
rect 4562 1113 4596 1147
rect 4642 1113 4676 1147
rect 4722 1113 4756 1147
rect 4802 1113 4836 1147
rect 5170 1113 5204 1147
rect 5250 1113 5284 1147
rect 5330 1113 5364 1147
rect 5410 1113 5444 1147
rect 5904 1113 5938 1147
rect 5984 1113 6018 1147
rect 6064 1113 6098 1147
rect 6144 1113 6178 1147
rect 7288 1134 7322 1194
rect 7448 1134 7482 1194
rect 7989 1113 8023 1147
rect 8069 1113 8103 1147
rect 8149 1113 8183 1147
rect 8229 1113 8263 1147
rect 8721 1113 8755 1147
rect 8801 1113 8835 1147
rect 8881 1113 8915 1147
rect 8961 1113 8995 1147
rect 9329 1113 9363 1147
rect 9409 1113 9443 1147
rect 9489 1113 9523 1147
rect 9569 1113 9603 1147
rect 9933 1113 9967 1147
rect 10013 1113 10047 1147
rect 10093 1113 10127 1147
rect 10173 1113 10207 1147
rect 10541 1113 10575 1147
rect 10621 1113 10655 1147
rect 10701 1113 10735 1147
rect 10781 1113 10815 1147
rect 11271 1113 11305 1147
rect 11351 1113 11385 1147
rect 11431 1113 11465 1147
rect 11511 1113 11545 1147
rect 11879 1113 11913 1147
rect 11959 1113 11993 1147
rect 12039 1113 12073 1147
rect 12119 1113 12153 1147
rect 12613 1113 12647 1147
rect 12693 1113 12727 1147
rect 12773 1113 12807 1147
rect 12853 1113 12887 1147
rect 577 174 611 208
rect 657 174 691 208
rect 737 174 771 208
rect 817 174 851 208
rect 1311 174 1345 208
rect 1391 174 1425 208
rect 1471 174 1505 208
rect 1551 174 1585 208
rect 1919 174 1953 208
rect 1999 174 2033 208
rect 2079 174 2113 208
rect 2159 174 2193 208
rect 2649 174 2683 208
rect 2729 174 2763 208
rect 2809 174 2843 208
rect 2889 174 2923 208
rect 3257 174 3291 208
rect 3337 174 3371 208
rect 3417 174 3451 208
rect 3497 174 3531 208
rect 3861 174 3895 208
rect 3941 174 3975 208
rect 4021 174 4055 208
rect 4101 174 4135 208
rect 4469 174 4503 208
rect 4549 174 4583 208
rect 4629 174 4663 208
rect 4709 174 4743 208
rect 5201 174 5235 208
rect 5281 174 5315 208
rect 5361 174 5395 208
rect 5441 174 5475 208
rect 5982 127 6016 187
rect 6142 127 6176 187
rect 7286 174 7320 208
rect 7366 174 7400 208
rect 7446 174 7480 208
rect 7526 174 7560 208
rect 8020 174 8054 208
rect 8100 174 8134 208
rect 8180 174 8214 208
rect 8260 174 8294 208
rect 8628 174 8662 208
rect 8708 174 8742 208
rect 8788 174 8822 208
rect 8868 174 8902 208
rect 9358 174 9392 208
rect 9438 174 9472 208
rect 9518 174 9552 208
rect 9598 174 9632 208
rect 9966 174 10000 208
rect 10046 174 10080 208
rect 10126 174 10160 208
rect 10206 174 10240 208
rect 10570 174 10604 208
rect 10650 174 10684 208
rect 10730 174 10764 208
rect 10810 174 10844 208
rect 11178 174 11212 208
rect 11258 174 11292 208
rect 11338 174 11372 208
rect 11418 174 11452 208
rect 11910 174 11944 208
rect 11990 174 12024 208
rect 12070 174 12104 208
rect 12150 174 12184 208
rect 12691 127 12725 187
rect 12851 127 12885 187
rect 5982 -11 6016 49
rect 6142 -11 6176 49
rect 12691 -11 12725 49
rect 12851 -11 12885 49
rect 5982 -149 6016 -89
rect 6142 -149 6176 -89
rect 12691 -149 12725 -89
rect 12851 -149 12885 -89
rect 5982 -287 6016 -227
rect 6142 -287 6176 -227
rect 12691 -287 12725 -227
rect 12851 -287 12885 -227
rect 5982 -425 6016 -365
rect 6142 -425 6176 -365
rect 12691 -425 12725 -365
rect 12851 -425 12885 -365
rect 5982 -563 6016 -503
rect 6142 -563 6176 -503
rect 12691 -563 12725 -503
rect 12851 -563 12885 -503
rect 5982 -701 6016 -641
rect 6142 -701 6176 -641
rect 12691 -701 12725 -641
rect 12851 -701 12885 -641
rect 244 -886 278 -826
rect 332 -886 366 -826
rect 5982 -839 6016 -779
rect 6142 -839 6176 -779
rect 940 -913 974 -879
rect 1674 -913 1708 -879
rect 1796 -913 1830 -879
rect 3012 -913 3046 -879
rect 3134 -913 3168 -879
rect 4224 -913 4258 -879
rect 4346 -913 4380 -879
rect 5078 -913 5112 -879
rect 6953 -886 6987 -826
rect 6062 -923 6096 -889
rect 7041 -886 7075 -826
rect 12691 -839 12725 -779
rect 12851 -839 12885 -779
rect 7649 -913 7683 -879
rect 8383 -913 8417 -879
rect 8505 -913 8539 -879
rect 9721 -913 9755 -879
rect 9843 -913 9877 -879
rect 10933 -913 10967 -879
rect 11055 -913 11089 -879
rect 11787 -913 11821 -879
rect 12771 -923 12805 -889
rect 52 -1024 86 -964
rect 148 -1024 182 -964
rect 244 -1024 278 -964
rect 332 -1024 366 -964
rect 896 -1023 930 -963
rect 985 -1023 1019 -963
rect 1630 -1023 1664 -963
rect 1732 -1023 1766 -963
rect 1840 -1023 1874 -963
rect 2968 -1023 3002 -963
rect 3072 -1023 3106 -963
rect 3178 -1023 3212 -963
rect 4180 -1023 4214 -963
rect 4283 -1023 4317 -963
rect 4390 -1023 4424 -963
rect 5032 -1023 5066 -963
rect 5122 -1023 5156 -963
rect 6761 -1024 6795 -964
rect 6857 -1024 6891 -964
rect 6953 -1024 6987 -964
rect 7041 -1024 7075 -964
rect 7605 -1023 7639 -963
rect 7694 -1023 7728 -963
rect 8339 -1023 8373 -963
rect 8441 -1023 8475 -963
rect 8549 -1023 8583 -963
rect 9677 -1023 9711 -963
rect 9781 -1023 9815 -963
rect 9887 -1023 9921 -963
rect 10889 -1023 10923 -963
rect 10992 -1023 11026 -963
rect 11099 -1023 11133 -963
rect 11741 -1023 11775 -963
rect 11831 -1023 11865 -963
rect 196 -1108 230 -1074
rect 403 -1110 437 -1076
rect 6905 -1108 6939 -1074
rect 7112 -1110 7146 -1076
rect 52 -1227 86 -1167
rect 148 -1227 182 -1167
rect 244 -1227 278 -1167
rect 332 -1227 366 -1167
rect 893 -1224 927 -1164
rect 1000 -1224 1034 -1164
rect 1107 -1224 1141 -1164
rect 2105 -1224 2139 -1164
rect 2214 -1224 2248 -1164
rect 2319 -1224 2353 -1164
rect 3317 -1224 3351 -1164
rect 3427 -1224 3461 -1164
rect 3531 -1224 3565 -1164
rect 4529 -1224 4563 -1164
rect 4638 -1224 4672 -1164
rect 4743 -1224 4777 -1164
rect 5387 -1224 5421 -1164
rect 5475 -1221 5509 -1161
rect 6262 -1251 6296 -1217
rect 6354 -1251 6388 -1217
rect 6446 -1222 6447 -1217
rect 6447 -1222 6480 -1217
rect 6538 -1222 6565 -1217
rect 6565 -1222 6572 -1217
rect 6446 -1251 6480 -1222
rect 6538 -1251 6572 -1222
rect 6630 -1251 6664 -1217
rect 6761 -1227 6795 -1167
rect 6857 -1227 6891 -1167
rect 6953 -1227 6987 -1167
rect 7041 -1227 7075 -1167
rect 7602 -1224 7636 -1164
rect 7709 -1224 7743 -1164
rect 7816 -1224 7850 -1164
rect 8814 -1224 8848 -1164
rect 8923 -1224 8957 -1164
rect 9028 -1224 9062 -1164
rect 10026 -1224 10060 -1164
rect 10136 -1224 10170 -1164
rect 10240 -1224 10274 -1164
rect 11238 -1224 11272 -1164
rect 11347 -1224 11381 -1164
rect 11452 -1224 11486 -1164
rect 12096 -1224 12130 -1164
rect 12184 -1221 12218 -1161
rect 12971 -1251 13005 -1217
rect 13063 -1251 13097 -1217
rect 13155 -1222 13156 -1217
rect 13156 -1222 13189 -1217
rect 13247 -1222 13274 -1217
rect 13274 -1222 13281 -1217
rect 13155 -1251 13189 -1222
rect 13247 -1251 13281 -1222
rect 13339 -1251 13373 -1217
rect 244 -1365 278 -1305
rect 332 -1365 366 -1305
rect 937 -1317 971 -1283
rect 1063 -1317 1097 -1283
rect 2149 -1317 2183 -1283
rect 2275 -1317 2309 -1283
rect 3361 -1317 3395 -1283
rect 3487 -1317 3521 -1283
rect 4573 -1317 4607 -1283
rect 4699 -1317 4733 -1283
rect 5431 -1314 5465 -1280
rect 5872 -1319 5906 -1285
rect 5873 -1412 5907 -1378
rect 6132 -1394 6166 -1360
rect 6170 -1487 6204 -1453
rect 6309 -1483 6313 -1452
rect 6313 -1483 6343 -1452
rect 6309 -1486 6343 -1483
rect 6073 -1557 6107 -1523
rect 152 -1719 186 -1685
rect 6029 -1676 6063 -1616
rect 6117 -1676 6151 -1616
rect 6029 -1814 6063 -1754
rect 6117 -1814 6151 -1754
rect 6393 -1583 6427 -1563
rect 6393 -1597 6427 -1583
rect 6953 -1365 6987 -1305
rect 7041 -1365 7075 -1305
rect 7646 -1317 7680 -1283
rect 7772 -1317 7806 -1283
rect 8858 -1317 8892 -1283
rect 8984 -1317 9018 -1283
rect 10070 -1317 10104 -1283
rect 10196 -1317 10230 -1283
rect 11282 -1317 11316 -1283
rect 11408 -1317 11442 -1283
rect 12140 -1314 12174 -1280
rect 12581 -1319 12615 -1285
rect 12582 -1412 12616 -1378
rect 12841 -1394 12875 -1360
rect 6583 -1483 6613 -1453
rect 6613 -1483 6617 -1453
rect 6583 -1487 6617 -1483
rect 12879 -1487 12913 -1453
rect 13018 -1483 13022 -1452
rect 13022 -1483 13052 -1452
rect 13018 -1486 13052 -1483
rect 6502 -1651 6533 -1618
rect 6533 -1651 6536 -1618
rect 6502 -1652 6536 -1651
rect 12782 -1557 12816 -1523
rect 6861 -1719 6895 -1685
rect 12738 -1676 12772 -1616
rect 12826 -1676 12860 -1616
rect 6262 -1795 6296 -1761
rect 6354 -1795 6388 -1761
rect 6446 -1790 6480 -1761
rect 6446 -1795 6455 -1790
rect 6455 -1795 6480 -1790
rect 6538 -1795 6572 -1761
rect 6630 -1795 6664 -1761
rect 12738 -1814 12772 -1754
rect 151 -1876 185 -1842
rect 12826 -1814 12860 -1754
rect 13102 -1583 13136 -1563
rect 13102 -1597 13136 -1583
rect 13292 -1483 13322 -1453
rect 13322 -1483 13326 -1453
rect 13292 -1487 13326 -1483
rect 13211 -1651 13242 -1618
rect 13242 -1651 13245 -1618
rect 13211 -1652 13245 -1651
rect 12971 -1795 13005 -1761
rect 13063 -1795 13097 -1761
rect 13155 -1790 13189 -1761
rect 13155 -1795 13164 -1790
rect 13164 -1795 13189 -1790
rect 13247 -1795 13281 -1761
rect 13339 -1795 13373 -1761
rect 6860 -1876 6894 -1842
rect 6029 -1952 6063 -1892
rect 6117 -1952 6151 -1892
rect 6438 -1948 6472 -1914
rect 12738 -1952 12772 -1892
rect 12826 -1952 12860 -1892
rect 151 -2046 185 -2012
rect 6029 -2090 6063 -2030
rect 6117 -2090 6151 -2030
rect 6860 -2046 6894 -2012
rect 12738 -2090 12772 -2030
rect 12826 -2090 12860 -2030
rect 6438 -2144 6472 -2110
rect 152 -2198 186 -2164
rect 6029 -2228 6063 -2168
rect 157 -2342 191 -2308
rect 6117 -2228 6151 -2168
rect 6861 -2198 6895 -2164
rect 12738 -2228 12772 -2168
rect 499 -2393 531 -2359
rect 531 -2393 533 -2359
rect 579 -2393 611 -2359
rect 611 -2393 613 -2359
rect 659 -2393 691 -2359
rect 691 -2393 693 -2359
rect 739 -2393 771 -2359
rect 771 -2393 773 -2359
rect 819 -2393 851 -2359
rect 851 -2393 853 -2359
rect 899 -2393 931 -2359
rect 931 -2393 933 -2359
rect 1101 -2393 1103 -2359
rect 1103 -2393 1135 -2359
rect 1181 -2393 1183 -2359
rect 1183 -2393 1215 -2359
rect 1261 -2393 1263 -2359
rect 1263 -2393 1295 -2359
rect 1341 -2393 1343 -2359
rect 1343 -2393 1375 -2359
rect 1421 -2393 1423 -2359
rect 1423 -2393 1455 -2359
rect 1501 -2393 1503 -2359
rect 1503 -2393 1535 -2359
rect 1711 -2393 1743 -2359
rect 1743 -2393 1745 -2359
rect 1791 -2393 1823 -2359
rect 1823 -2393 1825 -2359
rect 1871 -2393 1903 -2359
rect 1903 -2393 1905 -2359
rect 1951 -2393 1983 -2359
rect 1983 -2393 1985 -2359
rect 2031 -2393 2063 -2359
rect 2063 -2393 2065 -2359
rect 2111 -2393 2143 -2359
rect 2143 -2393 2145 -2359
rect 2313 -2393 2315 -2359
rect 2315 -2393 2347 -2359
rect 2393 -2393 2395 -2359
rect 2395 -2393 2427 -2359
rect 2473 -2393 2475 -2359
rect 2475 -2393 2507 -2359
rect 2553 -2393 2555 -2359
rect 2555 -2393 2587 -2359
rect 2633 -2393 2635 -2359
rect 2635 -2393 2667 -2359
rect 2713 -2393 2715 -2359
rect 2715 -2393 2747 -2359
rect 2923 -2393 2955 -2359
rect 2955 -2393 2957 -2359
rect 3003 -2393 3035 -2359
rect 3035 -2393 3037 -2359
rect 3083 -2393 3115 -2359
rect 3115 -2393 3117 -2359
rect 3163 -2393 3195 -2359
rect 3195 -2393 3197 -2359
rect 3243 -2393 3275 -2359
rect 3275 -2393 3277 -2359
rect 3323 -2393 3355 -2359
rect 3355 -2393 3357 -2359
rect 3525 -2393 3527 -2359
rect 3527 -2393 3559 -2359
rect 3605 -2393 3607 -2359
rect 3607 -2393 3639 -2359
rect 3685 -2393 3687 -2359
rect 3687 -2393 3719 -2359
rect 3765 -2393 3767 -2359
rect 3767 -2393 3799 -2359
rect 3845 -2393 3847 -2359
rect 3847 -2393 3879 -2359
rect 3925 -2393 3927 -2359
rect 3927 -2393 3959 -2359
rect 4135 -2393 4167 -2359
rect 4167 -2393 4169 -2359
rect 4215 -2393 4247 -2359
rect 4247 -2393 4249 -2359
rect 4295 -2393 4327 -2359
rect 4327 -2393 4329 -2359
rect 4375 -2393 4407 -2359
rect 4407 -2393 4409 -2359
rect 4455 -2393 4487 -2359
rect 4487 -2393 4489 -2359
rect 4535 -2393 4567 -2359
rect 4567 -2393 4569 -2359
rect 4737 -2393 4739 -2359
rect 4739 -2393 4771 -2359
rect 4817 -2393 4819 -2359
rect 4819 -2393 4851 -2359
rect 4897 -2393 4899 -2359
rect 4899 -2393 4931 -2359
rect 4977 -2393 4979 -2359
rect 4979 -2393 5011 -2359
rect 5057 -2393 5059 -2359
rect 5059 -2393 5091 -2359
rect 5137 -2393 5139 -2359
rect 5139 -2393 5171 -2359
rect 5469 -2390 5471 -2356
rect 5471 -2390 5503 -2356
rect 5549 -2390 5551 -2356
rect 5551 -2390 5583 -2356
rect 5629 -2390 5631 -2356
rect 5631 -2390 5663 -2356
rect 5709 -2390 5711 -2356
rect 5711 -2390 5743 -2356
rect 5789 -2390 5791 -2356
rect 5791 -2390 5823 -2356
rect 5869 -2390 5871 -2356
rect 5871 -2390 5903 -2356
rect 6029 -2366 6063 -2306
rect 6117 -2366 6151 -2306
rect 6438 -2319 6472 -2285
rect 6866 -2342 6900 -2308
rect 12826 -2228 12860 -2168
rect 7208 -2393 7240 -2359
rect 7240 -2393 7242 -2359
rect 7288 -2393 7320 -2359
rect 7320 -2393 7322 -2359
rect 7368 -2393 7400 -2359
rect 7400 -2393 7402 -2359
rect 7448 -2393 7480 -2359
rect 7480 -2393 7482 -2359
rect 7528 -2393 7560 -2359
rect 7560 -2393 7562 -2359
rect 7608 -2393 7640 -2359
rect 7640 -2393 7642 -2359
rect 7810 -2393 7812 -2359
rect 7812 -2393 7844 -2359
rect 7890 -2393 7892 -2359
rect 7892 -2393 7924 -2359
rect 7970 -2393 7972 -2359
rect 7972 -2393 8004 -2359
rect 8050 -2393 8052 -2359
rect 8052 -2393 8084 -2359
rect 8130 -2393 8132 -2359
rect 8132 -2393 8164 -2359
rect 8210 -2393 8212 -2359
rect 8212 -2393 8244 -2359
rect 8420 -2393 8452 -2359
rect 8452 -2393 8454 -2359
rect 8500 -2393 8532 -2359
rect 8532 -2393 8534 -2359
rect 8580 -2393 8612 -2359
rect 8612 -2393 8614 -2359
rect 8660 -2393 8692 -2359
rect 8692 -2393 8694 -2359
rect 8740 -2393 8772 -2359
rect 8772 -2393 8774 -2359
rect 8820 -2393 8852 -2359
rect 8852 -2393 8854 -2359
rect 9022 -2393 9024 -2359
rect 9024 -2393 9056 -2359
rect 9102 -2393 9104 -2359
rect 9104 -2393 9136 -2359
rect 9182 -2393 9184 -2359
rect 9184 -2393 9216 -2359
rect 9262 -2393 9264 -2359
rect 9264 -2393 9296 -2359
rect 9342 -2393 9344 -2359
rect 9344 -2393 9376 -2359
rect 9422 -2393 9424 -2359
rect 9424 -2393 9456 -2359
rect 9632 -2393 9664 -2359
rect 9664 -2393 9666 -2359
rect 9712 -2393 9744 -2359
rect 9744 -2393 9746 -2359
rect 9792 -2393 9824 -2359
rect 9824 -2393 9826 -2359
rect 9872 -2393 9904 -2359
rect 9904 -2393 9906 -2359
rect 9952 -2393 9984 -2359
rect 9984 -2393 9986 -2359
rect 10032 -2393 10064 -2359
rect 10064 -2393 10066 -2359
rect 10234 -2393 10236 -2359
rect 10236 -2393 10268 -2359
rect 10314 -2393 10316 -2359
rect 10316 -2393 10348 -2359
rect 10394 -2393 10396 -2359
rect 10396 -2393 10428 -2359
rect 10474 -2393 10476 -2359
rect 10476 -2393 10508 -2359
rect 10554 -2393 10556 -2359
rect 10556 -2393 10588 -2359
rect 10634 -2393 10636 -2359
rect 10636 -2393 10668 -2359
rect 10844 -2393 10876 -2359
rect 10876 -2393 10878 -2359
rect 10924 -2393 10956 -2359
rect 10956 -2393 10958 -2359
rect 11004 -2393 11036 -2359
rect 11036 -2393 11038 -2359
rect 11084 -2393 11116 -2359
rect 11116 -2393 11118 -2359
rect 11164 -2393 11196 -2359
rect 11196 -2393 11198 -2359
rect 11244 -2393 11276 -2359
rect 11276 -2393 11278 -2359
rect 11446 -2393 11448 -2359
rect 11448 -2393 11480 -2359
rect 11526 -2393 11528 -2359
rect 11528 -2393 11560 -2359
rect 11606 -2393 11608 -2359
rect 11608 -2393 11640 -2359
rect 11686 -2393 11688 -2359
rect 11688 -2393 11720 -2359
rect 11766 -2393 11768 -2359
rect 11768 -2393 11800 -2359
rect 11846 -2393 11848 -2359
rect 11848 -2393 11880 -2359
rect 12178 -2390 12180 -2356
rect 12180 -2390 12212 -2356
rect 12258 -2390 12260 -2356
rect 12260 -2390 12292 -2356
rect 12338 -2390 12340 -2356
rect 12340 -2390 12372 -2356
rect 12418 -2390 12420 -2356
rect 12420 -2390 12452 -2356
rect 12498 -2390 12500 -2356
rect 12500 -2390 12532 -2356
rect 12578 -2390 12580 -2356
rect 12580 -2390 12612 -2356
rect 12738 -2366 12772 -2306
rect 12826 -2366 12860 -2306
<< metal1 >>
rect 725 3732 815 3748
rect 7434 3732 7524 3748
rect 725 3721 744 3732
rect 707 3699 744 3721
rect 598 3687 644 3699
rect 598 3627 604 3687
rect 638 3627 644 3687
rect 598 3549 644 3627
rect 686 3687 744 3699
rect 686 3627 692 3687
rect 726 3680 744 3687
rect 796 3729 815 3732
rect 796 3723 1404 3729
rect 796 3680 842 3723
rect 726 3671 842 3680
rect 894 3671 922 3723
rect 974 3671 1002 3723
rect 1054 3671 1082 3723
rect 1134 3671 1162 3723
rect 1214 3671 1242 3723
rect 1294 3671 1404 3723
rect 726 3663 1404 3671
rect 1466 3726 6374 3732
rect 1466 3674 1574 3726
rect 1626 3674 1654 3726
rect 1706 3674 1734 3726
rect 1786 3674 1814 3726
rect 1866 3674 1894 3726
rect 1946 3674 1974 3726
rect 2026 3674 2178 3726
rect 2230 3674 2258 3726
rect 2310 3674 2338 3726
rect 2390 3674 2418 3726
rect 2470 3674 2498 3726
rect 2550 3674 2578 3726
rect 2630 3674 2786 3726
rect 2838 3674 2866 3726
rect 2918 3674 2946 3726
rect 2998 3674 3026 3726
rect 3078 3674 3106 3726
rect 3158 3674 3186 3726
rect 3238 3674 3390 3726
rect 3442 3674 3470 3726
rect 3522 3674 3550 3726
rect 3602 3674 3630 3726
rect 3682 3674 3710 3726
rect 3762 3674 3790 3726
rect 3842 3674 3998 3726
rect 4050 3674 4078 3726
rect 4130 3674 4158 3726
rect 4210 3674 4238 3726
rect 4290 3674 4318 3726
rect 4370 3674 4398 3726
rect 4450 3674 4602 3726
rect 4654 3674 4682 3726
rect 4734 3674 4762 3726
rect 4814 3674 4842 3726
rect 4894 3674 4922 3726
rect 4974 3674 5002 3726
rect 5054 3674 5210 3726
rect 5262 3674 5290 3726
rect 5342 3674 5370 3726
rect 5422 3674 5450 3726
rect 5502 3674 5530 3726
rect 5582 3674 5610 3726
rect 5662 3674 5814 3726
rect 5866 3674 5894 3726
rect 5946 3674 5974 3726
rect 6026 3674 6054 3726
rect 6106 3674 6134 3726
rect 6186 3674 6214 3726
rect 6266 3674 6374 3726
rect 7434 3721 7453 3732
rect 7416 3699 7453 3721
rect 1466 3666 6374 3674
rect 6534 3670 6624 3686
rect 726 3633 760 3663
rect 726 3627 732 3633
rect 686 3615 732 3627
rect 6534 3618 6553 3670
rect 6605 3618 6624 3670
rect 6534 3602 6624 3618
rect 7011 3673 7101 3689
rect 7011 3621 7030 3673
rect 7082 3621 7101 3673
rect 7011 3605 7101 3621
rect 7307 3687 7353 3699
rect 7307 3627 7313 3687
rect 7347 3627 7353 3687
rect 598 3489 604 3549
rect 638 3489 644 3549
rect 598 3477 644 3489
rect 686 3549 732 3561
rect 686 3489 692 3549
rect 726 3489 732 3549
rect 7307 3549 7353 3627
rect 7395 3687 7453 3699
rect 7395 3627 7401 3687
rect 7435 3680 7453 3687
rect 7505 3729 7524 3732
rect 7505 3723 8113 3729
rect 7505 3680 7551 3723
rect 7435 3671 7551 3680
rect 7603 3671 7631 3723
rect 7683 3671 7711 3723
rect 7763 3671 7791 3723
rect 7843 3671 7871 3723
rect 7923 3671 7951 3723
rect 8003 3671 8113 3723
rect 7435 3663 8113 3671
rect 8175 3726 13083 3732
rect 8175 3674 8283 3726
rect 8335 3674 8363 3726
rect 8415 3674 8443 3726
rect 8495 3674 8523 3726
rect 8575 3674 8603 3726
rect 8655 3674 8683 3726
rect 8735 3674 8887 3726
rect 8939 3674 8967 3726
rect 9019 3674 9047 3726
rect 9099 3674 9127 3726
rect 9179 3674 9207 3726
rect 9259 3674 9287 3726
rect 9339 3674 9495 3726
rect 9547 3674 9575 3726
rect 9627 3674 9655 3726
rect 9707 3674 9735 3726
rect 9787 3674 9815 3726
rect 9867 3674 9895 3726
rect 9947 3674 10099 3726
rect 10151 3674 10179 3726
rect 10231 3674 10259 3726
rect 10311 3674 10339 3726
rect 10391 3674 10419 3726
rect 10471 3674 10499 3726
rect 10551 3674 10707 3726
rect 10759 3674 10787 3726
rect 10839 3674 10867 3726
rect 10919 3674 10947 3726
rect 10999 3674 11027 3726
rect 11079 3674 11107 3726
rect 11159 3674 11311 3726
rect 11363 3674 11391 3726
rect 11443 3674 11471 3726
rect 11523 3674 11551 3726
rect 11603 3674 11631 3726
rect 11683 3674 11711 3726
rect 11763 3674 11919 3726
rect 11971 3674 11999 3726
rect 12051 3674 12079 3726
rect 12131 3674 12159 3726
rect 12211 3674 12239 3726
rect 12291 3674 12319 3726
rect 12371 3674 12523 3726
rect 12575 3674 12603 3726
rect 12655 3674 12683 3726
rect 12735 3674 12763 3726
rect 12815 3674 12843 3726
rect 12895 3674 12923 3726
rect 12975 3674 13083 3726
rect 8175 3666 13083 3674
rect 13243 3670 13333 3686
rect 7435 3633 7469 3663
rect 7435 3627 7441 3633
rect 7395 3615 7441 3627
rect 13243 3618 13262 3670
rect 13314 3618 13333 3670
rect 13243 3602 13333 3618
rect 598 3411 644 3423
rect 598 3351 604 3411
rect 638 3351 644 3411
rect 598 3273 644 3351
rect 686 3411 732 3489
rect 6539 3526 6629 3542
rect 6539 3474 6558 3526
rect 6610 3474 6629 3526
rect 6539 3458 6629 3474
rect 7000 3501 7090 3517
rect 7000 3449 7019 3501
rect 7071 3449 7090 3501
rect 7307 3489 7313 3549
rect 7347 3489 7353 3549
rect 7307 3477 7353 3489
rect 7395 3549 7441 3561
rect 7395 3489 7401 3549
rect 7435 3489 7441 3549
rect 7000 3433 7090 3449
rect 686 3351 692 3411
rect 726 3351 732 3411
rect 7307 3411 7353 3423
rect 686 3339 732 3351
rect 6540 3374 6630 3390
rect 6540 3322 6559 3374
rect 6611 3322 6630 3374
rect 7307 3351 7313 3411
rect 7347 3351 7353 3411
rect 6540 3306 6630 3322
rect 7000 3309 7090 3325
rect 598 3213 604 3273
rect 638 3213 644 3273
rect 598 3201 644 3213
rect 686 3273 732 3285
rect 686 3213 692 3273
rect 726 3213 732 3273
rect 7000 3257 7019 3309
rect 7071 3257 7090 3309
rect 7000 3241 7090 3257
rect 7307 3273 7353 3351
rect 7395 3411 7441 3489
rect 13248 3526 13338 3542
rect 13248 3474 13267 3526
rect 13319 3474 13338 3526
rect 13248 3458 13338 3474
rect 7395 3351 7401 3411
rect 7435 3351 7441 3411
rect 7395 3339 7441 3351
rect 13249 3374 13339 3390
rect 13249 3322 13268 3374
rect 13320 3322 13339 3374
rect 13249 3306 13339 3322
rect 62 3127 522 3147
rect 62 3116 127 3127
rect 62 3082 91 3116
rect 125 3082 127 3116
rect 62 3075 127 3082
rect 179 3126 402 3127
rect 179 3116 258 3126
rect 310 3116 402 3126
rect 179 3082 183 3116
rect 217 3082 258 3116
rect 310 3082 367 3116
rect 401 3082 402 3116
rect 179 3075 258 3082
rect 62 3074 258 3075
rect 310 3075 402 3082
rect 454 3116 522 3127
rect 454 3082 459 3116
rect 493 3082 522 3116
rect 454 3075 522 3082
rect 310 3074 522 3075
rect 62 3051 522 3074
rect 598 3135 644 3147
rect 598 3075 604 3135
rect 638 3075 644 3135
rect 598 2997 644 3075
rect 686 3135 732 3213
rect 6540 3204 6630 3220
rect 6540 3152 6559 3204
rect 6611 3152 6630 3204
rect 7307 3213 7313 3273
rect 7347 3213 7353 3273
rect 7307 3201 7353 3213
rect 7395 3273 7441 3285
rect 7395 3213 7401 3273
rect 7435 3213 7441 3273
rect 6540 3136 6630 3152
rect 686 3075 692 3135
rect 726 3075 732 3135
rect 686 3063 732 3075
rect 6771 3127 7231 3147
rect 6771 3116 6836 3127
rect 6771 3082 6800 3116
rect 6834 3082 6836 3116
rect 6771 3075 6836 3082
rect 6888 3126 7111 3127
rect 6888 3116 6967 3126
rect 7019 3116 7111 3126
rect 6888 3082 6892 3116
rect 6926 3082 6967 3116
rect 7019 3082 7076 3116
rect 7110 3082 7111 3116
rect 6888 3075 6967 3082
rect 6771 3074 6967 3075
rect 7019 3075 7111 3082
rect 7163 3116 7231 3127
rect 7163 3082 7168 3116
rect 7202 3082 7231 3116
rect 7163 3075 7231 3082
rect 7019 3074 7231 3075
rect 6539 3047 6629 3063
rect 6771 3051 7231 3074
rect 7307 3135 7353 3147
rect 7307 3075 7313 3135
rect 7347 3075 7353 3135
rect 207 2973 570 2980
rect 207 2939 219 2973
rect 253 2952 570 2973
rect 253 2939 265 2952
rect 207 2932 265 2939
rect 312 2918 379 2924
rect 312 2884 328 2918
rect 362 2905 379 2918
rect 362 2884 514 2905
rect 312 2877 514 2884
rect 392 2816 458 2818
rect 130 2811 184 2815
rect 129 2808 184 2811
rect 0 2774 138 2808
rect 172 2774 184 2808
rect 129 2771 184 2774
rect 129 2767 183 2771
rect 392 2764 400 2816
rect 452 2764 458 2816
rect 392 2763 458 2764
rect 486 2733 514 2877
rect 542 2820 570 2952
rect 598 2937 604 2997
rect 638 2937 644 2997
rect 598 2925 644 2937
rect 686 2997 789 3009
rect 686 2937 692 2997
rect 726 2937 789 2997
rect 6539 2995 6558 3047
rect 6610 2995 6629 3047
rect 6539 2979 6629 2995
rect 7307 2997 7353 3075
rect 7395 3135 7441 3213
rect 13249 3204 13339 3220
rect 13249 3152 13268 3204
rect 13320 3152 13339 3204
rect 13249 3136 13339 3152
rect 7395 3075 7401 3135
rect 7435 3075 7441 3135
rect 7395 3063 7441 3075
rect 13248 3047 13338 3063
rect 686 2925 789 2937
rect 6916 2973 7279 2980
rect 6916 2939 6928 2973
rect 6962 2952 7279 2973
rect 6962 2939 6974 2952
rect 6916 2932 6974 2939
rect 636 2878 705 2884
rect 636 2844 648 2878
rect 682 2844 705 2878
rect 636 2838 705 2844
rect 542 2808 591 2820
rect 542 2774 551 2808
rect 585 2774 591 2808
rect 542 2761 591 2774
rect 486 2715 629 2733
rect 486 2705 589 2715
rect 580 2681 589 2705
rect 623 2681 629 2715
rect 580 2668 629 2681
rect 62 2581 522 2603
rect 62 2572 145 2581
rect 197 2572 265 2581
rect 317 2572 408 2581
rect 460 2572 522 2581
rect 62 2538 91 2572
rect 125 2538 145 2572
rect 217 2538 265 2572
rect 317 2538 367 2572
rect 401 2538 408 2572
rect 493 2538 522 2572
rect 62 2529 145 2538
rect 197 2529 265 2538
rect 317 2529 408 2538
rect 460 2529 522 2538
rect 62 2507 522 2529
rect 657 2438 705 2838
rect 37 2391 705 2438
rect 657 2250 705 2391
rect 647 2244 705 2250
rect 406 2238 471 2239
rect 406 2237 412 2238
rect 310 2235 412 2237
rect 308 2189 412 2235
rect 406 2186 412 2189
rect 464 2186 471 2238
rect 647 2210 659 2244
rect 693 2210 705 2244
rect 647 2204 705 2210
rect 743 2435 789 2925
rect 7021 2918 7088 2924
rect 7021 2884 7037 2918
rect 7071 2905 7088 2918
rect 7071 2884 7223 2905
rect 7021 2877 7223 2884
rect 6457 2805 6547 2821
rect 7101 2816 7167 2818
rect 6839 2811 6893 2815
rect 6838 2808 6893 2811
rect 6457 2794 6476 2805
rect 6382 2753 6476 2794
rect 6528 2753 6547 2805
rect 6709 2774 6847 2808
rect 6881 2774 6893 2808
rect 6838 2771 6893 2774
rect 6838 2767 6892 2771
rect 7101 2764 7109 2816
rect 7161 2764 7167 2816
rect 7101 2763 7167 2764
rect 839 2738 888 2745
rect 839 2733 1458 2738
rect 839 2699 848 2733
rect 882 2699 1458 2733
rect 839 2691 1458 2699
rect 839 2686 888 2691
rect 840 2644 889 2652
rect 1409 2644 1458 2691
rect 6382 2735 6547 2753
rect 6382 2689 6429 2735
rect 7195 2733 7223 2877
rect 7251 2820 7279 2952
rect 7307 2937 7313 2997
rect 7347 2937 7353 2997
rect 7307 2925 7353 2937
rect 7395 2997 7498 3009
rect 7395 2937 7401 2997
rect 7435 2937 7498 2997
rect 13248 2995 13267 3047
rect 13319 2995 13338 3047
rect 13248 2979 13338 2995
rect 7395 2925 7498 2937
rect 7345 2878 7414 2884
rect 7345 2844 7357 2878
rect 7391 2844 7414 2878
rect 7345 2838 7414 2844
rect 7251 2808 7300 2820
rect 7251 2774 7260 2808
rect 7294 2774 7300 2808
rect 7251 2761 7300 2774
rect 7195 2715 7338 2733
rect 7195 2705 7298 2715
rect 6383 2686 6429 2689
rect 840 2640 1341 2644
rect 840 2606 849 2640
rect 883 2635 1341 2640
rect 883 2606 1290 2635
rect 840 2601 1290 2606
rect 1324 2601 1341 2635
rect 840 2598 1341 2601
rect 1409 2638 5830 2644
rect 1409 2604 2022 2638
rect 2056 2604 2148 2638
rect 2182 2604 3234 2638
rect 3268 2604 3360 2638
rect 3394 2604 4446 2638
rect 4480 2604 4572 2638
rect 4606 2604 5658 2638
rect 5692 2604 5784 2638
rect 5818 2604 5830 2638
rect 6383 2626 6389 2686
rect 6423 2626 6429 2686
rect 6383 2614 6429 2626
rect 6471 2686 6517 2698
rect 6471 2626 6477 2686
rect 6511 2626 6517 2686
rect 7289 2681 7298 2705
rect 7332 2681 7338 2715
rect 7289 2668 7338 2681
rect 6471 2617 6517 2626
rect 1409 2598 5830 2604
rect 840 2597 1336 2598
rect 1409 2597 1855 2598
rect 840 2593 889 2597
rect 1278 2595 1336 2597
rect 6471 2588 6709 2617
rect 1240 2546 1286 2554
rect 1217 2545 1296 2546
rect 1217 2481 1224 2545
rect 1288 2481 1296 2545
rect 1328 2545 1374 2557
rect 1972 2549 2018 2557
rect 1328 2485 1334 2545
rect 1368 2485 1374 2545
rect 1240 2470 1286 2481
rect 1328 2435 1374 2485
rect 1949 2548 2028 2549
rect 1949 2484 1956 2548
rect 2020 2484 2028 2548
rect 2077 2545 2123 2557
rect 2186 2549 2232 2557
rect 3184 2549 3230 2557
rect 2077 2485 2083 2545
rect 2117 2485 2123 2545
rect 1972 2473 2018 2484
rect 2077 2435 2123 2485
rect 2176 2548 2255 2549
rect 2176 2484 2184 2548
rect 2248 2484 2255 2548
rect 3161 2548 3240 2549
rect 3161 2484 3168 2548
rect 3232 2484 3240 2548
rect 3288 2545 3334 2557
rect 3398 2549 3444 2557
rect 4396 2549 4442 2557
rect 3288 2485 3294 2545
rect 3328 2485 3334 2545
rect 2186 2473 2232 2484
rect 3184 2473 3230 2484
rect 3288 2435 3334 2485
rect 3388 2548 3467 2549
rect 3388 2484 3396 2548
rect 3460 2484 3467 2548
rect 4373 2548 4452 2549
rect 4373 2484 4380 2548
rect 4444 2484 4452 2548
rect 4501 2545 4547 2557
rect 4610 2549 4656 2557
rect 5608 2549 5654 2557
rect 4501 2485 4507 2545
rect 4541 2485 4547 2545
rect 3398 2473 3444 2484
rect 4396 2473 4442 2484
rect 4501 2435 4547 2485
rect 4600 2548 4679 2549
rect 4600 2484 4608 2548
rect 4672 2484 4679 2548
rect 5585 2548 5664 2549
rect 5585 2484 5592 2548
rect 5656 2484 5664 2548
rect 5715 2545 5761 2557
rect 5822 2549 5868 2557
rect 5715 2485 5721 2545
rect 5755 2485 5761 2545
rect 4610 2473 4656 2484
rect 5608 2473 5654 2484
rect 5715 2435 5761 2485
rect 5812 2548 5891 2549
rect 5812 2484 5820 2548
rect 5884 2484 5891 2548
rect 6383 2548 6429 2560
rect 6383 2488 6389 2548
rect 6423 2488 6429 2548
rect 5822 2473 5868 2484
rect 6383 2476 6429 2488
rect 6471 2548 6517 2588
rect 6471 2488 6477 2548
rect 6511 2488 6517 2548
rect 6471 2476 6517 2488
rect 6545 2548 6635 2560
rect 6545 2544 6573 2548
rect 6607 2544 6635 2548
rect 6545 2492 6564 2544
rect 6616 2492 6635 2544
rect 6545 2488 6573 2492
rect 6607 2488 6635 2492
rect 6545 2476 6635 2488
rect 6663 2548 6709 2588
rect 6663 2488 6669 2548
rect 6703 2488 6709 2548
rect 6771 2581 7231 2603
rect 6771 2572 6854 2581
rect 6906 2572 6974 2581
rect 7026 2572 7117 2581
rect 7169 2572 7231 2581
rect 6771 2538 6800 2572
rect 6834 2538 6854 2572
rect 6926 2538 6974 2572
rect 7026 2538 7076 2572
rect 7110 2538 7117 2572
rect 7202 2538 7231 2572
rect 6771 2529 6854 2538
rect 6906 2529 6974 2538
rect 7026 2529 7117 2538
rect 7169 2529 7231 2538
rect 6771 2507 7231 2529
rect 6663 2476 6709 2488
rect 6302 2435 6368 2437
rect 743 2431 6368 2435
rect 743 2397 6318 2431
rect 6352 2397 6368 2431
rect 743 2393 6368 2397
rect 743 2172 789 2393
rect 1593 2346 1639 2356
rect 1571 2282 1580 2346
rect 1644 2282 1653 2346
rect 1571 2281 1653 2282
rect 1683 2344 1729 2393
rect 2325 2346 2371 2356
rect 1683 2284 1689 2344
rect 1723 2284 1729 2344
rect 1593 2272 1639 2281
rect 1683 2272 1729 2284
rect 2303 2282 2312 2346
rect 2376 2282 2385 2346
rect 2303 2281 2385 2282
rect 2432 2344 2478 2393
rect 2535 2346 2581 2356
rect 3537 2346 3583 2356
rect 2432 2284 2438 2344
rect 2472 2284 2478 2344
rect 2325 2272 2371 2281
rect 2432 2272 2478 2284
rect 2521 2282 2530 2346
rect 2594 2282 2603 2346
rect 2521 2281 2603 2282
rect 3515 2282 3524 2346
rect 3588 2282 3597 2346
rect 3515 2281 3597 2282
rect 3643 2344 3689 2393
rect 3747 2346 3793 2356
rect 4875 2346 4921 2356
rect 3643 2284 3649 2344
rect 3683 2284 3689 2344
rect 2535 2272 2581 2281
rect 3537 2272 3583 2281
rect 3643 2272 3689 2284
rect 3733 2282 3742 2346
rect 3806 2282 3815 2346
rect 3733 2281 3815 2282
rect 4853 2282 4862 2346
rect 4926 2282 4935 2346
rect 4853 2281 4935 2282
rect 4983 2344 5029 2393
rect 5085 2346 5131 2356
rect 4983 2284 4989 2344
rect 5023 2284 5029 2344
rect 3747 2272 3793 2281
rect 4875 2272 4921 2281
rect 4983 2272 5029 2284
rect 5071 2282 5080 2346
rect 5144 2282 5153 2346
rect 5071 2281 5153 2282
rect 5730 2344 5776 2393
rect 6306 2391 6368 2393
rect 6401 2428 6429 2476
rect 7366 2438 7414 2838
rect 6685 2435 7414 2438
rect 6513 2429 7414 2435
rect 6513 2428 6525 2429
rect 6401 2399 6525 2428
rect 6401 2357 6429 2399
rect 6513 2395 6525 2399
rect 6559 2395 7414 2429
rect 6513 2391 7414 2395
rect 6513 2389 6755 2391
rect 6685 2386 6755 2389
rect 5819 2346 5865 2356
rect 5730 2284 5736 2344
rect 5770 2284 5776 2344
rect 5085 2272 5131 2281
rect 5730 2272 5776 2284
rect 5805 2282 5814 2346
rect 5878 2282 5887 2346
rect 5805 2281 5887 2282
rect 6383 2345 6429 2357
rect 6383 2285 6389 2345
rect 6423 2285 6429 2345
rect 5819 2272 5865 2281
rect 6383 2273 6429 2285
rect 6471 2345 6517 2357
rect 6471 2285 6477 2345
rect 6511 2285 6517 2345
rect 6471 2245 6517 2285
rect 6545 2345 6635 2357
rect 6545 2341 6573 2345
rect 6607 2341 6635 2345
rect 6545 2289 6564 2341
rect 6616 2289 6635 2341
rect 6545 2285 6573 2289
rect 6607 2285 6635 2289
rect 6545 2273 6635 2285
rect 6663 2345 6709 2357
rect 6663 2285 6669 2345
rect 6703 2285 6709 2345
rect 6663 2245 6709 2285
rect 7366 2250 7414 2391
rect 5771 2240 5830 2243
rect 893 2186 900 2238
rect 952 2236 958 2238
rect 1631 2236 1689 2240
rect 952 2234 1689 2236
rect 952 2200 1643 2234
rect 1677 2219 1689 2234
rect 2363 2234 3759 2240
rect 1677 2200 1691 2219
rect 952 2189 1691 2200
rect 2363 2200 2375 2234
rect 2409 2200 2497 2234
rect 2531 2200 3587 2234
rect 3621 2200 3709 2234
rect 3743 2200 3759 2234
rect 2363 2194 3759 2200
rect 4913 2234 5097 2240
rect 4913 2200 4925 2234
rect 4959 2200 5047 2234
rect 5081 2200 5097 2234
rect 4913 2194 5097 2200
rect 5769 2234 5830 2240
rect 5769 2200 5781 2234
rect 5815 2200 5830 2234
rect 5769 2194 5830 2200
rect 952 2186 958 2189
rect 893 2185 958 2186
rect 1633 2184 1691 2189
rect 573 2160 619 2172
rect 573 2100 579 2160
rect 613 2100 619 2160
rect 573 2022 619 2100
rect 733 2160 789 2172
rect 733 2100 739 2160
rect 773 2100 789 2160
rect 733 2088 789 2100
rect 573 1962 579 2022
rect 613 1962 619 2022
rect 573 1950 619 1962
rect 733 2022 779 2034
rect 733 1962 739 2022
rect 773 1962 779 2022
rect 573 1884 619 1896
rect 573 1824 579 1884
rect 613 1824 619 1884
rect 573 1746 619 1824
rect 733 1884 779 1962
rect 733 1824 739 1884
rect 773 1824 779 1884
rect 733 1812 779 1824
rect 88 1700 186 1715
rect 88 1644 105 1700
rect 165 1644 186 1700
rect 573 1686 579 1746
rect 613 1686 619 1746
rect 573 1674 619 1686
rect 733 1746 779 1758
rect 733 1686 739 1746
rect 773 1686 779 1746
rect 88 1625 186 1644
rect 573 1608 619 1620
rect 573 1548 579 1608
rect 613 1548 619 1608
rect 573 1470 619 1548
rect 733 1608 779 1686
rect 733 1548 739 1608
rect 773 1548 779 1608
rect 733 1536 779 1548
rect 573 1410 579 1470
rect 613 1410 619 1470
rect 573 1398 619 1410
rect 733 1470 779 1482
rect 733 1410 739 1470
rect 773 1410 779 1470
rect 573 1332 619 1344
rect 573 1272 579 1332
rect 613 1272 619 1332
rect 573 1194 619 1272
rect 733 1332 779 1410
rect 733 1272 739 1332
rect 773 1272 779 1332
rect 733 1260 779 1272
rect 573 1134 579 1194
rect 613 1134 619 1194
rect 733 1194 779 1206
rect 733 1170 739 1194
rect 573 1122 619 1134
rect 694 1154 739 1170
rect 773 1170 779 1194
rect 773 1154 801 1170
rect 694 1102 730 1154
rect 782 1102 801 1154
rect 694 1086 801 1102
rect 1254 1157 1586 1163
rect 1254 1105 1272 1157
rect 1324 1105 1352 1157
rect 1404 1105 1432 1157
rect 1484 1105 1512 1157
rect 1564 1105 1586 1157
rect 1254 1095 1586 1105
rect 1986 1157 2318 1163
rect 1986 1105 2004 1157
rect 2056 1105 2084 1157
rect 2136 1105 2164 1157
rect 2216 1105 2244 1157
rect 2296 1105 2318 1157
rect 1986 1095 2318 1105
rect 2489 1047 2547 2194
rect 2588 1157 2920 1163
rect 2588 1105 2610 1157
rect 2662 1105 2690 1157
rect 2742 1105 2770 1157
rect 2822 1105 2850 1157
rect 2902 1105 2920 1157
rect 2588 1095 2920 1105
rect 3198 1157 3530 1163
rect 3198 1105 3216 1157
rect 3268 1105 3296 1157
rect 3348 1105 3376 1157
rect 3428 1105 3456 1157
rect 3508 1105 3530 1157
rect 3198 1095 3530 1105
rect 3800 1157 4132 1163
rect 3800 1105 3822 1157
rect 3874 1105 3902 1157
rect 3954 1105 3982 1157
rect 4034 1105 4062 1157
rect 4114 1105 4132 1157
rect 3800 1095 4132 1105
rect 4536 1157 4868 1163
rect 4536 1105 4554 1157
rect 4606 1105 4634 1157
rect 4686 1105 4714 1157
rect 4766 1105 4794 1157
rect 4846 1105 4868 1157
rect 4536 1095 4868 1105
rect 283 1019 2547 1047
rect 4915 991 4973 2194
rect 5138 1157 5470 1163
rect 5138 1105 5160 1157
rect 5212 1105 5240 1157
rect 5292 1105 5320 1157
rect 5372 1105 5400 1157
rect 5452 1105 5470 1157
rect 5138 1095 5470 1105
rect 283 963 4973 991
rect 5771 1062 5830 2194
rect 6383 2207 6429 2219
rect 6383 2147 6389 2207
rect 6423 2147 6429 2207
rect 6383 2095 6429 2147
rect 6471 2216 6709 2245
rect 7356 2244 7414 2250
rect 7115 2238 7180 2239
rect 7115 2237 7121 2238
rect 7019 2235 7121 2237
rect 6471 2207 6517 2216
rect 6471 2147 6477 2207
rect 6511 2147 6517 2207
rect 7017 2189 7121 2235
rect 7115 2186 7121 2189
rect 7173 2186 7180 2238
rect 7356 2210 7368 2244
rect 7402 2210 7414 2244
rect 7356 2204 7414 2210
rect 7452 2435 7498 2925
rect 13166 2805 13256 2821
rect 13166 2794 13185 2805
rect 13091 2753 13185 2794
rect 13237 2753 13256 2805
rect 7548 2738 7597 2745
rect 7548 2733 8167 2738
rect 7548 2699 7557 2733
rect 7591 2699 8167 2733
rect 7548 2691 8167 2699
rect 7548 2686 7597 2691
rect 7549 2644 7598 2652
rect 8118 2644 8167 2691
rect 13091 2735 13256 2753
rect 13091 2689 13138 2735
rect 13092 2686 13138 2689
rect 7549 2640 8050 2644
rect 7549 2606 7558 2640
rect 7592 2635 8050 2640
rect 7592 2606 7999 2635
rect 7549 2601 7999 2606
rect 8033 2601 8050 2635
rect 7549 2598 8050 2601
rect 8118 2638 12539 2644
rect 8118 2604 8731 2638
rect 8765 2604 8857 2638
rect 8891 2604 9943 2638
rect 9977 2604 10069 2638
rect 10103 2604 11155 2638
rect 11189 2604 11281 2638
rect 11315 2604 12367 2638
rect 12401 2604 12493 2638
rect 12527 2604 12539 2638
rect 13092 2626 13098 2686
rect 13132 2626 13138 2686
rect 13092 2614 13138 2626
rect 13180 2686 13226 2698
rect 13180 2626 13186 2686
rect 13220 2626 13226 2686
rect 13180 2617 13226 2626
rect 8118 2598 12539 2604
rect 7549 2597 8045 2598
rect 8118 2597 8564 2598
rect 7549 2593 7598 2597
rect 7987 2595 8045 2597
rect 13180 2588 13418 2617
rect 7949 2546 7995 2554
rect 7926 2545 8005 2546
rect 7926 2481 7933 2545
rect 7997 2481 8005 2545
rect 8037 2545 8083 2557
rect 8681 2549 8727 2557
rect 8037 2485 8043 2545
rect 8077 2485 8083 2545
rect 7949 2470 7995 2481
rect 8037 2435 8083 2485
rect 8658 2548 8737 2549
rect 8658 2484 8665 2548
rect 8729 2484 8737 2548
rect 8786 2545 8832 2557
rect 8895 2549 8941 2557
rect 9893 2549 9939 2557
rect 8786 2485 8792 2545
rect 8826 2485 8832 2545
rect 8681 2473 8727 2484
rect 8786 2435 8832 2485
rect 8885 2548 8964 2549
rect 8885 2484 8893 2548
rect 8957 2484 8964 2548
rect 9870 2548 9949 2549
rect 9870 2484 9877 2548
rect 9941 2484 9949 2548
rect 9997 2545 10043 2557
rect 10107 2549 10153 2557
rect 11105 2549 11151 2557
rect 9997 2485 10003 2545
rect 10037 2485 10043 2545
rect 8895 2473 8941 2484
rect 9893 2473 9939 2484
rect 9997 2435 10043 2485
rect 10097 2548 10176 2549
rect 10097 2484 10105 2548
rect 10169 2484 10176 2548
rect 11082 2548 11161 2549
rect 11082 2484 11089 2548
rect 11153 2484 11161 2548
rect 11210 2545 11256 2557
rect 11319 2549 11365 2557
rect 12317 2549 12363 2557
rect 11210 2485 11216 2545
rect 11250 2485 11256 2545
rect 10107 2473 10153 2484
rect 11105 2473 11151 2484
rect 11210 2435 11256 2485
rect 11309 2548 11388 2549
rect 11309 2484 11317 2548
rect 11381 2484 11388 2548
rect 12294 2548 12373 2549
rect 12294 2484 12301 2548
rect 12365 2484 12373 2548
rect 12424 2545 12470 2557
rect 12531 2549 12577 2557
rect 12424 2485 12430 2545
rect 12464 2485 12470 2545
rect 11319 2473 11365 2484
rect 12317 2473 12363 2484
rect 12424 2435 12470 2485
rect 12521 2548 12600 2549
rect 12521 2484 12529 2548
rect 12593 2484 12600 2548
rect 13092 2548 13138 2560
rect 13092 2488 13098 2548
rect 13132 2488 13138 2548
rect 12531 2473 12577 2484
rect 13092 2476 13138 2488
rect 13180 2548 13226 2588
rect 13180 2488 13186 2548
rect 13220 2488 13226 2548
rect 13180 2476 13226 2488
rect 13254 2548 13344 2560
rect 13254 2544 13282 2548
rect 13316 2544 13344 2548
rect 13254 2492 13273 2544
rect 13325 2492 13344 2544
rect 13254 2488 13282 2492
rect 13316 2488 13344 2492
rect 13254 2476 13344 2488
rect 13372 2548 13418 2588
rect 13372 2488 13378 2548
rect 13412 2488 13418 2548
rect 13372 2476 13418 2488
rect 13011 2435 13077 2437
rect 7452 2431 13077 2435
rect 7452 2397 13027 2431
rect 13061 2397 13077 2431
rect 7452 2393 13077 2397
rect 7452 2172 7498 2393
rect 8302 2346 8348 2356
rect 8280 2282 8289 2346
rect 8353 2282 8362 2346
rect 8280 2281 8362 2282
rect 8392 2344 8438 2393
rect 9034 2346 9080 2356
rect 8392 2284 8398 2344
rect 8432 2284 8438 2344
rect 8302 2272 8348 2281
rect 8392 2272 8438 2284
rect 9012 2282 9021 2346
rect 9085 2282 9094 2346
rect 9012 2281 9094 2282
rect 9141 2344 9187 2393
rect 9244 2346 9290 2356
rect 10246 2346 10292 2356
rect 9141 2284 9147 2344
rect 9181 2284 9187 2344
rect 9034 2272 9080 2281
rect 9141 2272 9187 2284
rect 9230 2282 9239 2346
rect 9303 2282 9312 2346
rect 9230 2281 9312 2282
rect 10224 2282 10233 2346
rect 10297 2282 10306 2346
rect 10224 2281 10306 2282
rect 10352 2344 10398 2393
rect 10456 2346 10502 2356
rect 11584 2346 11630 2356
rect 10352 2284 10358 2344
rect 10392 2284 10398 2344
rect 9244 2272 9290 2281
rect 10246 2272 10292 2281
rect 10352 2272 10398 2284
rect 10442 2282 10451 2346
rect 10515 2282 10524 2346
rect 10442 2281 10524 2282
rect 11562 2282 11571 2346
rect 11635 2282 11644 2346
rect 11562 2281 11644 2282
rect 11692 2344 11738 2393
rect 11794 2346 11840 2356
rect 11692 2284 11698 2344
rect 11732 2284 11738 2344
rect 10456 2272 10502 2281
rect 11584 2272 11630 2281
rect 11692 2272 11738 2284
rect 11780 2282 11789 2346
rect 11853 2282 11862 2346
rect 11780 2281 11862 2282
rect 12439 2344 12485 2393
rect 13015 2391 13077 2393
rect 13110 2428 13138 2476
rect 13222 2429 13492 2435
rect 13222 2428 13234 2429
rect 13110 2399 13234 2428
rect 13110 2357 13138 2399
rect 13222 2395 13234 2399
rect 13268 2395 13492 2429
rect 13222 2389 13492 2395
rect 12528 2346 12574 2356
rect 12439 2284 12445 2344
rect 12479 2284 12485 2344
rect 11794 2272 11840 2281
rect 12439 2272 12485 2284
rect 12514 2282 12523 2346
rect 12587 2282 12596 2346
rect 12514 2281 12596 2282
rect 13092 2345 13138 2357
rect 13092 2285 13098 2345
rect 13132 2285 13138 2345
rect 12528 2272 12574 2281
rect 13092 2273 13138 2285
rect 13180 2345 13226 2357
rect 13180 2285 13186 2345
rect 13220 2285 13226 2345
rect 13180 2245 13226 2285
rect 13254 2345 13344 2357
rect 13254 2341 13282 2345
rect 13316 2341 13344 2345
rect 13254 2289 13273 2341
rect 13325 2289 13344 2341
rect 13254 2285 13282 2289
rect 13316 2285 13344 2289
rect 13254 2273 13344 2285
rect 13372 2345 13418 2357
rect 13372 2285 13378 2345
rect 13412 2285 13418 2345
rect 13372 2245 13418 2285
rect 12480 2240 12539 2243
rect 7602 2186 7609 2238
rect 7661 2236 7667 2238
rect 8340 2236 8398 2240
rect 7661 2234 8398 2236
rect 7661 2200 8352 2234
rect 8386 2219 8398 2234
rect 9072 2234 10468 2240
rect 8386 2200 8400 2219
rect 7661 2189 8400 2200
rect 9072 2200 9084 2234
rect 9118 2200 9206 2234
rect 9240 2200 10296 2234
rect 10330 2200 10418 2234
rect 10452 2200 10468 2234
rect 9072 2194 10468 2200
rect 11622 2234 11806 2240
rect 11622 2200 11634 2234
rect 11668 2200 11756 2234
rect 11790 2200 11806 2234
rect 11622 2194 11806 2200
rect 12478 2234 12539 2240
rect 12478 2200 12490 2234
rect 12524 2200 12539 2234
rect 12478 2194 12539 2200
rect 7661 2186 7667 2189
rect 7602 2185 7667 2186
rect 8342 2184 8400 2189
rect 6471 2135 6517 2147
rect 7282 2160 7328 2172
rect 7282 2100 7288 2160
rect 7322 2100 7328 2160
rect 6383 2079 6544 2095
rect 6383 2027 6473 2079
rect 6525 2027 6544 2079
rect 6383 2011 6544 2027
rect 7282 2022 7328 2100
rect 7442 2160 7498 2172
rect 7442 2100 7448 2160
rect 7482 2100 7498 2160
rect 7442 2088 7498 2100
rect 7282 1962 7288 2022
rect 7322 1962 7328 2022
rect 7282 1950 7328 1962
rect 7442 2022 7488 2034
rect 7442 1962 7448 2022
rect 7482 1962 7488 2022
rect 7282 1884 7328 1896
rect 7282 1824 7288 1884
rect 7322 1824 7328 1884
rect 7282 1746 7328 1824
rect 7442 1884 7488 1962
rect 7442 1824 7448 1884
rect 7482 1824 7488 1884
rect 7442 1812 7488 1824
rect 7282 1686 7288 1746
rect 7322 1686 7328 1746
rect 7282 1674 7328 1686
rect 7442 1746 7488 1758
rect 7442 1686 7448 1746
rect 7482 1686 7488 1746
rect 7282 1608 7328 1620
rect 7282 1548 7288 1608
rect 7322 1548 7328 1608
rect 7282 1470 7328 1548
rect 7442 1608 7488 1686
rect 7442 1548 7448 1608
rect 7482 1548 7488 1608
rect 7442 1536 7488 1548
rect 7282 1410 7288 1470
rect 7322 1410 7328 1470
rect 7282 1398 7328 1410
rect 7442 1470 7488 1482
rect 7442 1410 7448 1470
rect 7482 1410 7488 1470
rect 7282 1332 7328 1344
rect 7282 1272 7288 1332
rect 7322 1272 7328 1332
rect 7282 1194 7328 1272
rect 7442 1332 7488 1410
rect 7442 1272 7448 1332
rect 7482 1272 7488 1332
rect 7442 1260 7488 1272
rect 5872 1157 6204 1163
rect 5872 1105 5894 1157
rect 5946 1105 5974 1157
rect 6026 1105 6054 1157
rect 6106 1105 6134 1157
rect 6186 1105 6204 1157
rect 7282 1134 7288 1194
rect 7322 1134 7328 1194
rect 7442 1194 7488 1206
rect 7442 1170 7448 1194
rect 7282 1122 7328 1134
rect 7403 1154 7448 1170
rect 7482 1170 7488 1194
rect 7482 1154 7510 1170
rect 5872 1095 6204 1105
rect 7403 1102 7439 1154
rect 7491 1102 7510 1154
rect 7403 1086 7510 1102
rect 7963 1157 8295 1163
rect 7963 1105 7981 1157
rect 8033 1105 8061 1157
rect 8113 1105 8141 1157
rect 8193 1105 8221 1157
rect 8273 1105 8295 1157
rect 7963 1095 8295 1105
rect 8695 1157 9027 1163
rect 8695 1105 8713 1157
rect 8765 1105 8793 1157
rect 8845 1105 8873 1157
rect 8925 1105 8953 1157
rect 9005 1105 9027 1157
rect 8695 1095 9027 1105
rect 5771 935 5829 1062
rect 283 907 5829 935
rect 9198 879 9256 2194
rect 9297 1157 9629 1163
rect 9297 1105 9319 1157
rect 9371 1105 9399 1157
rect 9451 1105 9479 1157
rect 9531 1105 9559 1157
rect 9611 1105 9629 1157
rect 9297 1095 9629 1105
rect 9907 1157 10239 1163
rect 9907 1105 9925 1157
rect 9977 1105 10005 1157
rect 10057 1105 10085 1157
rect 10137 1105 10165 1157
rect 10217 1105 10239 1157
rect 9907 1095 10239 1105
rect 10509 1157 10841 1163
rect 10509 1105 10531 1157
rect 10583 1105 10611 1157
rect 10663 1105 10691 1157
rect 10743 1105 10771 1157
rect 10823 1105 10841 1157
rect 10509 1095 10841 1105
rect 11245 1157 11577 1163
rect 11245 1105 11263 1157
rect 11315 1105 11343 1157
rect 11395 1105 11423 1157
rect 11475 1105 11503 1157
rect 11555 1105 11577 1157
rect 11245 1095 11577 1105
rect 283 851 9256 879
rect 11624 823 11682 2194
rect 11847 1157 12179 1163
rect 11847 1105 11869 1157
rect 11921 1105 11949 1157
rect 12001 1105 12029 1157
rect 12081 1105 12109 1157
rect 12161 1105 12179 1157
rect 11847 1095 12179 1105
rect 283 795 11682 823
rect 12480 1062 12539 2194
rect 13092 2207 13138 2219
rect 13092 2147 13098 2207
rect 13132 2147 13138 2207
rect 13092 2095 13138 2147
rect 13180 2216 13418 2245
rect 13180 2207 13226 2216
rect 13180 2147 13186 2207
rect 13220 2147 13226 2207
rect 13180 2135 13226 2147
rect 13092 2079 13253 2095
rect 13092 2027 13182 2079
rect 13234 2027 13253 2079
rect 13092 2011 13253 2027
rect 12581 1157 12913 1163
rect 12581 1105 12603 1157
rect 12655 1105 12683 1157
rect 12735 1105 12763 1157
rect 12815 1105 12843 1157
rect 12895 1105 12913 1157
rect 12581 1095 12913 1105
rect 12480 767 12538 1062
rect 283 739 12538 767
rect 283 685 12574 711
rect 283 684 12504 685
rect 283 632 900 684
rect 952 677 12504 684
rect 952 674 7609 677
rect 952 632 5800 674
rect 283 622 5800 632
rect 5853 624 7609 674
rect 7661 624 12504 677
rect 5853 622 12504 624
rect 283 621 12504 622
rect 12568 621 12574 685
rect 283 599 12574 621
rect 283 543 10975 571
rect 283 487 8549 515
rect 283 431 7693 459
rect 283 375 4266 403
rect 283 319 1840 347
rect 283 263 984 291
rect 551 216 883 226
rect 551 164 569 216
rect 621 164 649 216
rect 701 164 729 216
rect 781 164 809 216
rect 861 164 883 216
rect 551 158 883 164
rect 211 -706 372 -690
rect 211 -758 230 -706
rect 282 -758 372 -706
rect 211 -774 372 -758
rect 238 -826 284 -814
rect 238 -886 244 -826
rect 278 -886 284 -826
rect 238 -895 284 -886
rect 46 -924 284 -895
rect 326 -826 372 -774
rect 326 -886 332 -826
rect 366 -886 372 -826
rect 326 -898 372 -886
rect 925 -873 984 263
rect 1285 216 1617 226
rect 1285 164 1303 216
rect 1355 164 1383 216
rect 1435 164 1463 216
rect 1515 164 1543 216
rect 1595 164 1617 216
rect 1285 158 1617 164
rect 1782 -873 1840 319
rect 1887 216 2219 226
rect 1887 164 1909 216
rect 1961 164 1989 216
rect 2041 164 2069 216
rect 2121 164 2149 216
rect 2201 164 2219 216
rect 1887 158 2219 164
rect 2623 216 2955 226
rect 2623 164 2641 216
rect 2693 164 2721 216
rect 2773 164 2801 216
rect 2853 164 2881 216
rect 2933 164 2955 216
rect 2623 158 2955 164
rect 3225 216 3557 226
rect 3225 164 3247 216
rect 3299 164 3327 216
rect 3379 164 3407 216
rect 3459 164 3487 216
rect 3539 164 3557 216
rect 3225 158 3557 164
rect 3835 216 4167 226
rect 3835 164 3853 216
rect 3905 164 3933 216
rect 3985 164 4013 216
rect 4065 164 4093 216
rect 4145 164 4167 216
rect 3835 158 4167 164
rect 4208 -873 4266 375
rect 7635 259 7693 431
rect 4437 216 4769 226
rect 4437 164 4459 216
rect 4511 164 4539 216
rect 4591 164 4619 216
rect 4671 164 4699 216
rect 4751 164 4769 216
rect 4437 158 4769 164
rect 5169 216 5501 226
rect 5169 164 5191 216
rect 5243 164 5271 216
rect 5323 164 5351 216
rect 5403 164 5431 216
rect 5483 164 5501 216
rect 5169 158 5501 164
rect 5954 219 6061 235
rect 5954 167 5973 219
rect 6025 167 6061 219
rect 7260 216 7592 226
rect 5954 151 5982 167
rect 5976 127 5982 151
rect 6016 151 6061 167
rect 6136 187 6182 199
rect 6016 127 6022 151
rect 5976 115 6022 127
rect 6136 127 6142 187
rect 6176 127 6182 187
rect 7260 164 7278 216
rect 7330 164 7358 216
rect 7410 164 7438 216
rect 7490 164 7518 216
rect 7570 164 7592 216
rect 7260 158 7592 164
rect 5976 49 6022 61
rect 5976 -11 5982 49
rect 6016 -11 6022 49
rect 5976 -89 6022 -11
rect 6136 49 6182 127
rect 6136 -11 6142 49
rect 6176 -11 6182 49
rect 6136 -23 6182 -11
rect 5976 -149 5982 -89
rect 6016 -149 6022 -89
rect 5976 -161 6022 -149
rect 6136 -89 6182 -77
rect 6136 -149 6142 -89
rect 6176 -149 6182 -89
rect 5976 -227 6022 -215
rect 5976 -287 5982 -227
rect 6016 -287 6022 -227
rect 5976 -365 6022 -287
rect 6136 -227 6182 -149
rect 6136 -287 6142 -227
rect 6176 -287 6182 -227
rect 6136 -299 6182 -287
rect 5976 -425 5982 -365
rect 6016 -425 6022 -365
rect 5976 -437 6022 -425
rect 6136 -365 6182 -353
rect 6136 -425 6142 -365
rect 6176 -425 6182 -365
rect 5976 -503 6022 -491
rect 5976 -563 5982 -503
rect 6016 -563 6022 -503
rect 5976 -641 6022 -563
rect 6136 -503 6182 -425
rect 6136 -563 6142 -503
rect 6176 -563 6182 -503
rect 6136 -575 6182 -563
rect 5976 -701 5982 -641
rect 6016 -701 6022 -641
rect 5976 -713 6022 -701
rect 6136 -641 6182 -629
rect 6136 -701 6142 -641
rect 6176 -701 6182 -641
rect 5966 -779 6022 -767
rect 5966 -839 5982 -779
rect 6016 -839 6022 -779
rect 5966 -851 6022 -839
rect 6136 -779 6182 -701
rect 6920 -706 7081 -690
rect 6920 -758 6939 -706
rect 6991 -758 7081 -706
rect 6920 -774 7081 -758
rect 6136 -839 6142 -779
rect 6176 -839 6182 -779
rect 6136 -851 6182 -839
rect 6947 -826 6993 -814
rect 5064 -868 5122 -863
rect 5797 -865 5862 -864
rect 5797 -868 5803 -865
rect 925 -879 986 -873
rect 925 -913 940 -879
rect 974 -913 986 -879
rect 925 -919 986 -913
rect 1658 -879 1842 -873
rect 1658 -913 1674 -879
rect 1708 -913 1796 -879
rect 1830 -913 1842 -879
rect 1658 -919 1842 -913
rect 2996 -879 4392 -873
rect 2996 -913 3012 -879
rect 3046 -913 3134 -879
rect 3168 -913 4224 -879
rect 4258 -913 4346 -879
rect 4380 -913 4392 -879
rect 5064 -879 5803 -868
rect 5064 -898 5078 -879
rect 2996 -919 4392 -913
rect 5066 -913 5078 -898
rect 5112 -913 5803 -879
rect 5066 -915 5803 -913
rect 5066 -919 5124 -915
rect 5797 -917 5803 -915
rect 5855 -917 5862 -865
rect 925 -922 984 -919
rect 46 -964 92 -924
rect 46 -1024 52 -964
rect 86 -1024 92 -964
rect 46 -1036 92 -1024
rect 120 -964 210 -952
rect 120 -968 148 -964
rect 182 -968 210 -964
rect 120 -1020 139 -968
rect 191 -1020 210 -968
rect 120 -1024 148 -1020
rect 182 -1024 210 -1020
rect 120 -1036 210 -1024
rect 238 -964 284 -924
rect 238 -1024 244 -964
rect 278 -1024 284 -964
rect 238 -1036 284 -1024
rect 326 -964 372 -952
rect 890 -960 936 -951
rect 326 -1024 332 -964
rect 366 -1024 372 -964
rect 326 -1036 372 -1024
rect 868 -961 950 -960
rect 868 -1025 877 -961
rect 941 -1025 950 -961
rect 979 -963 1025 -951
rect 1624 -960 1670 -951
rect 979 -1023 985 -963
rect 1019 -1023 1025 -963
rect 890 -1035 936 -1025
rect 24 -1074 242 -1068
rect 24 -1108 196 -1074
rect 230 -1078 242 -1074
rect 326 -1078 354 -1036
rect 230 -1107 354 -1078
rect 230 -1108 242 -1107
rect 24 -1114 242 -1108
rect 326 -1155 354 -1107
rect 387 -1072 449 -1070
rect 979 -1072 1025 -1023
rect 1602 -961 1684 -960
rect 1602 -1025 1611 -961
rect 1675 -1025 1684 -961
rect 1726 -963 1772 -951
rect 1834 -960 1880 -951
rect 2962 -960 3008 -951
rect 1726 -1023 1732 -963
rect 1766 -1023 1772 -963
rect 1624 -1035 1670 -1025
rect 1726 -1072 1772 -1023
rect 1820 -961 1902 -960
rect 1820 -1025 1829 -961
rect 1893 -1025 1902 -961
rect 2940 -961 3022 -960
rect 2940 -1025 2949 -961
rect 3013 -1025 3022 -961
rect 3066 -963 3112 -951
rect 3172 -960 3218 -951
rect 4174 -960 4220 -951
rect 3066 -1023 3072 -963
rect 3106 -1023 3112 -963
rect 1834 -1035 1880 -1025
rect 2962 -1035 3008 -1025
rect 3066 -1072 3112 -1023
rect 3158 -961 3240 -960
rect 3158 -1025 3167 -961
rect 3231 -1025 3240 -961
rect 4152 -961 4234 -960
rect 4152 -1025 4161 -961
rect 4225 -1025 4234 -961
rect 4277 -963 4323 -951
rect 4384 -960 4430 -951
rect 4277 -1023 4283 -963
rect 4317 -1023 4323 -963
rect 3172 -1035 3218 -1025
rect 4174 -1035 4220 -1025
rect 4277 -1072 4323 -1023
rect 4370 -961 4452 -960
rect 4370 -1025 4379 -961
rect 4443 -1025 4452 -961
rect 5026 -963 5072 -951
rect 5116 -960 5162 -951
rect 5026 -1023 5032 -963
rect 5066 -1023 5072 -963
rect 4384 -1035 4430 -1025
rect 5026 -1072 5072 -1023
rect 5102 -961 5184 -960
rect 5102 -1025 5111 -961
rect 5175 -1025 5184 -961
rect 5116 -1035 5162 -1025
rect 5966 -1072 6012 -851
rect 387 -1076 6012 -1072
rect 387 -1110 403 -1076
rect 437 -1110 6012 -1076
rect 387 -1114 6012 -1110
rect 387 -1116 453 -1114
rect 46 -1167 92 -1155
rect 46 -1227 52 -1167
rect 86 -1227 92 -1167
rect 46 -1267 92 -1227
rect 120 -1167 210 -1155
rect 120 -1171 148 -1167
rect 182 -1171 210 -1167
rect 120 -1223 139 -1171
rect 191 -1223 210 -1171
rect 120 -1227 148 -1223
rect 182 -1227 210 -1223
rect 120 -1239 210 -1227
rect 238 -1167 284 -1155
rect 238 -1227 244 -1167
rect 278 -1227 284 -1167
rect 238 -1267 284 -1227
rect 326 -1167 372 -1155
rect 887 -1163 933 -1152
rect 326 -1227 332 -1167
rect 366 -1227 372 -1167
rect 326 -1239 372 -1227
rect 864 -1227 871 -1163
rect 935 -1227 943 -1163
rect 864 -1228 943 -1227
rect 994 -1164 1040 -1114
rect 1101 -1163 1147 -1152
rect 2099 -1163 2145 -1152
rect 994 -1224 1000 -1164
rect 1034 -1224 1040 -1164
rect 887 -1236 933 -1228
rect 994 -1236 1040 -1224
rect 1091 -1227 1099 -1163
rect 1163 -1227 1170 -1163
rect 1091 -1228 1170 -1227
rect 2076 -1227 2083 -1163
rect 2147 -1227 2155 -1163
rect 2076 -1228 2155 -1227
rect 2208 -1164 2254 -1114
rect 2313 -1163 2359 -1152
rect 3311 -1163 3357 -1152
rect 2208 -1224 2214 -1164
rect 2248 -1224 2254 -1164
rect 1101 -1236 1147 -1228
rect 2099 -1236 2145 -1228
rect 2208 -1236 2254 -1224
rect 2303 -1227 2311 -1163
rect 2375 -1227 2382 -1163
rect 2303 -1228 2382 -1227
rect 3288 -1227 3295 -1163
rect 3359 -1227 3367 -1163
rect 3288 -1228 3367 -1227
rect 3421 -1164 3467 -1114
rect 3525 -1163 3571 -1152
rect 4523 -1163 4569 -1152
rect 3421 -1224 3427 -1164
rect 3461 -1224 3467 -1164
rect 2313 -1236 2359 -1228
rect 3311 -1236 3357 -1228
rect 3421 -1236 3467 -1224
rect 3515 -1227 3523 -1163
rect 3587 -1227 3594 -1163
rect 3515 -1228 3594 -1227
rect 4500 -1227 4507 -1163
rect 4571 -1227 4579 -1163
rect 4500 -1228 4579 -1227
rect 4632 -1164 4678 -1114
rect 4737 -1163 4783 -1152
rect 4632 -1224 4638 -1164
rect 4672 -1224 4678 -1164
rect 3525 -1236 3571 -1228
rect 4523 -1236 4569 -1228
rect 4632 -1236 4678 -1224
rect 4727 -1227 4735 -1163
rect 4799 -1227 4806 -1163
rect 4727 -1228 4806 -1227
rect 5381 -1164 5427 -1114
rect 5469 -1160 5515 -1149
rect 5381 -1224 5387 -1164
rect 5421 -1224 5427 -1164
rect 4737 -1236 4783 -1228
rect 5381 -1236 5427 -1224
rect 5459 -1224 5467 -1160
rect 5531 -1224 5538 -1160
rect 5459 -1225 5538 -1224
rect 5469 -1233 5515 -1225
rect 46 -1296 284 -1267
rect 5419 -1276 5477 -1274
rect 5866 -1276 5915 -1272
rect 4900 -1277 5346 -1276
rect 5419 -1277 5915 -1276
rect 925 -1283 5346 -1277
rect 238 -1305 284 -1296
rect 238 -1365 244 -1305
rect 278 -1365 284 -1305
rect 238 -1377 284 -1365
rect 326 -1305 372 -1293
rect 326 -1365 332 -1305
rect 366 -1365 372 -1305
rect 925 -1317 937 -1283
rect 971 -1317 1063 -1283
rect 1097 -1317 2149 -1283
rect 2183 -1317 2275 -1283
rect 2309 -1317 3361 -1283
rect 3395 -1317 3487 -1283
rect 3521 -1317 4573 -1283
rect 4607 -1317 4699 -1283
rect 4733 -1317 5346 -1283
rect 925 -1323 5346 -1317
rect 5414 -1280 5915 -1277
rect 5414 -1314 5431 -1280
rect 5465 -1285 5915 -1280
rect 5465 -1314 5872 -1285
rect 5414 -1319 5872 -1314
rect 5906 -1319 5915 -1285
rect 5414 -1323 5915 -1319
rect 326 -1368 372 -1365
rect 326 -1414 373 -1368
rect 208 -1432 373 -1414
rect 5297 -1370 5346 -1323
rect 5866 -1331 5915 -1323
rect 5867 -1370 5916 -1365
rect 5297 -1378 5916 -1370
rect 5297 -1412 5873 -1378
rect 5907 -1412 5916 -1378
rect 5297 -1417 5916 -1412
rect 5867 -1424 5916 -1417
rect 208 -1484 227 -1432
rect 279 -1473 373 -1432
rect 279 -1484 298 -1473
rect 208 -1500 298 -1484
rect 5966 -1604 6012 -1114
rect 6050 -889 6108 -883
rect 6050 -923 6062 -889
rect 6096 -923 6108 -889
rect 6284 -917 6291 -865
rect 6343 -868 6349 -865
rect 6343 -914 6447 -868
rect 6947 -886 6953 -826
rect 6987 -886 6993 -826
rect 6947 -895 6993 -886
rect 6343 -916 6445 -914
rect 6343 -917 6349 -916
rect 6284 -918 6349 -917
rect 6050 -929 6108 -923
rect 6755 -924 6993 -895
rect 7035 -826 7081 -774
rect 7035 -886 7041 -826
rect 7075 -886 7081 -826
rect 7035 -898 7081 -886
rect 7634 -873 7693 259
rect 7994 216 8326 226
rect 7994 164 8012 216
rect 8064 164 8092 216
rect 8144 164 8172 216
rect 8224 164 8252 216
rect 8304 164 8326 216
rect 7994 158 8326 164
rect 8491 -873 8549 487
rect 8596 216 8928 226
rect 8596 164 8618 216
rect 8670 164 8698 216
rect 8750 164 8778 216
rect 8830 164 8858 216
rect 8910 164 8928 216
rect 8596 158 8928 164
rect 9332 216 9664 226
rect 9332 164 9350 216
rect 9402 164 9430 216
rect 9482 164 9510 216
rect 9562 164 9590 216
rect 9642 164 9664 216
rect 9332 158 9664 164
rect 9934 216 10266 226
rect 9934 164 9956 216
rect 10008 164 10036 216
rect 10088 164 10116 216
rect 10168 164 10196 216
rect 10248 164 10266 216
rect 9934 158 10266 164
rect 10544 216 10876 226
rect 10544 164 10562 216
rect 10614 164 10642 216
rect 10694 164 10722 216
rect 10774 164 10802 216
rect 10854 164 10876 216
rect 10544 158 10876 164
rect 10917 -873 10975 543
rect 11146 216 11478 226
rect 11146 164 11168 216
rect 11220 164 11248 216
rect 11300 164 11328 216
rect 11380 164 11408 216
rect 11460 164 11478 216
rect 11146 158 11478 164
rect 11878 216 12210 226
rect 11878 164 11900 216
rect 11952 164 11980 216
rect 12032 164 12060 216
rect 12112 164 12140 216
rect 12192 164 12210 216
rect 11878 158 12210 164
rect 12663 219 12770 235
rect 12663 167 12682 219
rect 12734 167 12770 219
rect 12663 151 12691 167
rect 12685 127 12691 151
rect 12725 151 12770 167
rect 12845 187 12891 199
rect 12725 127 12731 151
rect 12685 115 12731 127
rect 12845 127 12851 187
rect 12885 127 12891 187
rect 12685 49 12731 61
rect 12685 -11 12691 49
rect 12725 -11 12731 49
rect 12685 -89 12731 -11
rect 12845 49 12891 127
rect 12845 -11 12851 49
rect 12885 -11 12891 49
rect 12845 -23 12891 -11
rect 12685 -149 12691 -89
rect 12725 -149 12731 -89
rect 12685 -161 12731 -149
rect 12845 -89 12891 -77
rect 12845 -149 12851 -89
rect 12885 -149 12891 -89
rect 12685 -227 12731 -215
rect 12685 -287 12691 -227
rect 12725 -287 12731 -227
rect 12685 -365 12731 -287
rect 12845 -227 12891 -149
rect 12845 -287 12851 -227
rect 12885 -287 12891 -227
rect 12845 -299 12891 -287
rect 12685 -425 12691 -365
rect 12725 -425 12731 -365
rect 12685 -437 12731 -425
rect 12845 -365 12891 -353
rect 12845 -425 12851 -365
rect 12885 -425 12891 -365
rect 12685 -503 12731 -491
rect 12685 -563 12691 -503
rect 12725 -563 12731 -503
rect 12685 -641 12731 -563
rect 12845 -503 12891 -425
rect 12845 -563 12851 -503
rect 12885 -563 12891 -503
rect 12845 -575 12891 -563
rect 12685 -701 12691 -641
rect 12725 -701 12731 -641
rect 12685 -713 12731 -701
rect 12845 -641 12891 -629
rect 12845 -701 12851 -641
rect 12885 -701 12891 -641
rect 12675 -779 12731 -767
rect 12675 -839 12691 -779
rect 12725 -839 12731 -779
rect 12675 -851 12731 -839
rect 12845 -779 12891 -701
rect 12845 -839 12851 -779
rect 12885 -839 12891 -779
rect 12845 -851 12891 -839
rect 11773 -868 11831 -863
rect 12506 -865 12571 -864
rect 12506 -868 12512 -865
rect 7634 -879 7695 -873
rect 7634 -913 7649 -879
rect 7683 -913 7695 -879
rect 7634 -919 7695 -913
rect 8367 -879 8551 -873
rect 8367 -913 8383 -879
rect 8417 -913 8505 -879
rect 8539 -913 8551 -879
rect 8367 -919 8551 -913
rect 9705 -879 11101 -873
rect 9705 -913 9721 -879
rect 9755 -913 9843 -879
rect 9877 -913 10933 -879
rect 10967 -913 11055 -879
rect 11089 -913 11101 -879
rect 11773 -879 12512 -868
rect 11773 -898 11787 -879
rect 9705 -919 11101 -913
rect 11775 -913 11787 -898
rect 11821 -913 12512 -879
rect 11775 -915 12512 -913
rect 11775 -919 11833 -915
rect 12506 -917 12512 -915
rect 12564 -917 12571 -865
rect 7634 -922 7693 -919
rect 6050 -1070 6098 -929
rect 6755 -964 6801 -924
rect 6755 -1024 6761 -964
rect 6795 -1024 6801 -964
rect 6755 -1036 6801 -1024
rect 6829 -964 6919 -952
rect 6829 -968 6857 -964
rect 6891 -968 6919 -964
rect 6829 -1020 6848 -968
rect 6900 -1020 6919 -968
rect 6829 -1024 6857 -1020
rect 6891 -1024 6919 -1020
rect 6829 -1036 6919 -1024
rect 6947 -964 6993 -924
rect 6947 -1024 6953 -964
rect 6987 -1024 6993 -964
rect 6947 -1036 6993 -1024
rect 7035 -964 7081 -952
rect 7599 -960 7645 -951
rect 7035 -1024 7041 -964
rect 7075 -1024 7081 -964
rect 7035 -1036 7081 -1024
rect 7577 -961 7659 -960
rect 7577 -1025 7586 -961
rect 7650 -1025 7659 -961
rect 7688 -963 7734 -951
rect 8333 -960 8379 -951
rect 7688 -1023 7694 -963
rect 7728 -1023 7734 -963
rect 7599 -1035 7645 -1025
rect 6708 -1070 6951 -1068
rect 6050 -1074 6951 -1070
rect 6050 -1108 6905 -1074
rect 6939 -1078 6951 -1074
rect 7035 -1078 7063 -1036
rect 6939 -1107 7063 -1078
rect 6939 -1108 6951 -1107
rect 6050 -1114 6951 -1108
rect 6050 -1117 6770 -1114
rect 6050 -1517 6098 -1117
rect 7035 -1155 7063 -1107
rect 7096 -1072 7158 -1070
rect 7688 -1072 7734 -1023
rect 8311 -961 8393 -960
rect 8311 -1025 8320 -961
rect 8384 -1025 8393 -961
rect 8435 -963 8481 -951
rect 8543 -960 8589 -951
rect 9671 -960 9717 -951
rect 8435 -1023 8441 -963
rect 8475 -1023 8481 -963
rect 8333 -1035 8379 -1025
rect 8435 -1072 8481 -1023
rect 8529 -961 8611 -960
rect 8529 -1025 8538 -961
rect 8602 -1025 8611 -961
rect 9649 -961 9731 -960
rect 9649 -1025 9658 -961
rect 9722 -1025 9731 -961
rect 9775 -963 9821 -951
rect 9881 -960 9927 -951
rect 10883 -960 10929 -951
rect 9775 -1023 9781 -963
rect 9815 -1023 9821 -963
rect 8543 -1035 8589 -1025
rect 9671 -1035 9717 -1025
rect 9775 -1072 9821 -1023
rect 9867 -961 9949 -960
rect 9867 -1025 9876 -961
rect 9940 -1025 9949 -961
rect 10861 -961 10943 -960
rect 10861 -1025 10870 -961
rect 10934 -1025 10943 -961
rect 10986 -963 11032 -951
rect 11093 -960 11139 -951
rect 10986 -1023 10992 -963
rect 11026 -1023 11032 -963
rect 9881 -1035 9927 -1025
rect 10883 -1035 10929 -1025
rect 10986 -1072 11032 -1023
rect 11079 -961 11161 -960
rect 11079 -1025 11088 -961
rect 11152 -1025 11161 -961
rect 11735 -963 11781 -951
rect 11825 -960 11871 -951
rect 11735 -1023 11741 -963
rect 11775 -1023 11781 -963
rect 11093 -1035 11139 -1025
rect 11735 -1072 11781 -1023
rect 11811 -961 11893 -960
rect 11811 -1025 11820 -961
rect 11884 -1025 11893 -961
rect 11825 -1035 11871 -1025
rect 12675 -1072 12721 -851
rect 7096 -1076 12721 -1072
rect 7096 -1110 7112 -1076
rect 7146 -1110 12721 -1076
rect 7096 -1114 12721 -1110
rect 7096 -1116 7162 -1114
rect 6755 -1167 6801 -1155
rect 6233 -1208 6693 -1186
rect 6233 -1217 6295 -1208
rect 6347 -1217 6438 -1208
rect 6490 -1217 6558 -1208
rect 6610 -1217 6693 -1208
rect 6233 -1251 6262 -1217
rect 6347 -1251 6354 -1217
rect 6388 -1251 6438 -1217
rect 6490 -1251 6538 -1217
rect 6610 -1251 6630 -1217
rect 6664 -1251 6693 -1217
rect 6233 -1260 6295 -1251
rect 6347 -1260 6438 -1251
rect 6490 -1260 6558 -1251
rect 6610 -1260 6693 -1251
rect 6233 -1282 6693 -1260
rect 6755 -1227 6761 -1167
rect 6795 -1227 6801 -1167
rect 6755 -1267 6801 -1227
rect 6829 -1167 6919 -1155
rect 6829 -1171 6857 -1167
rect 6891 -1171 6919 -1167
rect 6829 -1223 6848 -1171
rect 6900 -1223 6919 -1171
rect 6829 -1227 6857 -1223
rect 6891 -1227 6919 -1223
rect 6829 -1239 6919 -1227
rect 6947 -1167 6993 -1155
rect 6947 -1227 6953 -1167
rect 6987 -1227 6993 -1167
rect 6947 -1267 6993 -1227
rect 7035 -1167 7081 -1155
rect 7596 -1163 7642 -1152
rect 7035 -1227 7041 -1167
rect 7075 -1227 7081 -1167
rect 7035 -1239 7081 -1227
rect 7573 -1227 7580 -1163
rect 7644 -1227 7652 -1163
rect 7573 -1228 7652 -1227
rect 7703 -1164 7749 -1114
rect 7810 -1163 7856 -1152
rect 8808 -1163 8854 -1152
rect 7703 -1224 7709 -1164
rect 7743 -1224 7749 -1164
rect 7596 -1236 7642 -1228
rect 7703 -1236 7749 -1224
rect 7800 -1227 7808 -1163
rect 7872 -1227 7879 -1163
rect 7800 -1228 7879 -1227
rect 8785 -1227 8792 -1163
rect 8856 -1227 8864 -1163
rect 8785 -1228 8864 -1227
rect 8917 -1164 8963 -1114
rect 9022 -1163 9068 -1152
rect 10020 -1163 10066 -1152
rect 8917 -1224 8923 -1164
rect 8957 -1224 8963 -1164
rect 7810 -1236 7856 -1228
rect 8808 -1236 8854 -1228
rect 8917 -1236 8963 -1224
rect 9012 -1227 9020 -1163
rect 9084 -1227 9091 -1163
rect 9012 -1228 9091 -1227
rect 9997 -1227 10004 -1163
rect 10068 -1227 10076 -1163
rect 9997 -1228 10076 -1227
rect 10130 -1164 10176 -1114
rect 10234 -1163 10280 -1152
rect 11232 -1163 11278 -1152
rect 10130 -1224 10136 -1164
rect 10170 -1224 10176 -1164
rect 9022 -1236 9068 -1228
rect 10020 -1236 10066 -1228
rect 10130 -1236 10176 -1224
rect 10224 -1227 10232 -1163
rect 10296 -1227 10303 -1163
rect 10224 -1228 10303 -1227
rect 11209 -1227 11216 -1163
rect 11280 -1227 11288 -1163
rect 11209 -1228 11288 -1227
rect 11341 -1164 11387 -1114
rect 11446 -1163 11492 -1152
rect 11341 -1224 11347 -1164
rect 11381 -1224 11387 -1164
rect 10234 -1236 10280 -1228
rect 11232 -1236 11278 -1228
rect 11341 -1236 11387 -1224
rect 11436 -1227 11444 -1163
rect 11508 -1227 11515 -1163
rect 11436 -1228 11515 -1227
rect 12090 -1164 12136 -1114
rect 12178 -1160 12224 -1149
rect 12090 -1224 12096 -1164
rect 12130 -1224 12136 -1164
rect 11446 -1236 11492 -1228
rect 12090 -1236 12136 -1224
rect 12168 -1224 12176 -1160
rect 12240 -1224 12247 -1160
rect 12168 -1225 12247 -1224
rect 12178 -1233 12224 -1225
rect 6755 -1296 6993 -1267
rect 12128 -1276 12186 -1274
rect 12575 -1276 12624 -1272
rect 11609 -1277 12055 -1276
rect 12128 -1277 12624 -1276
rect 7634 -1283 12055 -1277
rect 6947 -1305 6993 -1296
rect 6126 -1360 6175 -1347
rect 6126 -1394 6132 -1360
rect 6166 -1384 6175 -1360
rect 6947 -1365 6953 -1305
rect 6987 -1365 6993 -1305
rect 6947 -1377 6993 -1365
rect 7035 -1305 7081 -1293
rect 7035 -1365 7041 -1305
rect 7075 -1365 7081 -1305
rect 7634 -1317 7646 -1283
rect 7680 -1317 7772 -1283
rect 7806 -1317 8858 -1283
rect 8892 -1317 8984 -1283
rect 9018 -1317 10070 -1283
rect 10104 -1317 10196 -1283
rect 10230 -1317 11282 -1283
rect 11316 -1317 11408 -1283
rect 11442 -1317 12055 -1283
rect 7634 -1323 12055 -1317
rect 12123 -1280 12624 -1277
rect 12123 -1314 12140 -1280
rect 12174 -1285 12624 -1280
rect 12174 -1314 12581 -1285
rect 12123 -1319 12581 -1314
rect 12615 -1319 12624 -1285
rect 12123 -1323 12624 -1319
rect 7035 -1368 7081 -1365
rect 6166 -1394 6269 -1384
rect 6126 -1412 6269 -1394
rect 6164 -1453 6213 -1440
rect 6164 -1487 6170 -1453
rect 6204 -1487 6213 -1453
rect 6164 -1499 6213 -1487
rect 6050 -1523 6119 -1517
rect 6050 -1557 6073 -1523
rect 6107 -1557 6119 -1523
rect 6050 -1563 6119 -1557
rect 5966 -1616 6069 -1604
rect 126 -1674 216 -1658
rect 126 -1726 145 -1674
rect 197 -1726 216 -1674
rect 5966 -1676 6029 -1616
rect 6063 -1676 6069 -1616
rect 5966 -1688 6069 -1676
rect 6111 -1616 6157 -1604
rect 6111 -1676 6117 -1616
rect 6151 -1676 6157 -1616
rect 6185 -1631 6213 -1499
rect 6241 -1556 6269 -1412
rect 7035 -1414 7082 -1368
rect 6917 -1432 7082 -1414
rect 12006 -1370 12055 -1323
rect 12575 -1331 12624 -1323
rect 12576 -1370 12625 -1365
rect 12006 -1378 12625 -1370
rect 12006 -1412 12582 -1378
rect 12616 -1412 12625 -1378
rect 12006 -1417 12625 -1412
rect 12576 -1424 12625 -1417
rect 6297 -1443 6363 -1442
rect 6297 -1495 6303 -1443
rect 6355 -1495 6363 -1443
rect 6572 -1450 6626 -1446
rect 6571 -1453 6626 -1450
rect 6571 -1487 6583 -1453
rect 6617 -1487 6755 -1453
rect 6917 -1484 6936 -1432
rect 6988 -1473 7082 -1432
rect 6988 -1484 7007 -1473
rect 6571 -1490 6626 -1487
rect 6571 -1494 6625 -1490
rect 6297 -1497 6363 -1495
rect 6917 -1500 7007 -1484
rect 6241 -1563 6443 -1556
rect 6241 -1584 6393 -1563
rect 6376 -1597 6393 -1584
rect 6427 -1597 6443 -1563
rect 6376 -1603 6443 -1597
rect 12675 -1604 12721 -1114
rect 12759 -889 12817 -883
rect 12759 -923 12771 -889
rect 12805 -923 12817 -889
rect 12993 -917 13000 -865
rect 13052 -868 13058 -865
rect 13052 -914 13156 -868
rect 13052 -916 13154 -914
rect 13052 -917 13058 -916
rect 12993 -918 13058 -917
rect 12759 -929 12817 -923
rect 12759 -1070 12807 -929
rect 13446 -1070 13492 2389
rect 12759 -1117 13492 -1070
rect 12759 -1517 12807 -1117
rect 12942 -1208 13402 -1186
rect 12942 -1217 13004 -1208
rect 13056 -1217 13147 -1208
rect 13199 -1217 13267 -1208
rect 13319 -1217 13402 -1208
rect 12942 -1251 12971 -1217
rect 13056 -1251 13063 -1217
rect 13097 -1251 13147 -1217
rect 13199 -1251 13247 -1217
rect 13319 -1251 13339 -1217
rect 13373 -1251 13402 -1217
rect 12942 -1260 13004 -1251
rect 13056 -1260 13147 -1251
rect 13199 -1260 13267 -1251
rect 13319 -1260 13402 -1251
rect 12942 -1282 13402 -1260
rect 12835 -1360 12884 -1347
rect 12835 -1394 12841 -1360
rect 12875 -1384 12884 -1360
rect 12875 -1394 12978 -1384
rect 12835 -1412 12978 -1394
rect 12873 -1453 12922 -1440
rect 12873 -1487 12879 -1453
rect 12913 -1487 12922 -1453
rect 12873 -1499 12922 -1487
rect 12759 -1523 12828 -1517
rect 12759 -1557 12782 -1523
rect 12816 -1557 12828 -1523
rect 12759 -1563 12828 -1557
rect 6490 -1618 6548 -1611
rect 6490 -1631 6502 -1618
rect 6185 -1652 6502 -1631
rect 6536 -1652 6548 -1618
rect 6185 -1659 6548 -1652
rect 12675 -1616 12778 -1604
rect 126 -1742 216 -1726
rect 6023 -1754 6069 -1742
rect 6023 -1814 6029 -1754
rect 6063 -1814 6069 -1754
rect 125 -1831 215 -1815
rect 125 -1883 144 -1831
rect 196 -1883 215 -1831
rect 125 -1899 215 -1883
rect 6023 -1892 6069 -1814
rect 6111 -1754 6157 -1676
rect 6835 -1674 6925 -1658
rect 6835 -1726 6854 -1674
rect 6906 -1726 6925 -1674
rect 12675 -1676 12738 -1616
rect 12772 -1676 12778 -1616
rect 12675 -1688 12778 -1676
rect 12820 -1616 12866 -1604
rect 12820 -1676 12826 -1616
rect 12860 -1676 12866 -1616
rect 12894 -1631 12922 -1499
rect 12950 -1556 12978 -1412
rect 13006 -1443 13072 -1442
rect 13006 -1495 13012 -1443
rect 13064 -1495 13072 -1443
rect 13281 -1450 13335 -1446
rect 13280 -1453 13335 -1450
rect 13280 -1487 13292 -1453
rect 13326 -1487 13464 -1453
rect 13280 -1490 13335 -1487
rect 13280 -1494 13334 -1490
rect 13006 -1497 13072 -1495
rect 12950 -1563 13152 -1556
rect 12950 -1584 13102 -1563
rect 13085 -1597 13102 -1584
rect 13136 -1597 13152 -1563
rect 13085 -1603 13152 -1597
rect 13199 -1618 13257 -1611
rect 13199 -1631 13211 -1618
rect 12894 -1652 13211 -1631
rect 13245 -1652 13257 -1618
rect 12894 -1659 13257 -1652
rect 6111 -1814 6117 -1754
rect 6151 -1814 6157 -1754
rect 6111 -1826 6157 -1814
rect 6233 -1753 6693 -1730
rect 6835 -1742 6925 -1726
rect 6233 -1754 6445 -1753
rect 6233 -1761 6301 -1754
rect 6233 -1795 6262 -1761
rect 6296 -1795 6301 -1761
rect 6233 -1806 6301 -1795
rect 6353 -1761 6445 -1754
rect 6497 -1754 6693 -1753
rect 6497 -1761 6576 -1754
rect 6353 -1795 6354 -1761
rect 6388 -1795 6445 -1761
rect 6497 -1795 6538 -1761
rect 6572 -1795 6576 -1761
rect 6353 -1805 6445 -1795
rect 6497 -1805 6576 -1795
rect 6353 -1806 6576 -1805
rect 6628 -1761 6693 -1754
rect 6628 -1795 6630 -1761
rect 6664 -1795 6693 -1761
rect 6628 -1806 6693 -1795
rect 6233 -1826 6693 -1806
rect 12732 -1754 12778 -1742
rect 12732 -1814 12738 -1754
rect 12772 -1814 12778 -1754
rect 6834 -1831 6924 -1815
rect 6023 -1952 6029 -1892
rect 6063 -1952 6069 -1892
rect 6023 -1964 6069 -1952
rect 6111 -1892 6157 -1880
rect 6834 -1883 6853 -1831
rect 6905 -1883 6924 -1831
rect 6111 -1952 6117 -1892
rect 6151 -1952 6157 -1892
rect 125 -2001 215 -1985
rect 125 -2053 144 -2001
rect 196 -2053 215 -2001
rect 125 -2069 215 -2053
rect 6023 -2030 6069 -2018
rect 6023 -2090 6029 -2030
rect 6063 -2090 6069 -2030
rect 126 -2153 216 -2137
rect 126 -2205 145 -2153
rect 197 -2205 216 -2153
rect 126 -2221 216 -2205
rect 6023 -2168 6069 -2090
rect 6111 -2030 6157 -1952
rect 6412 -1903 6502 -1887
rect 6834 -1899 6924 -1883
rect 12732 -1892 12778 -1814
rect 12820 -1754 12866 -1676
rect 12820 -1814 12826 -1754
rect 12860 -1814 12866 -1754
rect 12820 -1826 12866 -1814
rect 12942 -1753 13402 -1730
rect 12942 -1754 13154 -1753
rect 12942 -1761 13010 -1754
rect 12942 -1795 12971 -1761
rect 13005 -1795 13010 -1761
rect 12942 -1806 13010 -1795
rect 13062 -1761 13154 -1754
rect 13206 -1754 13402 -1753
rect 13206 -1761 13285 -1754
rect 13062 -1795 13063 -1761
rect 13097 -1795 13154 -1761
rect 13206 -1795 13247 -1761
rect 13281 -1795 13285 -1761
rect 13062 -1805 13154 -1795
rect 13206 -1805 13285 -1795
rect 13062 -1806 13285 -1805
rect 13337 -1761 13402 -1754
rect 13337 -1795 13339 -1761
rect 13373 -1795 13402 -1761
rect 13337 -1806 13402 -1795
rect 12942 -1826 13402 -1806
rect 6412 -1955 6431 -1903
rect 6483 -1955 6502 -1903
rect 6412 -1971 6502 -1955
rect 12732 -1952 12738 -1892
rect 12772 -1952 12778 -1892
rect 12732 -1964 12778 -1952
rect 12820 -1892 12866 -1880
rect 12820 -1952 12826 -1892
rect 12860 -1952 12866 -1892
rect 6111 -2090 6117 -2030
rect 6151 -2090 6157 -2030
rect 6834 -2001 6924 -1985
rect 6834 -2053 6853 -2001
rect 6905 -2053 6924 -2001
rect 6834 -2069 6924 -2053
rect 12732 -2030 12778 -2018
rect 6111 -2102 6157 -2090
rect 6412 -2099 6502 -2083
rect 6412 -2151 6431 -2099
rect 6483 -2151 6502 -2099
rect 12732 -2090 12738 -2030
rect 12772 -2090 12778 -2030
rect 6023 -2228 6029 -2168
rect 6063 -2228 6069 -2168
rect 6023 -2240 6069 -2228
rect 6111 -2168 6157 -2156
rect 6412 -2167 6502 -2151
rect 6835 -2153 6925 -2137
rect 6111 -2228 6117 -2168
rect 6151 -2228 6157 -2168
rect 6835 -2205 6854 -2153
rect 6906 -2205 6925 -2153
rect 6835 -2221 6925 -2205
rect 12732 -2168 12778 -2090
rect 12820 -2030 12866 -1952
rect 12820 -2090 12826 -2030
rect 12860 -2090 12866 -2030
rect 12820 -2102 12866 -2090
rect 131 -2297 221 -2281
rect 131 -2349 150 -2297
rect 202 -2349 221 -2297
rect 6023 -2306 6069 -2294
rect 6023 -2312 6029 -2306
rect 5995 -2342 6029 -2312
rect 131 -2365 221 -2349
rect 381 -2353 5289 -2345
rect 381 -2405 489 -2353
rect 541 -2405 569 -2353
rect 621 -2405 649 -2353
rect 701 -2405 729 -2353
rect 781 -2405 809 -2353
rect 861 -2405 889 -2353
rect 941 -2405 1093 -2353
rect 1145 -2405 1173 -2353
rect 1225 -2405 1253 -2353
rect 1305 -2405 1333 -2353
rect 1385 -2405 1413 -2353
rect 1465 -2405 1493 -2353
rect 1545 -2405 1701 -2353
rect 1753 -2405 1781 -2353
rect 1833 -2405 1861 -2353
rect 1913 -2405 1941 -2353
rect 1993 -2405 2021 -2353
rect 2073 -2405 2101 -2353
rect 2153 -2405 2305 -2353
rect 2357 -2405 2385 -2353
rect 2437 -2405 2465 -2353
rect 2517 -2405 2545 -2353
rect 2597 -2405 2625 -2353
rect 2677 -2405 2705 -2353
rect 2757 -2405 2913 -2353
rect 2965 -2405 2993 -2353
rect 3045 -2405 3073 -2353
rect 3125 -2405 3153 -2353
rect 3205 -2405 3233 -2353
rect 3285 -2405 3313 -2353
rect 3365 -2405 3517 -2353
rect 3569 -2405 3597 -2353
rect 3649 -2405 3677 -2353
rect 3729 -2405 3757 -2353
rect 3809 -2405 3837 -2353
rect 3889 -2405 3917 -2353
rect 3969 -2405 4125 -2353
rect 4177 -2405 4205 -2353
rect 4257 -2405 4285 -2353
rect 4337 -2405 4365 -2353
rect 4417 -2405 4445 -2353
rect 4497 -2405 4525 -2353
rect 4577 -2405 4729 -2353
rect 4781 -2405 4809 -2353
rect 4861 -2405 4889 -2353
rect 4941 -2405 4969 -2353
rect 5021 -2405 5049 -2353
rect 5101 -2405 5129 -2353
rect 5181 -2405 5289 -2353
rect 381 -2411 5289 -2405
rect 5351 -2350 6029 -2342
rect 5351 -2402 5461 -2350
rect 5513 -2402 5541 -2350
rect 5593 -2402 5621 -2350
rect 5673 -2402 5701 -2350
rect 5753 -2402 5781 -2350
rect 5833 -2402 5861 -2350
rect 5913 -2359 6029 -2350
rect 5913 -2402 5959 -2359
rect 5351 -2408 5959 -2402
rect 5940 -2411 5959 -2408
rect 6011 -2366 6029 -2359
rect 6063 -2366 6069 -2306
rect 6011 -2378 6069 -2366
rect 6111 -2306 6157 -2228
rect 12732 -2228 12738 -2168
rect 12772 -2228 12778 -2168
rect 12732 -2240 12778 -2228
rect 12820 -2168 12866 -2156
rect 12820 -2228 12826 -2168
rect 12860 -2228 12866 -2168
rect 6111 -2366 6117 -2306
rect 6151 -2366 6157 -2306
rect 6412 -2274 6502 -2258
rect 6412 -2326 6431 -2274
rect 6483 -2326 6502 -2274
rect 6412 -2342 6502 -2326
rect 6840 -2297 6930 -2281
rect 6840 -2349 6859 -2297
rect 6911 -2349 6930 -2297
rect 12732 -2306 12778 -2294
rect 12732 -2312 12738 -2306
rect 12704 -2342 12738 -2312
rect 6840 -2365 6930 -2349
rect 7090 -2353 11998 -2345
rect 6111 -2378 6157 -2366
rect 6011 -2400 6048 -2378
rect 6011 -2411 6030 -2400
rect 7090 -2405 7198 -2353
rect 7250 -2405 7278 -2353
rect 7330 -2405 7358 -2353
rect 7410 -2405 7438 -2353
rect 7490 -2405 7518 -2353
rect 7570 -2405 7598 -2353
rect 7650 -2405 7802 -2353
rect 7854 -2405 7882 -2353
rect 7934 -2405 7962 -2353
rect 8014 -2405 8042 -2353
rect 8094 -2405 8122 -2353
rect 8174 -2405 8202 -2353
rect 8254 -2405 8410 -2353
rect 8462 -2405 8490 -2353
rect 8542 -2405 8570 -2353
rect 8622 -2405 8650 -2353
rect 8702 -2405 8730 -2353
rect 8782 -2405 8810 -2353
rect 8862 -2405 9014 -2353
rect 9066 -2405 9094 -2353
rect 9146 -2405 9174 -2353
rect 9226 -2405 9254 -2353
rect 9306 -2405 9334 -2353
rect 9386 -2405 9414 -2353
rect 9466 -2405 9622 -2353
rect 9674 -2405 9702 -2353
rect 9754 -2405 9782 -2353
rect 9834 -2405 9862 -2353
rect 9914 -2405 9942 -2353
rect 9994 -2405 10022 -2353
rect 10074 -2405 10226 -2353
rect 10278 -2405 10306 -2353
rect 10358 -2405 10386 -2353
rect 10438 -2405 10466 -2353
rect 10518 -2405 10546 -2353
rect 10598 -2405 10626 -2353
rect 10678 -2405 10834 -2353
rect 10886 -2405 10914 -2353
rect 10966 -2405 10994 -2353
rect 11046 -2405 11074 -2353
rect 11126 -2405 11154 -2353
rect 11206 -2405 11234 -2353
rect 11286 -2405 11438 -2353
rect 11490 -2405 11518 -2353
rect 11570 -2405 11598 -2353
rect 11650 -2405 11678 -2353
rect 11730 -2405 11758 -2353
rect 11810 -2405 11838 -2353
rect 11890 -2405 11998 -2353
rect 7090 -2411 11998 -2405
rect 12060 -2350 12738 -2342
rect 12060 -2402 12170 -2350
rect 12222 -2402 12250 -2350
rect 12302 -2402 12330 -2350
rect 12382 -2402 12410 -2350
rect 12462 -2402 12490 -2350
rect 12542 -2402 12570 -2350
rect 12622 -2359 12738 -2350
rect 12622 -2402 12668 -2359
rect 12060 -2408 12668 -2402
rect 12649 -2411 12668 -2408
rect 12720 -2366 12738 -2359
rect 12772 -2366 12778 -2306
rect 12720 -2378 12778 -2366
rect 12820 -2306 12866 -2228
rect 12820 -2366 12826 -2306
rect 12860 -2366 12866 -2306
rect 12820 -2378 12866 -2366
rect 12720 -2400 12757 -2378
rect 12720 -2411 12739 -2400
rect 5940 -2427 6030 -2411
rect 12649 -2427 12739 -2411
<< via1 >>
rect 744 3680 796 3732
rect 842 3711 894 3723
rect 842 3677 852 3711
rect 852 3677 886 3711
rect 886 3677 894 3711
rect 842 3671 894 3677
rect 922 3711 974 3723
rect 922 3677 932 3711
rect 932 3677 966 3711
rect 966 3677 974 3711
rect 922 3671 974 3677
rect 1002 3711 1054 3723
rect 1002 3677 1012 3711
rect 1012 3677 1046 3711
rect 1046 3677 1054 3711
rect 1002 3671 1054 3677
rect 1082 3711 1134 3723
rect 1082 3677 1092 3711
rect 1092 3677 1126 3711
rect 1126 3677 1134 3711
rect 1082 3671 1134 3677
rect 1162 3711 1214 3723
rect 1162 3677 1172 3711
rect 1172 3677 1206 3711
rect 1206 3677 1214 3711
rect 1162 3671 1214 3677
rect 1242 3711 1294 3723
rect 1242 3677 1252 3711
rect 1252 3677 1286 3711
rect 1286 3677 1294 3711
rect 1242 3671 1294 3677
rect 1574 3714 1626 3726
rect 1574 3680 1584 3714
rect 1584 3680 1618 3714
rect 1618 3680 1626 3714
rect 1574 3674 1626 3680
rect 1654 3714 1706 3726
rect 1654 3680 1664 3714
rect 1664 3680 1698 3714
rect 1698 3680 1706 3714
rect 1654 3674 1706 3680
rect 1734 3714 1786 3726
rect 1734 3680 1744 3714
rect 1744 3680 1778 3714
rect 1778 3680 1786 3714
rect 1734 3674 1786 3680
rect 1814 3714 1866 3726
rect 1814 3680 1824 3714
rect 1824 3680 1858 3714
rect 1858 3680 1866 3714
rect 1814 3674 1866 3680
rect 1894 3714 1946 3726
rect 1894 3680 1904 3714
rect 1904 3680 1938 3714
rect 1938 3680 1946 3714
rect 1894 3674 1946 3680
rect 1974 3714 2026 3726
rect 1974 3680 1984 3714
rect 1984 3680 2018 3714
rect 2018 3680 2026 3714
rect 1974 3674 2026 3680
rect 2178 3714 2230 3726
rect 2178 3680 2186 3714
rect 2186 3680 2220 3714
rect 2220 3680 2230 3714
rect 2178 3674 2230 3680
rect 2258 3714 2310 3726
rect 2258 3680 2266 3714
rect 2266 3680 2300 3714
rect 2300 3680 2310 3714
rect 2258 3674 2310 3680
rect 2338 3714 2390 3726
rect 2338 3680 2346 3714
rect 2346 3680 2380 3714
rect 2380 3680 2390 3714
rect 2338 3674 2390 3680
rect 2418 3714 2470 3726
rect 2418 3680 2426 3714
rect 2426 3680 2460 3714
rect 2460 3680 2470 3714
rect 2418 3674 2470 3680
rect 2498 3714 2550 3726
rect 2498 3680 2506 3714
rect 2506 3680 2540 3714
rect 2540 3680 2550 3714
rect 2498 3674 2550 3680
rect 2578 3714 2630 3726
rect 2578 3680 2586 3714
rect 2586 3680 2620 3714
rect 2620 3680 2630 3714
rect 2578 3674 2630 3680
rect 2786 3714 2838 3726
rect 2786 3680 2796 3714
rect 2796 3680 2830 3714
rect 2830 3680 2838 3714
rect 2786 3674 2838 3680
rect 2866 3714 2918 3726
rect 2866 3680 2876 3714
rect 2876 3680 2910 3714
rect 2910 3680 2918 3714
rect 2866 3674 2918 3680
rect 2946 3714 2998 3726
rect 2946 3680 2956 3714
rect 2956 3680 2990 3714
rect 2990 3680 2998 3714
rect 2946 3674 2998 3680
rect 3026 3714 3078 3726
rect 3026 3680 3036 3714
rect 3036 3680 3070 3714
rect 3070 3680 3078 3714
rect 3026 3674 3078 3680
rect 3106 3714 3158 3726
rect 3106 3680 3116 3714
rect 3116 3680 3150 3714
rect 3150 3680 3158 3714
rect 3106 3674 3158 3680
rect 3186 3714 3238 3726
rect 3186 3680 3196 3714
rect 3196 3680 3230 3714
rect 3230 3680 3238 3714
rect 3186 3674 3238 3680
rect 3390 3714 3442 3726
rect 3390 3680 3398 3714
rect 3398 3680 3432 3714
rect 3432 3680 3442 3714
rect 3390 3674 3442 3680
rect 3470 3714 3522 3726
rect 3470 3680 3478 3714
rect 3478 3680 3512 3714
rect 3512 3680 3522 3714
rect 3470 3674 3522 3680
rect 3550 3714 3602 3726
rect 3550 3680 3558 3714
rect 3558 3680 3592 3714
rect 3592 3680 3602 3714
rect 3550 3674 3602 3680
rect 3630 3714 3682 3726
rect 3630 3680 3638 3714
rect 3638 3680 3672 3714
rect 3672 3680 3682 3714
rect 3630 3674 3682 3680
rect 3710 3714 3762 3726
rect 3710 3680 3718 3714
rect 3718 3680 3752 3714
rect 3752 3680 3762 3714
rect 3710 3674 3762 3680
rect 3790 3714 3842 3726
rect 3790 3680 3798 3714
rect 3798 3680 3832 3714
rect 3832 3680 3842 3714
rect 3790 3674 3842 3680
rect 3998 3714 4050 3726
rect 3998 3680 4008 3714
rect 4008 3680 4042 3714
rect 4042 3680 4050 3714
rect 3998 3674 4050 3680
rect 4078 3714 4130 3726
rect 4078 3680 4088 3714
rect 4088 3680 4122 3714
rect 4122 3680 4130 3714
rect 4078 3674 4130 3680
rect 4158 3714 4210 3726
rect 4158 3680 4168 3714
rect 4168 3680 4202 3714
rect 4202 3680 4210 3714
rect 4158 3674 4210 3680
rect 4238 3714 4290 3726
rect 4238 3680 4248 3714
rect 4248 3680 4282 3714
rect 4282 3680 4290 3714
rect 4238 3674 4290 3680
rect 4318 3714 4370 3726
rect 4318 3680 4328 3714
rect 4328 3680 4362 3714
rect 4362 3680 4370 3714
rect 4318 3674 4370 3680
rect 4398 3714 4450 3726
rect 4398 3680 4408 3714
rect 4408 3680 4442 3714
rect 4442 3680 4450 3714
rect 4398 3674 4450 3680
rect 4602 3714 4654 3726
rect 4602 3680 4610 3714
rect 4610 3680 4644 3714
rect 4644 3680 4654 3714
rect 4602 3674 4654 3680
rect 4682 3714 4734 3726
rect 4682 3680 4690 3714
rect 4690 3680 4724 3714
rect 4724 3680 4734 3714
rect 4682 3674 4734 3680
rect 4762 3714 4814 3726
rect 4762 3680 4770 3714
rect 4770 3680 4804 3714
rect 4804 3680 4814 3714
rect 4762 3674 4814 3680
rect 4842 3714 4894 3726
rect 4842 3680 4850 3714
rect 4850 3680 4884 3714
rect 4884 3680 4894 3714
rect 4842 3674 4894 3680
rect 4922 3714 4974 3726
rect 4922 3680 4930 3714
rect 4930 3680 4964 3714
rect 4964 3680 4974 3714
rect 4922 3674 4974 3680
rect 5002 3714 5054 3726
rect 5002 3680 5010 3714
rect 5010 3680 5044 3714
rect 5044 3680 5054 3714
rect 5002 3674 5054 3680
rect 5210 3714 5262 3726
rect 5210 3680 5220 3714
rect 5220 3680 5254 3714
rect 5254 3680 5262 3714
rect 5210 3674 5262 3680
rect 5290 3714 5342 3726
rect 5290 3680 5300 3714
rect 5300 3680 5334 3714
rect 5334 3680 5342 3714
rect 5290 3674 5342 3680
rect 5370 3714 5422 3726
rect 5370 3680 5380 3714
rect 5380 3680 5414 3714
rect 5414 3680 5422 3714
rect 5370 3674 5422 3680
rect 5450 3714 5502 3726
rect 5450 3680 5460 3714
rect 5460 3680 5494 3714
rect 5494 3680 5502 3714
rect 5450 3674 5502 3680
rect 5530 3714 5582 3726
rect 5530 3680 5540 3714
rect 5540 3680 5574 3714
rect 5574 3680 5582 3714
rect 5530 3674 5582 3680
rect 5610 3714 5662 3726
rect 5610 3680 5620 3714
rect 5620 3680 5654 3714
rect 5654 3680 5662 3714
rect 5610 3674 5662 3680
rect 5814 3714 5866 3726
rect 5814 3680 5822 3714
rect 5822 3680 5856 3714
rect 5856 3680 5866 3714
rect 5814 3674 5866 3680
rect 5894 3714 5946 3726
rect 5894 3680 5902 3714
rect 5902 3680 5936 3714
rect 5936 3680 5946 3714
rect 5894 3674 5946 3680
rect 5974 3714 6026 3726
rect 5974 3680 5982 3714
rect 5982 3680 6016 3714
rect 6016 3680 6026 3714
rect 5974 3674 6026 3680
rect 6054 3714 6106 3726
rect 6054 3680 6062 3714
rect 6062 3680 6096 3714
rect 6096 3680 6106 3714
rect 6054 3674 6106 3680
rect 6134 3714 6186 3726
rect 6134 3680 6142 3714
rect 6142 3680 6176 3714
rect 6176 3680 6186 3714
rect 6134 3674 6186 3680
rect 6214 3714 6266 3726
rect 6214 3680 6222 3714
rect 6222 3680 6256 3714
rect 6256 3680 6266 3714
rect 6214 3674 6266 3680
rect 6553 3663 6605 3670
rect 6553 3629 6564 3663
rect 6564 3629 6598 3663
rect 6598 3629 6605 3663
rect 6553 3618 6605 3629
rect 7030 3666 7082 3673
rect 7030 3632 7041 3666
rect 7041 3632 7075 3666
rect 7075 3632 7082 3666
rect 7030 3621 7082 3632
rect 7453 3680 7505 3732
rect 7551 3711 7603 3723
rect 7551 3677 7561 3711
rect 7561 3677 7595 3711
rect 7595 3677 7603 3711
rect 7551 3671 7603 3677
rect 7631 3711 7683 3723
rect 7631 3677 7641 3711
rect 7641 3677 7675 3711
rect 7675 3677 7683 3711
rect 7631 3671 7683 3677
rect 7711 3711 7763 3723
rect 7711 3677 7721 3711
rect 7721 3677 7755 3711
rect 7755 3677 7763 3711
rect 7711 3671 7763 3677
rect 7791 3711 7843 3723
rect 7791 3677 7801 3711
rect 7801 3677 7835 3711
rect 7835 3677 7843 3711
rect 7791 3671 7843 3677
rect 7871 3711 7923 3723
rect 7871 3677 7881 3711
rect 7881 3677 7915 3711
rect 7915 3677 7923 3711
rect 7871 3671 7923 3677
rect 7951 3711 8003 3723
rect 7951 3677 7961 3711
rect 7961 3677 7995 3711
rect 7995 3677 8003 3711
rect 7951 3671 8003 3677
rect 8283 3714 8335 3726
rect 8283 3680 8293 3714
rect 8293 3680 8327 3714
rect 8327 3680 8335 3714
rect 8283 3674 8335 3680
rect 8363 3714 8415 3726
rect 8363 3680 8373 3714
rect 8373 3680 8407 3714
rect 8407 3680 8415 3714
rect 8363 3674 8415 3680
rect 8443 3714 8495 3726
rect 8443 3680 8453 3714
rect 8453 3680 8487 3714
rect 8487 3680 8495 3714
rect 8443 3674 8495 3680
rect 8523 3714 8575 3726
rect 8523 3680 8533 3714
rect 8533 3680 8567 3714
rect 8567 3680 8575 3714
rect 8523 3674 8575 3680
rect 8603 3714 8655 3726
rect 8603 3680 8613 3714
rect 8613 3680 8647 3714
rect 8647 3680 8655 3714
rect 8603 3674 8655 3680
rect 8683 3714 8735 3726
rect 8683 3680 8693 3714
rect 8693 3680 8727 3714
rect 8727 3680 8735 3714
rect 8683 3674 8735 3680
rect 8887 3714 8939 3726
rect 8887 3680 8895 3714
rect 8895 3680 8929 3714
rect 8929 3680 8939 3714
rect 8887 3674 8939 3680
rect 8967 3714 9019 3726
rect 8967 3680 8975 3714
rect 8975 3680 9009 3714
rect 9009 3680 9019 3714
rect 8967 3674 9019 3680
rect 9047 3714 9099 3726
rect 9047 3680 9055 3714
rect 9055 3680 9089 3714
rect 9089 3680 9099 3714
rect 9047 3674 9099 3680
rect 9127 3714 9179 3726
rect 9127 3680 9135 3714
rect 9135 3680 9169 3714
rect 9169 3680 9179 3714
rect 9127 3674 9179 3680
rect 9207 3714 9259 3726
rect 9207 3680 9215 3714
rect 9215 3680 9249 3714
rect 9249 3680 9259 3714
rect 9207 3674 9259 3680
rect 9287 3714 9339 3726
rect 9287 3680 9295 3714
rect 9295 3680 9329 3714
rect 9329 3680 9339 3714
rect 9287 3674 9339 3680
rect 9495 3714 9547 3726
rect 9495 3680 9505 3714
rect 9505 3680 9539 3714
rect 9539 3680 9547 3714
rect 9495 3674 9547 3680
rect 9575 3714 9627 3726
rect 9575 3680 9585 3714
rect 9585 3680 9619 3714
rect 9619 3680 9627 3714
rect 9575 3674 9627 3680
rect 9655 3714 9707 3726
rect 9655 3680 9665 3714
rect 9665 3680 9699 3714
rect 9699 3680 9707 3714
rect 9655 3674 9707 3680
rect 9735 3714 9787 3726
rect 9735 3680 9745 3714
rect 9745 3680 9779 3714
rect 9779 3680 9787 3714
rect 9735 3674 9787 3680
rect 9815 3714 9867 3726
rect 9815 3680 9825 3714
rect 9825 3680 9859 3714
rect 9859 3680 9867 3714
rect 9815 3674 9867 3680
rect 9895 3714 9947 3726
rect 9895 3680 9905 3714
rect 9905 3680 9939 3714
rect 9939 3680 9947 3714
rect 9895 3674 9947 3680
rect 10099 3714 10151 3726
rect 10099 3680 10107 3714
rect 10107 3680 10141 3714
rect 10141 3680 10151 3714
rect 10099 3674 10151 3680
rect 10179 3714 10231 3726
rect 10179 3680 10187 3714
rect 10187 3680 10221 3714
rect 10221 3680 10231 3714
rect 10179 3674 10231 3680
rect 10259 3714 10311 3726
rect 10259 3680 10267 3714
rect 10267 3680 10301 3714
rect 10301 3680 10311 3714
rect 10259 3674 10311 3680
rect 10339 3714 10391 3726
rect 10339 3680 10347 3714
rect 10347 3680 10381 3714
rect 10381 3680 10391 3714
rect 10339 3674 10391 3680
rect 10419 3714 10471 3726
rect 10419 3680 10427 3714
rect 10427 3680 10461 3714
rect 10461 3680 10471 3714
rect 10419 3674 10471 3680
rect 10499 3714 10551 3726
rect 10499 3680 10507 3714
rect 10507 3680 10541 3714
rect 10541 3680 10551 3714
rect 10499 3674 10551 3680
rect 10707 3714 10759 3726
rect 10707 3680 10717 3714
rect 10717 3680 10751 3714
rect 10751 3680 10759 3714
rect 10707 3674 10759 3680
rect 10787 3714 10839 3726
rect 10787 3680 10797 3714
rect 10797 3680 10831 3714
rect 10831 3680 10839 3714
rect 10787 3674 10839 3680
rect 10867 3714 10919 3726
rect 10867 3680 10877 3714
rect 10877 3680 10911 3714
rect 10911 3680 10919 3714
rect 10867 3674 10919 3680
rect 10947 3714 10999 3726
rect 10947 3680 10957 3714
rect 10957 3680 10991 3714
rect 10991 3680 10999 3714
rect 10947 3674 10999 3680
rect 11027 3714 11079 3726
rect 11027 3680 11037 3714
rect 11037 3680 11071 3714
rect 11071 3680 11079 3714
rect 11027 3674 11079 3680
rect 11107 3714 11159 3726
rect 11107 3680 11117 3714
rect 11117 3680 11151 3714
rect 11151 3680 11159 3714
rect 11107 3674 11159 3680
rect 11311 3714 11363 3726
rect 11311 3680 11319 3714
rect 11319 3680 11353 3714
rect 11353 3680 11363 3714
rect 11311 3674 11363 3680
rect 11391 3714 11443 3726
rect 11391 3680 11399 3714
rect 11399 3680 11433 3714
rect 11433 3680 11443 3714
rect 11391 3674 11443 3680
rect 11471 3714 11523 3726
rect 11471 3680 11479 3714
rect 11479 3680 11513 3714
rect 11513 3680 11523 3714
rect 11471 3674 11523 3680
rect 11551 3714 11603 3726
rect 11551 3680 11559 3714
rect 11559 3680 11593 3714
rect 11593 3680 11603 3714
rect 11551 3674 11603 3680
rect 11631 3714 11683 3726
rect 11631 3680 11639 3714
rect 11639 3680 11673 3714
rect 11673 3680 11683 3714
rect 11631 3674 11683 3680
rect 11711 3714 11763 3726
rect 11711 3680 11719 3714
rect 11719 3680 11753 3714
rect 11753 3680 11763 3714
rect 11711 3674 11763 3680
rect 11919 3714 11971 3726
rect 11919 3680 11929 3714
rect 11929 3680 11963 3714
rect 11963 3680 11971 3714
rect 11919 3674 11971 3680
rect 11999 3714 12051 3726
rect 11999 3680 12009 3714
rect 12009 3680 12043 3714
rect 12043 3680 12051 3714
rect 11999 3674 12051 3680
rect 12079 3714 12131 3726
rect 12079 3680 12089 3714
rect 12089 3680 12123 3714
rect 12123 3680 12131 3714
rect 12079 3674 12131 3680
rect 12159 3714 12211 3726
rect 12159 3680 12169 3714
rect 12169 3680 12203 3714
rect 12203 3680 12211 3714
rect 12159 3674 12211 3680
rect 12239 3714 12291 3726
rect 12239 3680 12249 3714
rect 12249 3680 12283 3714
rect 12283 3680 12291 3714
rect 12239 3674 12291 3680
rect 12319 3714 12371 3726
rect 12319 3680 12329 3714
rect 12329 3680 12363 3714
rect 12363 3680 12371 3714
rect 12319 3674 12371 3680
rect 12523 3714 12575 3726
rect 12523 3680 12531 3714
rect 12531 3680 12565 3714
rect 12565 3680 12575 3714
rect 12523 3674 12575 3680
rect 12603 3714 12655 3726
rect 12603 3680 12611 3714
rect 12611 3680 12645 3714
rect 12645 3680 12655 3714
rect 12603 3674 12655 3680
rect 12683 3714 12735 3726
rect 12683 3680 12691 3714
rect 12691 3680 12725 3714
rect 12725 3680 12735 3714
rect 12683 3674 12735 3680
rect 12763 3714 12815 3726
rect 12763 3680 12771 3714
rect 12771 3680 12805 3714
rect 12805 3680 12815 3714
rect 12763 3674 12815 3680
rect 12843 3714 12895 3726
rect 12843 3680 12851 3714
rect 12851 3680 12885 3714
rect 12885 3680 12895 3714
rect 12843 3674 12895 3680
rect 12923 3714 12975 3726
rect 12923 3680 12931 3714
rect 12931 3680 12965 3714
rect 12965 3680 12975 3714
rect 12923 3674 12975 3680
rect 13262 3663 13314 3670
rect 13262 3629 13273 3663
rect 13273 3629 13307 3663
rect 13307 3629 13314 3663
rect 13262 3618 13314 3629
rect 6558 3519 6610 3526
rect 6558 3485 6569 3519
rect 6569 3485 6603 3519
rect 6603 3485 6610 3519
rect 6558 3474 6610 3485
rect 7019 3494 7071 3501
rect 7019 3460 7030 3494
rect 7030 3460 7064 3494
rect 7064 3460 7071 3494
rect 7019 3449 7071 3460
rect 6559 3367 6611 3374
rect 6559 3333 6570 3367
rect 6570 3333 6604 3367
rect 6604 3333 6611 3367
rect 6559 3322 6611 3333
rect 7019 3302 7071 3309
rect 7019 3268 7030 3302
rect 7030 3268 7064 3302
rect 7064 3268 7071 3302
rect 7019 3257 7071 3268
rect 13267 3519 13319 3526
rect 13267 3485 13278 3519
rect 13278 3485 13312 3519
rect 13312 3485 13319 3519
rect 13267 3474 13319 3485
rect 13268 3367 13320 3374
rect 13268 3333 13279 3367
rect 13279 3333 13313 3367
rect 13313 3333 13320 3367
rect 13268 3322 13320 3333
rect 127 3075 179 3127
rect 258 3116 310 3126
rect 258 3082 275 3116
rect 275 3082 309 3116
rect 309 3082 310 3116
rect 258 3074 310 3082
rect 402 3075 454 3127
rect 6559 3197 6611 3204
rect 6559 3163 6570 3197
rect 6570 3163 6604 3197
rect 6604 3163 6611 3197
rect 6559 3152 6611 3163
rect 6836 3075 6888 3127
rect 6967 3116 7019 3126
rect 6967 3082 6984 3116
rect 6984 3082 7018 3116
rect 7018 3082 7019 3116
rect 6967 3074 7019 3082
rect 7111 3075 7163 3127
rect 400 2807 452 2816
rect 400 2773 412 2807
rect 412 2773 446 2807
rect 446 2773 452 2807
rect 400 2764 452 2773
rect 6558 3040 6610 3047
rect 6558 3006 6569 3040
rect 6569 3006 6603 3040
rect 6603 3006 6610 3040
rect 6558 2995 6610 3006
rect 13268 3197 13320 3204
rect 13268 3163 13279 3197
rect 13279 3163 13313 3197
rect 13313 3163 13320 3197
rect 13268 3152 13320 3163
rect 145 2572 197 2581
rect 265 2572 317 2581
rect 408 2572 460 2581
rect 145 2538 183 2572
rect 183 2538 197 2572
rect 265 2538 275 2572
rect 275 2538 309 2572
rect 309 2538 317 2572
rect 408 2538 459 2572
rect 459 2538 460 2572
rect 145 2529 197 2538
rect 265 2529 317 2538
rect 408 2529 460 2538
rect 412 2186 464 2238
rect 6476 2753 6528 2805
rect 7109 2807 7161 2816
rect 7109 2773 7121 2807
rect 7121 2773 7155 2807
rect 7155 2773 7161 2807
rect 7109 2764 7161 2773
rect 13267 3040 13319 3047
rect 13267 3006 13278 3040
rect 13278 3006 13312 3040
rect 13312 3006 13319 3040
rect 13267 2995 13319 3006
rect 1224 2542 1288 2545
rect 1224 2482 1246 2542
rect 1246 2482 1280 2542
rect 1280 2482 1288 2542
rect 1224 2481 1288 2482
rect 1956 2545 2020 2548
rect 1956 2485 1978 2545
rect 1978 2485 2012 2545
rect 2012 2485 2020 2545
rect 1956 2484 2020 2485
rect 2184 2545 2248 2548
rect 2184 2485 2192 2545
rect 2192 2485 2226 2545
rect 2226 2485 2248 2545
rect 2184 2484 2248 2485
rect 3168 2545 3232 2548
rect 3168 2485 3190 2545
rect 3190 2485 3224 2545
rect 3224 2485 3232 2545
rect 3168 2484 3232 2485
rect 3396 2545 3460 2548
rect 3396 2485 3404 2545
rect 3404 2485 3438 2545
rect 3438 2485 3460 2545
rect 3396 2484 3460 2485
rect 4380 2545 4444 2548
rect 4380 2485 4402 2545
rect 4402 2485 4436 2545
rect 4436 2485 4444 2545
rect 4380 2484 4444 2485
rect 4608 2545 4672 2548
rect 4608 2485 4616 2545
rect 4616 2485 4650 2545
rect 4650 2485 4672 2545
rect 4608 2484 4672 2485
rect 5592 2545 5656 2548
rect 5592 2485 5614 2545
rect 5614 2485 5648 2545
rect 5648 2485 5656 2545
rect 5592 2484 5656 2485
rect 5820 2545 5884 2548
rect 5820 2485 5828 2545
rect 5828 2485 5862 2545
rect 5862 2485 5884 2545
rect 5820 2484 5884 2485
rect 6564 2492 6573 2544
rect 6573 2492 6607 2544
rect 6607 2492 6616 2544
rect 6854 2572 6906 2581
rect 6974 2572 7026 2581
rect 7117 2572 7169 2581
rect 6854 2538 6892 2572
rect 6892 2538 6906 2572
rect 6974 2538 6984 2572
rect 6984 2538 7018 2572
rect 7018 2538 7026 2572
rect 7117 2538 7168 2572
rect 7168 2538 7169 2572
rect 6854 2529 6906 2538
rect 6974 2529 7026 2538
rect 7117 2529 7169 2538
rect 1580 2344 1644 2346
rect 1580 2284 1599 2344
rect 1599 2284 1633 2344
rect 1633 2284 1644 2344
rect 1580 2282 1644 2284
rect 2312 2344 2376 2346
rect 2312 2284 2331 2344
rect 2331 2284 2365 2344
rect 2365 2284 2376 2344
rect 2312 2282 2376 2284
rect 2530 2344 2594 2346
rect 2530 2284 2541 2344
rect 2541 2284 2575 2344
rect 2575 2284 2594 2344
rect 2530 2282 2594 2284
rect 3524 2344 3588 2346
rect 3524 2284 3543 2344
rect 3543 2284 3577 2344
rect 3577 2284 3588 2344
rect 3524 2282 3588 2284
rect 3742 2344 3806 2346
rect 3742 2284 3753 2344
rect 3753 2284 3787 2344
rect 3787 2284 3806 2344
rect 3742 2282 3806 2284
rect 4862 2344 4926 2346
rect 4862 2284 4881 2344
rect 4881 2284 4915 2344
rect 4915 2284 4926 2344
rect 4862 2282 4926 2284
rect 5080 2344 5144 2346
rect 5080 2284 5091 2344
rect 5091 2284 5125 2344
rect 5125 2284 5144 2344
rect 5080 2282 5144 2284
rect 5814 2344 5878 2346
rect 5814 2284 5825 2344
rect 5825 2284 5859 2344
rect 5859 2284 5878 2344
rect 5814 2282 5878 2284
rect 6564 2289 6573 2341
rect 6573 2289 6607 2341
rect 6607 2289 6616 2341
rect 900 2186 952 2238
rect 105 1649 163 1700
rect 163 1649 165 1700
rect 105 1644 165 1649
rect 730 1134 739 1154
rect 739 1134 773 1154
rect 773 1134 782 1154
rect 730 1102 782 1134
rect 1272 1147 1324 1157
rect 1272 1113 1280 1147
rect 1280 1113 1314 1147
rect 1314 1113 1324 1147
rect 1272 1105 1324 1113
rect 1352 1147 1404 1157
rect 1352 1113 1360 1147
rect 1360 1113 1394 1147
rect 1394 1113 1404 1147
rect 1352 1105 1404 1113
rect 1432 1147 1484 1157
rect 1432 1113 1440 1147
rect 1440 1113 1474 1147
rect 1474 1113 1484 1147
rect 1432 1105 1484 1113
rect 1512 1147 1564 1157
rect 1512 1113 1520 1147
rect 1520 1113 1554 1147
rect 1554 1113 1564 1147
rect 1512 1105 1564 1113
rect 2004 1147 2056 1157
rect 2004 1113 2012 1147
rect 2012 1113 2046 1147
rect 2046 1113 2056 1147
rect 2004 1105 2056 1113
rect 2084 1147 2136 1157
rect 2084 1113 2092 1147
rect 2092 1113 2126 1147
rect 2126 1113 2136 1147
rect 2084 1105 2136 1113
rect 2164 1147 2216 1157
rect 2164 1113 2172 1147
rect 2172 1113 2206 1147
rect 2206 1113 2216 1147
rect 2164 1105 2216 1113
rect 2244 1147 2296 1157
rect 2244 1113 2252 1147
rect 2252 1113 2286 1147
rect 2286 1113 2296 1147
rect 2244 1105 2296 1113
rect 2610 1147 2662 1157
rect 2610 1113 2620 1147
rect 2620 1113 2654 1147
rect 2654 1113 2662 1147
rect 2610 1105 2662 1113
rect 2690 1147 2742 1157
rect 2690 1113 2700 1147
rect 2700 1113 2734 1147
rect 2734 1113 2742 1147
rect 2690 1105 2742 1113
rect 2770 1147 2822 1157
rect 2770 1113 2780 1147
rect 2780 1113 2814 1147
rect 2814 1113 2822 1147
rect 2770 1105 2822 1113
rect 2850 1147 2902 1157
rect 2850 1113 2860 1147
rect 2860 1113 2894 1147
rect 2894 1113 2902 1147
rect 2850 1105 2902 1113
rect 3216 1147 3268 1157
rect 3216 1113 3224 1147
rect 3224 1113 3258 1147
rect 3258 1113 3268 1147
rect 3216 1105 3268 1113
rect 3296 1147 3348 1157
rect 3296 1113 3304 1147
rect 3304 1113 3338 1147
rect 3338 1113 3348 1147
rect 3296 1105 3348 1113
rect 3376 1147 3428 1157
rect 3376 1113 3384 1147
rect 3384 1113 3418 1147
rect 3418 1113 3428 1147
rect 3376 1105 3428 1113
rect 3456 1147 3508 1157
rect 3456 1113 3464 1147
rect 3464 1113 3498 1147
rect 3498 1113 3508 1147
rect 3456 1105 3508 1113
rect 3822 1147 3874 1157
rect 3822 1113 3832 1147
rect 3832 1113 3866 1147
rect 3866 1113 3874 1147
rect 3822 1105 3874 1113
rect 3902 1147 3954 1157
rect 3902 1113 3912 1147
rect 3912 1113 3946 1147
rect 3946 1113 3954 1147
rect 3902 1105 3954 1113
rect 3982 1147 4034 1157
rect 3982 1113 3992 1147
rect 3992 1113 4026 1147
rect 4026 1113 4034 1147
rect 3982 1105 4034 1113
rect 4062 1147 4114 1157
rect 4062 1113 4072 1147
rect 4072 1113 4106 1147
rect 4106 1113 4114 1147
rect 4062 1105 4114 1113
rect 4554 1147 4606 1157
rect 4554 1113 4562 1147
rect 4562 1113 4596 1147
rect 4596 1113 4606 1147
rect 4554 1105 4606 1113
rect 4634 1147 4686 1157
rect 4634 1113 4642 1147
rect 4642 1113 4676 1147
rect 4676 1113 4686 1147
rect 4634 1105 4686 1113
rect 4714 1147 4766 1157
rect 4714 1113 4722 1147
rect 4722 1113 4756 1147
rect 4756 1113 4766 1147
rect 4714 1105 4766 1113
rect 4794 1147 4846 1157
rect 4794 1113 4802 1147
rect 4802 1113 4836 1147
rect 4836 1113 4846 1147
rect 4794 1105 4846 1113
rect 5160 1147 5212 1157
rect 5160 1113 5170 1147
rect 5170 1113 5204 1147
rect 5204 1113 5212 1147
rect 5160 1105 5212 1113
rect 5240 1147 5292 1157
rect 5240 1113 5250 1147
rect 5250 1113 5284 1147
rect 5284 1113 5292 1147
rect 5240 1105 5292 1113
rect 5320 1147 5372 1157
rect 5320 1113 5330 1147
rect 5330 1113 5364 1147
rect 5364 1113 5372 1147
rect 5320 1105 5372 1113
rect 5400 1147 5452 1157
rect 5400 1113 5410 1147
rect 5410 1113 5444 1147
rect 5444 1113 5452 1147
rect 5400 1105 5452 1113
rect 7121 2186 7173 2238
rect 13185 2753 13237 2805
rect 7933 2542 7997 2545
rect 7933 2482 7955 2542
rect 7955 2482 7989 2542
rect 7989 2482 7997 2542
rect 7933 2481 7997 2482
rect 8665 2545 8729 2548
rect 8665 2485 8687 2545
rect 8687 2485 8721 2545
rect 8721 2485 8729 2545
rect 8665 2484 8729 2485
rect 8893 2545 8957 2548
rect 8893 2485 8901 2545
rect 8901 2485 8935 2545
rect 8935 2485 8957 2545
rect 8893 2484 8957 2485
rect 9877 2545 9941 2548
rect 9877 2485 9899 2545
rect 9899 2485 9933 2545
rect 9933 2485 9941 2545
rect 9877 2484 9941 2485
rect 10105 2545 10169 2548
rect 10105 2485 10113 2545
rect 10113 2485 10147 2545
rect 10147 2485 10169 2545
rect 10105 2484 10169 2485
rect 11089 2545 11153 2548
rect 11089 2485 11111 2545
rect 11111 2485 11145 2545
rect 11145 2485 11153 2545
rect 11089 2484 11153 2485
rect 11317 2545 11381 2548
rect 11317 2485 11325 2545
rect 11325 2485 11359 2545
rect 11359 2485 11381 2545
rect 11317 2484 11381 2485
rect 12301 2545 12365 2548
rect 12301 2485 12323 2545
rect 12323 2485 12357 2545
rect 12357 2485 12365 2545
rect 12301 2484 12365 2485
rect 12529 2545 12593 2548
rect 12529 2485 12537 2545
rect 12537 2485 12571 2545
rect 12571 2485 12593 2545
rect 12529 2484 12593 2485
rect 13273 2492 13282 2544
rect 13282 2492 13316 2544
rect 13316 2492 13325 2544
rect 8289 2344 8353 2346
rect 8289 2284 8308 2344
rect 8308 2284 8342 2344
rect 8342 2284 8353 2344
rect 8289 2282 8353 2284
rect 9021 2344 9085 2346
rect 9021 2284 9040 2344
rect 9040 2284 9074 2344
rect 9074 2284 9085 2344
rect 9021 2282 9085 2284
rect 9239 2344 9303 2346
rect 9239 2284 9250 2344
rect 9250 2284 9284 2344
rect 9284 2284 9303 2344
rect 9239 2282 9303 2284
rect 10233 2344 10297 2346
rect 10233 2284 10252 2344
rect 10252 2284 10286 2344
rect 10286 2284 10297 2344
rect 10233 2282 10297 2284
rect 10451 2344 10515 2346
rect 10451 2284 10462 2344
rect 10462 2284 10496 2344
rect 10496 2284 10515 2344
rect 10451 2282 10515 2284
rect 11571 2344 11635 2346
rect 11571 2284 11590 2344
rect 11590 2284 11624 2344
rect 11624 2284 11635 2344
rect 11571 2282 11635 2284
rect 11789 2344 11853 2346
rect 11789 2284 11800 2344
rect 11800 2284 11834 2344
rect 11834 2284 11853 2344
rect 11789 2282 11853 2284
rect 12523 2344 12587 2346
rect 12523 2284 12534 2344
rect 12534 2284 12568 2344
rect 12568 2284 12587 2344
rect 12523 2282 12587 2284
rect 13273 2289 13282 2341
rect 13282 2289 13316 2341
rect 13316 2289 13325 2341
rect 7609 2186 7661 2238
rect 6473 2027 6525 2079
rect 5894 1147 5946 1157
rect 5894 1113 5904 1147
rect 5904 1113 5938 1147
rect 5938 1113 5946 1147
rect 5894 1105 5946 1113
rect 5974 1147 6026 1157
rect 5974 1113 5984 1147
rect 5984 1113 6018 1147
rect 6018 1113 6026 1147
rect 5974 1105 6026 1113
rect 6054 1147 6106 1157
rect 6054 1113 6064 1147
rect 6064 1113 6098 1147
rect 6098 1113 6106 1147
rect 6054 1105 6106 1113
rect 6134 1147 6186 1157
rect 6134 1113 6144 1147
rect 6144 1113 6178 1147
rect 6178 1113 6186 1147
rect 6134 1105 6186 1113
rect 7439 1134 7448 1154
rect 7448 1134 7482 1154
rect 7482 1134 7491 1154
rect 7439 1102 7491 1134
rect 7981 1147 8033 1157
rect 7981 1113 7989 1147
rect 7989 1113 8023 1147
rect 8023 1113 8033 1147
rect 7981 1105 8033 1113
rect 8061 1147 8113 1157
rect 8061 1113 8069 1147
rect 8069 1113 8103 1147
rect 8103 1113 8113 1147
rect 8061 1105 8113 1113
rect 8141 1147 8193 1157
rect 8141 1113 8149 1147
rect 8149 1113 8183 1147
rect 8183 1113 8193 1147
rect 8141 1105 8193 1113
rect 8221 1147 8273 1157
rect 8221 1113 8229 1147
rect 8229 1113 8263 1147
rect 8263 1113 8273 1147
rect 8221 1105 8273 1113
rect 8713 1147 8765 1157
rect 8713 1113 8721 1147
rect 8721 1113 8755 1147
rect 8755 1113 8765 1147
rect 8713 1105 8765 1113
rect 8793 1147 8845 1157
rect 8793 1113 8801 1147
rect 8801 1113 8835 1147
rect 8835 1113 8845 1147
rect 8793 1105 8845 1113
rect 8873 1147 8925 1157
rect 8873 1113 8881 1147
rect 8881 1113 8915 1147
rect 8915 1113 8925 1147
rect 8873 1105 8925 1113
rect 8953 1147 9005 1157
rect 8953 1113 8961 1147
rect 8961 1113 8995 1147
rect 8995 1113 9005 1147
rect 8953 1105 9005 1113
rect 9319 1147 9371 1157
rect 9319 1113 9329 1147
rect 9329 1113 9363 1147
rect 9363 1113 9371 1147
rect 9319 1105 9371 1113
rect 9399 1147 9451 1157
rect 9399 1113 9409 1147
rect 9409 1113 9443 1147
rect 9443 1113 9451 1147
rect 9399 1105 9451 1113
rect 9479 1147 9531 1157
rect 9479 1113 9489 1147
rect 9489 1113 9523 1147
rect 9523 1113 9531 1147
rect 9479 1105 9531 1113
rect 9559 1147 9611 1157
rect 9559 1113 9569 1147
rect 9569 1113 9603 1147
rect 9603 1113 9611 1147
rect 9559 1105 9611 1113
rect 9925 1147 9977 1157
rect 9925 1113 9933 1147
rect 9933 1113 9967 1147
rect 9967 1113 9977 1147
rect 9925 1105 9977 1113
rect 10005 1147 10057 1157
rect 10005 1113 10013 1147
rect 10013 1113 10047 1147
rect 10047 1113 10057 1147
rect 10005 1105 10057 1113
rect 10085 1147 10137 1157
rect 10085 1113 10093 1147
rect 10093 1113 10127 1147
rect 10127 1113 10137 1147
rect 10085 1105 10137 1113
rect 10165 1147 10217 1157
rect 10165 1113 10173 1147
rect 10173 1113 10207 1147
rect 10207 1113 10217 1147
rect 10165 1105 10217 1113
rect 10531 1147 10583 1157
rect 10531 1113 10541 1147
rect 10541 1113 10575 1147
rect 10575 1113 10583 1147
rect 10531 1105 10583 1113
rect 10611 1147 10663 1157
rect 10611 1113 10621 1147
rect 10621 1113 10655 1147
rect 10655 1113 10663 1147
rect 10611 1105 10663 1113
rect 10691 1147 10743 1157
rect 10691 1113 10701 1147
rect 10701 1113 10735 1147
rect 10735 1113 10743 1147
rect 10691 1105 10743 1113
rect 10771 1147 10823 1157
rect 10771 1113 10781 1147
rect 10781 1113 10815 1147
rect 10815 1113 10823 1147
rect 10771 1105 10823 1113
rect 11263 1147 11315 1157
rect 11263 1113 11271 1147
rect 11271 1113 11305 1147
rect 11305 1113 11315 1147
rect 11263 1105 11315 1113
rect 11343 1147 11395 1157
rect 11343 1113 11351 1147
rect 11351 1113 11385 1147
rect 11385 1113 11395 1147
rect 11343 1105 11395 1113
rect 11423 1147 11475 1157
rect 11423 1113 11431 1147
rect 11431 1113 11465 1147
rect 11465 1113 11475 1147
rect 11423 1105 11475 1113
rect 11503 1147 11555 1157
rect 11503 1113 11511 1147
rect 11511 1113 11545 1147
rect 11545 1113 11555 1147
rect 11503 1105 11555 1113
rect 11869 1147 11921 1157
rect 11869 1113 11879 1147
rect 11879 1113 11913 1147
rect 11913 1113 11921 1147
rect 11869 1105 11921 1113
rect 11949 1147 12001 1157
rect 11949 1113 11959 1147
rect 11959 1113 11993 1147
rect 11993 1113 12001 1147
rect 11949 1105 12001 1113
rect 12029 1147 12081 1157
rect 12029 1113 12039 1147
rect 12039 1113 12073 1147
rect 12073 1113 12081 1147
rect 12029 1105 12081 1113
rect 12109 1147 12161 1157
rect 12109 1113 12119 1147
rect 12119 1113 12153 1147
rect 12153 1113 12161 1147
rect 12109 1105 12161 1113
rect 13182 2027 13234 2079
rect 12603 1147 12655 1157
rect 12603 1113 12613 1147
rect 12613 1113 12647 1147
rect 12647 1113 12655 1147
rect 12603 1105 12655 1113
rect 12683 1147 12735 1157
rect 12683 1113 12693 1147
rect 12693 1113 12727 1147
rect 12727 1113 12735 1147
rect 12683 1105 12735 1113
rect 12763 1147 12815 1157
rect 12763 1113 12773 1147
rect 12773 1113 12807 1147
rect 12807 1113 12815 1147
rect 12763 1105 12815 1113
rect 12843 1147 12895 1157
rect 12843 1113 12853 1147
rect 12853 1113 12887 1147
rect 12887 1113 12895 1147
rect 12843 1105 12895 1113
rect 900 632 952 684
rect 5800 622 5853 674
rect 7609 624 7661 677
rect 12504 621 12568 685
rect 569 208 621 216
rect 569 174 577 208
rect 577 174 611 208
rect 611 174 621 208
rect 569 164 621 174
rect 649 208 701 216
rect 649 174 657 208
rect 657 174 691 208
rect 691 174 701 208
rect 649 164 701 174
rect 729 208 781 216
rect 729 174 737 208
rect 737 174 771 208
rect 771 174 781 208
rect 729 164 781 174
rect 809 208 861 216
rect 809 174 817 208
rect 817 174 851 208
rect 851 174 861 208
rect 809 164 861 174
rect 230 -758 282 -706
rect 1303 208 1355 216
rect 1303 174 1311 208
rect 1311 174 1345 208
rect 1345 174 1355 208
rect 1303 164 1355 174
rect 1383 208 1435 216
rect 1383 174 1391 208
rect 1391 174 1425 208
rect 1425 174 1435 208
rect 1383 164 1435 174
rect 1463 208 1515 216
rect 1463 174 1471 208
rect 1471 174 1505 208
rect 1505 174 1515 208
rect 1463 164 1515 174
rect 1543 208 1595 216
rect 1543 174 1551 208
rect 1551 174 1585 208
rect 1585 174 1595 208
rect 1543 164 1595 174
rect 1909 208 1961 216
rect 1909 174 1919 208
rect 1919 174 1953 208
rect 1953 174 1961 208
rect 1909 164 1961 174
rect 1989 208 2041 216
rect 1989 174 1999 208
rect 1999 174 2033 208
rect 2033 174 2041 208
rect 1989 164 2041 174
rect 2069 208 2121 216
rect 2069 174 2079 208
rect 2079 174 2113 208
rect 2113 174 2121 208
rect 2069 164 2121 174
rect 2149 208 2201 216
rect 2149 174 2159 208
rect 2159 174 2193 208
rect 2193 174 2201 208
rect 2149 164 2201 174
rect 2641 208 2693 216
rect 2641 174 2649 208
rect 2649 174 2683 208
rect 2683 174 2693 208
rect 2641 164 2693 174
rect 2721 208 2773 216
rect 2721 174 2729 208
rect 2729 174 2763 208
rect 2763 174 2773 208
rect 2721 164 2773 174
rect 2801 208 2853 216
rect 2801 174 2809 208
rect 2809 174 2843 208
rect 2843 174 2853 208
rect 2801 164 2853 174
rect 2881 208 2933 216
rect 2881 174 2889 208
rect 2889 174 2923 208
rect 2923 174 2933 208
rect 2881 164 2933 174
rect 3247 208 3299 216
rect 3247 174 3257 208
rect 3257 174 3291 208
rect 3291 174 3299 208
rect 3247 164 3299 174
rect 3327 208 3379 216
rect 3327 174 3337 208
rect 3337 174 3371 208
rect 3371 174 3379 208
rect 3327 164 3379 174
rect 3407 208 3459 216
rect 3407 174 3417 208
rect 3417 174 3451 208
rect 3451 174 3459 208
rect 3407 164 3459 174
rect 3487 208 3539 216
rect 3487 174 3497 208
rect 3497 174 3531 208
rect 3531 174 3539 208
rect 3487 164 3539 174
rect 3853 208 3905 216
rect 3853 174 3861 208
rect 3861 174 3895 208
rect 3895 174 3905 208
rect 3853 164 3905 174
rect 3933 208 3985 216
rect 3933 174 3941 208
rect 3941 174 3975 208
rect 3975 174 3985 208
rect 3933 164 3985 174
rect 4013 208 4065 216
rect 4013 174 4021 208
rect 4021 174 4055 208
rect 4055 174 4065 208
rect 4013 164 4065 174
rect 4093 208 4145 216
rect 4093 174 4101 208
rect 4101 174 4135 208
rect 4135 174 4145 208
rect 4093 164 4145 174
rect 4459 208 4511 216
rect 4459 174 4469 208
rect 4469 174 4503 208
rect 4503 174 4511 208
rect 4459 164 4511 174
rect 4539 208 4591 216
rect 4539 174 4549 208
rect 4549 174 4583 208
rect 4583 174 4591 208
rect 4539 164 4591 174
rect 4619 208 4671 216
rect 4619 174 4629 208
rect 4629 174 4663 208
rect 4663 174 4671 208
rect 4619 164 4671 174
rect 4699 208 4751 216
rect 4699 174 4709 208
rect 4709 174 4743 208
rect 4743 174 4751 208
rect 4699 164 4751 174
rect 5191 208 5243 216
rect 5191 174 5201 208
rect 5201 174 5235 208
rect 5235 174 5243 208
rect 5191 164 5243 174
rect 5271 208 5323 216
rect 5271 174 5281 208
rect 5281 174 5315 208
rect 5315 174 5323 208
rect 5271 164 5323 174
rect 5351 208 5403 216
rect 5351 174 5361 208
rect 5361 174 5395 208
rect 5395 174 5403 208
rect 5351 164 5403 174
rect 5431 208 5483 216
rect 5431 174 5441 208
rect 5441 174 5475 208
rect 5475 174 5483 208
rect 5431 164 5483 174
rect 5973 187 6025 219
rect 5973 167 5982 187
rect 5982 167 6016 187
rect 6016 167 6025 187
rect 7278 208 7330 216
rect 7278 174 7286 208
rect 7286 174 7320 208
rect 7320 174 7330 208
rect 7278 164 7330 174
rect 7358 208 7410 216
rect 7358 174 7366 208
rect 7366 174 7400 208
rect 7400 174 7410 208
rect 7358 164 7410 174
rect 7438 208 7490 216
rect 7438 174 7446 208
rect 7446 174 7480 208
rect 7480 174 7490 208
rect 7438 164 7490 174
rect 7518 208 7570 216
rect 7518 174 7526 208
rect 7526 174 7560 208
rect 7560 174 7570 208
rect 7518 164 7570 174
rect 6939 -758 6991 -706
rect 5803 -917 5855 -865
rect 139 -1020 148 -968
rect 148 -1020 182 -968
rect 182 -1020 191 -968
rect 877 -963 941 -961
rect 877 -1023 896 -963
rect 896 -1023 930 -963
rect 930 -1023 941 -963
rect 877 -1025 941 -1023
rect 1611 -963 1675 -961
rect 1611 -1023 1630 -963
rect 1630 -1023 1664 -963
rect 1664 -1023 1675 -963
rect 1611 -1025 1675 -1023
rect 1829 -963 1893 -961
rect 1829 -1023 1840 -963
rect 1840 -1023 1874 -963
rect 1874 -1023 1893 -963
rect 1829 -1025 1893 -1023
rect 2949 -963 3013 -961
rect 2949 -1023 2968 -963
rect 2968 -1023 3002 -963
rect 3002 -1023 3013 -963
rect 2949 -1025 3013 -1023
rect 3167 -963 3231 -961
rect 3167 -1023 3178 -963
rect 3178 -1023 3212 -963
rect 3212 -1023 3231 -963
rect 3167 -1025 3231 -1023
rect 4161 -963 4225 -961
rect 4161 -1023 4180 -963
rect 4180 -1023 4214 -963
rect 4214 -1023 4225 -963
rect 4161 -1025 4225 -1023
rect 4379 -963 4443 -961
rect 4379 -1023 4390 -963
rect 4390 -1023 4424 -963
rect 4424 -1023 4443 -963
rect 4379 -1025 4443 -1023
rect 5111 -963 5175 -961
rect 5111 -1023 5122 -963
rect 5122 -1023 5156 -963
rect 5156 -1023 5175 -963
rect 5111 -1025 5175 -1023
rect 139 -1223 148 -1171
rect 148 -1223 182 -1171
rect 182 -1223 191 -1171
rect 871 -1164 935 -1163
rect 871 -1224 893 -1164
rect 893 -1224 927 -1164
rect 927 -1224 935 -1164
rect 871 -1227 935 -1224
rect 1099 -1164 1163 -1163
rect 1099 -1224 1107 -1164
rect 1107 -1224 1141 -1164
rect 1141 -1224 1163 -1164
rect 1099 -1227 1163 -1224
rect 2083 -1164 2147 -1163
rect 2083 -1224 2105 -1164
rect 2105 -1224 2139 -1164
rect 2139 -1224 2147 -1164
rect 2083 -1227 2147 -1224
rect 2311 -1164 2375 -1163
rect 2311 -1224 2319 -1164
rect 2319 -1224 2353 -1164
rect 2353 -1224 2375 -1164
rect 2311 -1227 2375 -1224
rect 3295 -1164 3359 -1163
rect 3295 -1224 3317 -1164
rect 3317 -1224 3351 -1164
rect 3351 -1224 3359 -1164
rect 3295 -1227 3359 -1224
rect 3523 -1164 3587 -1163
rect 3523 -1224 3531 -1164
rect 3531 -1224 3565 -1164
rect 3565 -1224 3587 -1164
rect 3523 -1227 3587 -1224
rect 4507 -1164 4571 -1163
rect 4507 -1224 4529 -1164
rect 4529 -1224 4563 -1164
rect 4563 -1224 4571 -1164
rect 4507 -1227 4571 -1224
rect 4735 -1164 4799 -1163
rect 4735 -1224 4743 -1164
rect 4743 -1224 4777 -1164
rect 4777 -1224 4799 -1164
rect 4735 -1227 4799 -1224
rect 5467 -1161 5531 -1160
rect 5467 -1221 5475 -1161
rect 5475 -1221 5509 -1161
rect 5509 -1221 5531 -1161
rect 5467 -1224 5531 -1221
rect 227 -1484 279 -1432
rect 6291 -917 6343 -865
rect 8012 208 8064 216
rect 8012 174 8020 208
rect 8020 174 8054 208
rect 8054 174 8064 208
rect 8012 164 8064 174
rect 8092 208 8144 216
rect 8092 174 8100 208
rect 8100 174 8134 208
rect 8134 174 8144 208
rect 8092 164 8144 174
rect 8172 208 8224 216
rect 8172 174 8180 208
rect 8180 174 8214 208
rect 8214 174 8224 208
rect 8172 164 8224 174
rect 8252 208 8304 216
rect 8252 174 8260 208
rect 8260 174 8294 208
rect 8294 174 8304 208
rect 8252 164 8304 174
rect 8618 208 8670 216
rect 8618 174 8628 208
rect 8628 174 8662 208
rect 8662 174 8670 208
rect 8618 164 8670 174
rect 8698 208 8750 216
rect 8698 174 8708 208
rect 8708 174 8742 208
rect 8742 174 8750 208
rect 8698 164 8750 174
rect 8778 208 8830 216
rect 8778 174 8788 208
rect 8788 174 8822 208
rect 8822 174 8830 208
rect 8778 164 8830 174
rect 8858 208 8910 216
rect 8858 174 8868 208
rect 8868 174 8902 208
rect 8902 174 8910 208
rect 8858 164 8910 174
rect 9350 208 9402 216
rect 9350 174 9358 208
rect 9358 174 9392 208
rect 9392 174 9402 208
rect 9350 164 9402 174
rect 9430 208 9482 216
rect 9430 174 9438 208
rect 9438 174 9472 208
rect 9472 174 9482 208
rect 9430 164 9482 174
rect 9510 208 9562 216
rect 9510 174 9518 208
rect 9518 174 9552 208
rect 9552 174 9562 208
rect 9510 164 9562 174
rect 9590 208 9642 216
rect 9590 174 9598 208
rect 9598 174 9632 208
rect 9632 174 9642 208
rect 9590 164 9642 174
rect 9956 208 10008 216
rect 9956 174 9966 208
rect 9966 174 10000 208
rect 10000 174 10008 208
rect 9956 164 10008 174
rect 10036 208 10088 216
rect 10036 174 10046 208
rect 10046 174 10080 208
rect 10080 174 10088 208
rect 10036 164 10088 174
rect 10116 208 10168 216
rect 10116 174 10126 208
rect 10126 174 10160 208
rect 10160 174 10168 208
rect 10116 164 10168 174
rect 10196 208 10248 216
rect 10196 174 10206 208
rect 10206 174 10240 208
rect 10240 174 10248 208
rect 10196 164 10248 174
rect 10562 208 10614 216
rect 10562 174 10570 208
rect 10570 174 10604 208
rect 10604 174 10614 208
rect 10562 164 10614 174
rect 10642 208 10694 216
rect 10642 174 10650 208
rect 10650 174 10684 208
rect 10684 174 10694 208
rect 10642 164 10694 174
rect 10722 208 10774 216
rect 10722 174 10730 208
rect 10730 174 10764 208
rect 10764 174 10774 208
rect 10722 164 10774 174
rect 10802 208 10854 216
rect 10802 174 10810 208
rect 10810 174 10844 208
rect 10844 174 10854 208
rect 10802 164 10854 174
rect 11168 208 11220 216
rect 11168 174 11178 208
rect 11178 174 11212 208
rect 11212 174 11220 208
rect 11168 164 11220 174
rect 11248 208 11300 216
rect 11248 174 11258 208
rect 11258 174 11292 208
rect 11292 174 11300 208
rect 11248 164 11300 174
rect 11328 208 11380 216
rect 11328 174 11338 208
rect 11338 174 11372 208
rect 11372 174 11380 208
rect 11328 164 11380 174
rect 11408 208 11460 216
rect 11408 174 11418 208
rect 11418 174 11452 208
rect 11452 174 11460 208
rect 11408 164 11460 174
rect 11900 208 11952 216
rect 11900 174 11910 208
rect 11910 174 11944 208
rect 11944 174 11952 208
rect 11900 164 11952 174
rect 11980 208 12032 216
rect 11980 174 11990 208
rect 11990 174 12024 208
rect 12024 174 12032 208
rect 11980 164 12032 174
rect 12060 208 12112 216
rect 12060 174 12070 208
rect 12070 174 12104 208
rect 12104 174 12112 208
rect 12060 164 12112 174
rect 12140 208 12192 216
rect 12140 174 12150 208
rect 12150 174 12184 208
rect 12184 174 12192 208
rect 12140 164 12192 174
rect 12682 187 12734 219
rect 12682 167 12691 187
rect 12691 167 12725 187
rect 12725 167 12734 187
rect 12512 -917 12564 -865
rect 6848 -1020 6857 -968
rect 6857 -1020 6891 -968
rect 6891 -1020 6900 -968
rect 7586 -963 7650 -961
rect 7586 -1023 7605 -963
rect 7605 -1023 7639 -963
rect 7639 -1023 7650 -963
rect 7586 -1025 7650 -1023
rect 8320 -963 8384 -961
rect 8320 -1023 8339 -963
rect 8339 -1023 8373 -963
rect 8373 -1023 8384 -963
rect 8320 -1025 8384 -1023
rect 8538 -963 8602 -961
rect 8538 -1023 8549 -963
rect 8549 -1023 8583 -963
rect 8583 -1023 8602 -963
rect 8538 -1025 8602 -1023
rect 9658 -963 9722 -961
rect 9658 -1023 9677 -963
rect 9677 -1023 9711 -963
rect 9711 -1023 9722 -963
rect 9658 -1025 9722 -1023
rect 9876 -963 9940 -961
rect 9876 -1023 9887 -963
rect 9887 -1023 9921 -963
rect 9921 -1023 9940 -963
rect 9876 -1025 9940 -1023
rect 10870 -963 10934 -961
rect 10870 -1023 10889 -963
rect 10889 -1023 10923 -963
rect 10923 -1023 10934 -963
rect 10870 -1025 10934 -1023
rect 11088 -963 11152 -961
rect 11088 -1023 11099 -963
rect 11099 -1023 11133 -963
rect 11133 -1023 11152 -963
rect 11088 -1025 11152 -1023
rect 11820 -963 11884 -961
rect 11820 -1023 11831 -963
rect 11831 -1023 11865 -963
rect 11865 -1023 11884 -963
rect 11820 -1025 11884 -1023
rect 6295 -1217 6347 -1208
rect 6438 -1217 6490 -1208
rect 6558 -1217 6610 -1208
rect 6295 -1251 6296 -1217
rect 6296 -1251 6347 -1217
rect 6438 -1251 6446 -1217
rect 6446 -1251 6480 -1217
rect 6480 -1251 6490 -1217
rect 6558 -1251 6572 -1217
rect 6572 -1251 6610 -1217
rect 6295 -1260 6347 -1251
rect 6438 -1260 6490 -1251
rect 6558 -1260 6610 -1251
rect 6848 -1223 6857 -1171
rect 6857 -1223 6891 -1171
rect 6891 -1223 6900 -1171
rect 7580 -1164 7644 -1163
rect 7580 -1224 7602 -1164
rect 7602 -1224 7636 -1164
rect 7636 -1224 7644 -1164
rect 7580 -1227 7644 -1224
rect 7808 -1164 7872 -1163
rect 7808 -1224 7816 -1164
rect 7816 -1224 7850 -1164
rect 7850 -1224 7872 -1164
rect 7808 -1227 7872 -1224
rect 8792 -1164 8856 -1163
rect 8792 -1224 8814 -1164
rect 8814 -1224 8848 -1164
rect 8848 -1224 8856 -1164
rect 8792 -1227 8856 -1224
rect 9020 -1164 9084 -1163
rect 9020 -1224 9028 -1164
rect 9028 -1224 9062 -1164
rect 9062 -1224 9084 -1164
rect 9020 -1227 9084 -1224
rect 10004 -1164 10068 -1163
rect 10004 -1224 10026 -1164
rect 10026 -1224 10060 -1164
rect 10060 -1224 10068 -1164
rect 10004 -1227 10068 -1224
rect 10232 -1164 10296 -1163
rect 10232 -1224 10240 -1164
rect 10240 -1224 10274 -1164
rect 10274 -1224 10296 -1164
rect 10232 -1227 10296 -1224
rect 11216 -1164 11280 -1163
rect 11216 -1224 11238 -1164
rect 11238 -1224 11272 -1164
rect 11272 -1224 11280 -1164
rect 11216 -1227 11280 -1224
rect 11444 -1164 11508 -1163
rect 11444 -1224 11452 -1164
rect 11452 -1224 11486 -1164
rect 11486 -1224 11508 -1164
rect 11444 -1227 11508 -1224
rect 12176 -1161 12240 -1160
rect 12176 -1221 12184 -1161
rect 12184 -1221 12218 -1161
rect 12218 -1221 12240 -1161
rect 12176 -1224 12240 -1221
rect 145 -1685 197 -1674
rect 145 -1719 152 -1685
rect 152 -1719 186 -1685
rect 186 -1719 197 -1685
rect 145 -1726 197 -1719
rect 6303 -1452 6355 -1443
rect 6303 -1486 6309 -1452
rect 6309 -1486 6343 -1452
rect 6343 -1486 6355 -1452
rect 6303 -1495 6355 -1486
rect 6936 -1484 6988 -1432
rect 13000 -917 13052 -865
rect 13004 -1217 13056 -1208
rect 13147 -1217 13199 -1208
rect 13267 -1217 13319 -1208
rect 13004 -1251 13005 -1217
rect 13005 -1251 13056 -1217
rect 13147 -1251 13155 -1217
rect 13155 -1251 13189 -1217
rect 13189 -1251 13199 -1217
rect 13267 -1251 13281 -1217
rect 13281 -1251 13319 -1217
rect 13004 -1260 13056 -1251
rect 13147 -1260 13199 -1251
rect 13267 -1260 13319 -1251
rect 144 -1842 196 -1831
rect 144 -1876 151 -1842
rect 151 -1876 185 -1842
rect 185 -1876 196 -1842
rect 144 -1883 196 -1876
rect 6854 -1685 6906 -1674
rect 6854 -1719 6861 -1685
rect 6861 -1719 6895 -1685
rect 6895 -1719 6906 -1685
rect 6854 -1726 6906 -1719
rect 13012 -1452 13064 -1443
rect 13012 -1486 13018 -1452
rect 13018 -1486 13052 -1452
rect 13052 -1486 13064 -1452
rect 13012 -1495 13064 -1486
rect 6301 -1806 6353 -1754
rect 6445 -1761 6497 -1753
rect 6445 -1795 6446 -1761
rect 6446 -1795 6480 -1761
rect 6480 -1795 6497 -1761
rect 6445 -1805 6497 -1795
rect 6576 -1806 6628 -1754
rect 6853 -1842 6905 -1831
rect 6853 -1876 6860 -1842
rect 6860 -1876 6894 -1842
rect 6894 -1876 6905 -1842
rect 6853 -1883 6905 -1876
rect 144 -2012 196 -2001
rect 144 -2046 151 -2012
rect 151 -2046 185 -2012
rect 185 -2046 196 -2012
rect 144 -2053 196 -2046
rect 145 -2164 197 -2153
rect 145 -2198 152 -2164
rect 152 -2198 186 -2164
rect 186 -2198 197 -2164
rect 145 -2205 197 -2198
rect 13010 -1806 13062 -1754
rect 13154 -1761 13206 -1753
rect 13154 -1795 13155 -1761
rect 13155 -1795 13189 -1761
rect 13189 -1795 13206 -1761
rect 13154 -1805 13206 -1795
rect 13285 -1806 13337 -1754
rect 6431 -1914 6483 -1903
rect 6431 -1948 6438 -1914
rect 6438 -1948 6472 -1914
rect 6472 -1948 6483 -1914
rect 6431 -1955 6483 -1948
rect 6853 -2012 6905 -2001
rect 6853 -2046 6860 -2012
rect 6860 -2046 6894 -2012
rect 6894 -2046 6905 -2012
rect 6853 -2053 6905 -2046
rect 6431 -2110 6483 -2099
rect 6431 -2144 6438 -2110
rect 6438 -2144 6472 -2110
rect 6472 -2144 6483 -2110
rect 6431 -2151 6483 -2144
rect 6854 -2164 6906 -2153
rect 6854 -2198 6861 -2164
rect 6861 -2198 6895 -2164
rect 6895 -2198 6906 -2164
rect 6854 -2205 6906 -2198
rect 150 -2308 202 -2297
rect 150 -2342 157 -2308
rect 157 -2342 191 -2308
rect 191 -2342 202 -2308
rect 150 -2349 202 -2342
rect 489 -2359 541 -2353
rect 489 -2393 499 -2359
rect 499 -2393 533 -2359
rect 533 -2393 541 -2359
rect 489 -2405 541 -2393
rect 569 -2359 621 -2353
rect 569 -2393 579 -2359
rect 579 -2393 613 -2359
rect 613 -2393 621 -2359
rect 569 -2405 621 -2393
rect 649 -2359 701 -2353
rect 649 -2393 659 -2359
rect 659 -2393 693 -2359
rect 693 -2393 701 -2359
rect 649 -2405 701 -2393
rect 729 -2359 781 -2353
rect 729 -2393 739 -2359
rect 739 -2393 773 -2359
rect 773 -2393 781 -2359
rect 729 -2405 781 -2393
rect 809 -2359 861 -2353
rect 809 -2393 819 -2359
rect 819 -2393 853 -2359
rect 853 -2393 861 -2359
rect 809 -2405 861 -2393
rect 889 -2359 941 -2353
rect 889 -2393 899 -2359
rect 899 -2393 933 -2359
rect 933 -2393 941 -2359
rect 889 -2405 941 -2393
rect 1093 -2359 1145 -2353
rect 1093 -2393 1101 -2359
rect 1101 -2393 1135 -2359
rect 1135 -2393 1145 -2359
rect 1093 -2405 1145 -2393
rect 1173 -2359 1225 -2353
rect 1173 -2393 1181 -2359
rect 1181 -2393 1215 -2359
rect 1215 -2393 1225 -2359
rect 1173 -2405 1225 -2393
rect 1253 -2359 1305 -2353
rect 1253 -2393 1261 -2359
rect 1261 -2393 1295 -2359
rect 1295 -2393 1305 -2359
rect 1253 -2405 1305 -2393
rect 1333 -2359 1385 -2353
rect 1333 -2393 1341 -2359
rect 1341 -2393 1375 -2359
rect 1375 -2393 1385 -2359
rect 1333 -2405 1385 -2393
rect 1413 -2359 1465 -2353
rect 1413 -2393 1421 -2359
rect 1421 -2393 1455 -2359
rect 1455 -2393 1465 -2359
rect 1413 -2405 1465 -2393
rect 1493 -2359 1545 -2353
rect 1493 -2393 1501 -2359
rect 1501 -2393 1535 -2359
rect 1535 -2393 1545 -2359
rect 1493 -2405 1545 -2393
rect 1701 -2359 1753 -2353
rect 1701 -2393 1711 -2359
rect 1711 -2393 1745 -2359
rect 1745 -2393 1753 -2359
rect 1701 -2405 1753 -2393
rect 1781 -2359 1833 -2353
rect 1781 -2393 1791 -2359
rect 1791 -2393 1825 -2359
rect 1825 -2393 1833 -2359
rect 1781 -2405 1833 -2393
rect 1861 -2359 1913 -2353
rect 1861 -2393 1871 -2359
rect 1871 -2393 1905 -2359
rect 1905 -2393 1913 -2359
rect 1861 -2405 1913 -2393
rect 1941 -2359 1993 -2353
rect 1941 -2393 1951 -2359
rect 1951 -2393 1985 -2359
rect 1985 -2393 1993 -2359
rect 1941 -2405 1993 -2393
rect 2021 -2359 2073 -2353
rect 2021 -2393 2031 -2359
rect 2031 -2393 2065 -2359
rect 2065 -2393 2073 -2359
rect 2021 -2405 2073 -2393
rect 2101 -2359 2153 -2353
rect 2101 -2393 2111 -2359
rect 2111 -2393 2145 -2359
rect 2145 -2393 2153 -2359
rect 2101 -2405 2153 -2393
rect 2305 -2359 2357 -2353
rect 2305 -2393 2313 -2359
rect 2313 -2393 2347 -2359
rect 2347 -2393 2357 -2359
rect 2305 -2405 2357 -2393
rect 2385 -2359 2437 -2353
rect 2385 -2393 2393 -2359
rect 2393 -2393 2427 -2359
rect 2427 -2393 2437 -2359
rect 2385 -2405 2437 -2393
rect 2465 -2359 2517 -2353
rect 2465 -2393 2473 -2359
rect 2473 -2393 2507 -2359
rect 2507 -2393 2517 -2359
rect 2465 -2405 2517 -2393
rect 2545 -2359 2597 -2353
rect 2545 -2393 2553 -2359
rect 2553 -2393 2587 -2359
rect 2587 -2393 2597 -2359
rect 2545 -2405 2597 -2393
rect 2625 -2359 2677 -2353
rect 2625 -2393 2633 -2359
rect 2633 -2393 2667 -2359
rect 2667 -2393 2677 -2359
rect 2625 -2405 2677 -2393
rect 2705 -2359 2757 -2353
rect 2705 -2393 2713 -2359
rect 2713 -2393 2747 -2359
rect 2747 -2393 2757 -2359
rect 2705 -2405 2757 -2393
rect 2913 -2359 2965 -2353
rect 2913 -2393 2923 -2359
rect 2923 -2393 2957 -2359
rect 2957 -2393 2965 -2359
rect 2913 -2405 2965 -2393
rect 2993 -2359 3045 -2353
rect 2993 -2393 3003 -2359
rect 3003 -2393 3037 -2359
rect 3037 -2393 3045 -2359
rect 2993 -2405 3045 -2393
rect 3073 -2359 3125 -2353
rect 3073 -2393 3083 -2359
rect 3083 -2393 3117 -2359
rect 3117 -2393 3125 -2359
rect 3073 -2405 3125 -2393
rect 3153 -2359 3205 -2353
rect 3153 -2393 3163 -2359
rect 3163 -2393 3197 -2359
rect 3197 -2393 3205 -2359
rect 3153 -2405 3205 -2393
rect 3233 -2359 3285 -2353
rect 3233 -2393 3243 -2359
rect 3243 -2393 3277 -2359
rect 3277 -2393 3285 -2359
rect 3233 -2405 3285 -2393
rect 3313 -2359 3365 -2353
rect 3313 -2393 3323 -2359
rect 3323 -2393 3357 -2359
rect 3357 -2393 3365 -2359
rect 3313 -2405 3365 -2393
rect 3517 -2359 3569 -2353
rect 3517 -2393 3525 -2359
rect 3525 -2393 3559 -2359
rect 3559 -2393 3569 -2359
rect 3517 -2405 3569 -2393
rect 3597 -2359 3649 -2353
rect 3597 -2393 3605 -2359
rect 3605 -2393 3639 -2359
rect 3639 -2393 3649 -2359
rect 3597 -2405 3649 -2393
rect 3677 -2359 3729 -2353
rect 3677 -2393 3685 -2359
rect 3685 -2393 3719 -2359
rect 3719 -2393 3729 -2359
rect 3677 -2405 3729 -2393
rect 3757 -2359 3809 -2353
rect 3757 -2393 3765 -2359
rect 3765 -2393 3799 -2359
rect 3799 -2393 3809 -2359
rect 3757 -2405 3809 -2393
rect 3837 -2359 3889 -2353
rect 3837 -2393 3845 -2359
rect 3845 -2393 3879 -2359
rect 3879 -2393 3889 -2359
rect 3837 -2405 3889 -2393
rect 3917 -2359 3969 -2353
rect 3917 -2393 3925 -2359
rect 3925 -2393 3959 -2359
rect 3959 -2393 3969 -2359
rect 3917 -2405 3969 -2393
rect 4125 -2359 4177 -2353
rect 4125 -2393 4135 -2359
rect 4135 -2393 4169 -2359
rect 4169 -2393 4177 -2359
rect 4125 -2405 4177 -2393
rect 4205 -2359 4257 -2353
rect 4205 -2393 4215 -2359
rect 4215 -2393 4249 -2359
rect 4249 -2393 4257 -2359
rect 4205 -2405 4257 -2393
rect 4285 -2359 4337 -2353
rect 4285 -2393 4295 -2359
rect 4295 -2393 4329 -2359
rect 4329 -2393 4337 -2359
rect 4285 -2405 4337 -2393
rect 4365 -2359 4417 -2353
rect 4365 -2393 4375 -2359
rect 4375 -2393 4409 -2359
rect 4409 -2393 4417 -2359
rect 4365 -2405 4417 -2393
rect 4445 -2359 4497 -2353
rect 4445 -2393 4455 -2359
rect 4455 -2393 4489 -2359
rect 4489 -2393 4497 -2359
rect 4445 -2405 4497 -2393
rect 4525 -2359 4577 -2353
rect 4525 -2393 4535 -2359
rect 4535 -2393 4569 -2359
rect 4569 -2393 4577 -2359
rect 4525 -2405 4577 -2393
rect 4729 -2359 4781 -2353
rect 4729 -2393 4737 -2359
rect 4737 -2393 4771 -2359
rect 4771 -2393 4781 -2359
rect 4729 -2405 4781 -2393
rect 4809 -2359 4861 -2353
rect 4809 -2393 4817 -2359
rect 4817 -2393 4851 -2359
rect 4851 -2393 4861 -2359
rect 4809 -2405 4861 -2393
rect 4889 -2359 4941 -2353
rect 4889 -2393 4897 -2359
rect 4897 -2393 4931 -2359
rect 4931 -2393 4941 -2359
rect 4889 -2405 4941 -2393
rect 4969 -2359 5021 -2353
rect 4969 -2393 4977 -2359
rect 4977 -2393 5011 -2359
rect 5011 -2393 5021 -2359
rect 4969 -2405 5021 -2393
rect 5049 -2359 5101 -2353
rect 5049 -2393 5057 -2359
rect 5057 -2393 5091 -2359
rect 5091 -2393 5101 -2359
rect 5049 -2405 5101 -2393
rect 5129 -2359 5181 -2353
rect 5129 -2393 5137 -2359
rect 5137 -2393 5171 -2359
rect 5171 -2393 5181 -2359
rect 5129 -2405 5181 -2393
rect 5461 -2356 5513 -2350
rect 5461 -2390 5469 -2356
rect 5469 -2390 5503 -2356
rect 5503 -2390 5513 -2356
rect 5461 -2402 5513 -2390
rect 5541 -2356 5593 -2350
rect 5541 -2390 5549 -2356
rect 5549 -2390 5583 -2356
rect 5583 -2390 5593 -2356
rect 5541 -2402 5593 -2390
rect 5621 -2356 5673 -2350
rect 5621 -2390 5629 -2356
rect 5629 -2390 5663 -2356
rect 5663 -2390 5673 -2356
rect 5621 -2402 5673 -2390
rect 5701 -2356 5753 -2350
rect 5701 -2390 5709 -2356
rect 5709 -2390 5743 -2356
rect 5743 -2390 5753 -2356
rect 5701 -2402 5753 -2390
rect 5781 -2356 5833 -2350
rect 5781 -2390 5789 -2356
rect 5789 -2390 5823 -2356
rect 5823 -2390 5833 -2356
rect 5781 -2402 5833 -2390
rect 5861 -2356 5913 -2350
rect 5861 -2390 5869 -2356
rect 5869 -2390 5903 -2356
rect 5903 -2390 5913 -2356
rect 5861 -2402 5913 -2390
rect 5959 -2411 6011 -2359
rect 6431 -2285 6483 -2274
rect 6431 -2319 6438 -2285
rect 6438 -2319 6472 -2285
rect 6472 -2319 6483 -2285
rect 6431 -2326 6483 -2319
rect 6859 -2308 6911 -2297
rect 6859 -2342 6866 -2308
rect 6866 -2342 6900 -2308
rect 6900 -2342 6911 -2308
rect 6859 -2349 6911 -2342
rect 7198 -2359 7250 -2353
rect 7198 -2393 7208 -2359
rect 7208 -2393 7242 -2359
rect 7242 -2393 7250 -2359
rect 7198 -2405 7250 -2393
rect 7278 -2359 7330 -2353
rect 7278 -2393 7288 -2359
rect 7288 -2393 7322 -2359
rect 7322 -2393 7330 -2359
rect 7278 -2405 7330 -2393
rect 7358 -2359 7410 -2353
rect 7358 -2393 7368 -2359
rect 7368 -2393 7402 -2359
rect 7402 -2393 7410 -2359
rect 7358 -2405 7410 -2393
rect 7438 -2359 7490 -2353
rect 7438 -2393 7448 -2359
rect 7448 -2393 7482 -2359
rect 7482 -2393 7490 -2359
rect 7438 -2405 7490 -2393
rect 7518 -2359 7570 -2353
rect 7518 -2393 7528 -2359
rect 7528 -2393 7562 -2359
rect 7562 -2393 7570 -2359
rect 7518 -2405 7570 -2393
rect 7598 -2359 7650 -2353
rect 7598 -2393 7608 -2359
rect 7608 -2393 7642 -2359
rect 7642 -2393 7650 -2359
rect 7598 -2405 7650 -2393
rect 7802 -2359 7854 -2353
rect 7802 -2393 7810 -2359
rect 7810 -2393 7844 -2359
rect 7844 -2393 7854 -2359
rect 7802 -2405 7854 -2393
rect 7882 -2359 7934 -2353
rect 7882 -2393 7890 -2359
rect 7890 -2393 7924 -2359
rect 7924 -2393 7934 -2359
rect 7882 -2405 7934 -2393
rect 7962 -2359 8014 -2353
rect 7962 -2393 7970 -2359
rect 7970 -2393 8004 -2359
rect 8004 -2393 8014 -2359
rect 7962 -2405 8014 -2393
rect 8042 -2359 8094 -2353
rect 8042 -2393 8050 -2359
rect 8050 -2393 8084 -2359
rect 8084 -2393 8094 -2359
rect 8042 -2405 8094 -2393
rect 8122 -2359 8174 -2353
rect 8122 -2393 8130 -2359
rect 8130 -2393 8164 -2359
rect 8164 -2393 8174 -2359
rect 8122 -2405 8174 -2393
rect 8202 -2359 8254 -2353
rect 8202 -2393 8210 -2359
rect 8210 -2393 8244 -2359
rect 8244 -2393 8254 -2359
rect 8202 -2405 8254 -2393
rect 8410 -2359 8462 -2353
rect 8410 -2393 8420 -2359
rect 8420 -2393 8454 -2359
rect 8454 -2393 8462 -2359
rect 8410 -2405 8462 -2393
rect 8490 -2359 8542 -2353
rect 8490 -2393 8500 -2359
rect 8500 -2393 8534 -2359
rect 8534 -2393 8542 -2359
rect 8490 -2405 8542 -2393
rect 8570 -2359 8622 -2353
rect 8570 -2393 8580 -2359
rect 8580 -2393 8614 -2359
rect 8614 -2393 8622 -2359
rect 8570 -2405 8622 -2393
rect 8650 -2359 8702 -2353
rect 8650 -2393 8660 -2359
rect 8660 -2393 8694 -2359
rect 8694 -2393 8702 -2359
rect 8650 -2405 8702 -2393
rect 8730 -2359 8782 -2353
rect 8730 -2393 8740 -2359
rect 8740 -2393 8774 -2359
rect 8774 -2393 8782 -2359
rect 8730 -2405 8782 -2393
rect 8810 -2359 8862 -2353
rect 8810 -2393 8820 -2359
rect 8820 -2393 8854 -2359
rect 8854 -2393 8862 -2359
rect 8810 -2405 8862 -2393
rect 9014 -2359 9066 -2353
rect 9014 -2393 9022 -2359
rect 9022 -2393 9056 -2359
rect 9056 -2393 9066 -2359
rect 9014 -2405 9066 -2393
rect 9094 -2359 9146 -2353
rect 9094 -2393 9102 -2359
rect 9102 -2393 9136 -2359
rect 9136 -2393 9146 -2359
rect 9094 -2405 9146 -2393
rect 9174 -2359 9226 -2353
rect 9174 -2393 9182 -2359
rect 9182 -2393 9216 -2359
rect 9216 -2393 9226 -2359
rect 9174 -2405 9226 -2393
rect 9254 -2359 9306 -2353
rect 9254 -2393 9262 -2359
rect 9262 -2393 9296 -2359
rect 9296 -2393 9306 -2359
rect 9254 -2405 9306 -2393
rect 9334 -2359 9386 -2353
rect 9334 -2393 9342 -2359
rect 9342 -2393 9376 -2359
rect 9376 -2393 9386 -2359
rect 9334 -2405 9386 -2393
rect 9414 -2359 9466 -2353
rect 9414 -2393 9422 -2359
rect 9422 -2393 9456 -2359
rect 9456 -2393 9466 -2359
rect 9414 -2405 9466 -2393
rect 9622 -2359 9674 -2353
rect 9622 -2393 9632 -2359
rect 9632 -2393 9666 -2359
rect 9666 -2393 9674 -2359
rect 9622 -2405 9674 -2393
rect 9702 -2359 9754 -2353
rect 9702 -2393 9712 -2359
rect 9712 -2393 9746 -2359
rect 9746 -2393 9754 -2359
rect 9702 -2405 9754 -2393
rect 9782 -2359 9834 -2353
rect 9782 -2393 9792 -2359
rect 9792 -2393 9826 -2359
rect 9826 -2393 9834 -2359
rect 9782 -2405 9834 -2393
rect 9862 -2359 9914 -2353
rect 9862 -2393 9872 -2359
rect 9872 -2393 9906 -2359
rect 9906 -2393 9914 -2359
rect 9862 -2405 9914 -2393
rect 9942 -2359 9994 -2353
rect 9942 -2393 9952 -2359
rect 9952 -2393 9986 -2359
rect 9986 -2393 9994 -2359
rect 9942 -2405 9994 -2393
rect 10022 -2359 10074 -2353
rect 10022 -2393 10032 -2359
rect 10032 -2393 10066 -2359
rect 10066 -2393 10074 -2359
rect 10022 -2405 10074 -2393
rect 10226 -2359 10278 -2353
rect 10226 -2393 10234 -2359
rect 10234 -2393 10268 -2359
rect 10268 -2393 10278 -2359
rect 10226 -2405 10278 -2393
rect 10306 -2359 10358 -2353
rect 10306 -2393 10314 -2359
rect 10314 -2393 10348 -2359
rect 10348 -2393 10358 -2359
rect 10306 -2405 10358 -2393
rect 10386 -2359 10438 -2353
rect 10386 -2393 10394 -2359
rect 10394 -2393 10428 -2359
rect 10428 -2393 10438 -2359
rect 10386 -2405 10438 -2393
rect 10466 -2359 10518 -2353
rect 10466 -2393 10474 -2359
rect 10474 -2393 10508 -2359
rect 10508 -2393 10518 -2359
rect 10466 -2405 10518 -2393
rect 10546 -2359 10598 -2353
rect 10546 -2393 10554 -2359
rect 10554 -2393 10588 -2359
rect 10588 -2393 10598 -2359
rect 10546 -2405 10598 -2393
rect 10626 -2359 10678 -2353
rect 10626 -2393 10634 -2359
rect 10634 -2393 10668 -2359
rect 10668 -2393 10678 -2359
rect 10626 -2405 10678 -2393
rect 10834 -2359 10886 -2353
rect 10834 -2393 10844 -2359
rect 10844 -2393 10878 -2359
rect 10878 -2393 10886 -2359
rect 10834 -2405 10886 -2393
rect 10914 -2359 10966 -2353
rect 10914 -2393 10924 -2359
rect 10924 -2393 10958 -2359
rect 10958 -2393 10966 -2359
rect 10914 -2405 10966 -2393
rect 10994 -2359 11046 -2353
rect 10994 -2393 11004 -2359
rect 11004 -2393 11038 -2359
rect 11038 -2393 11046 -2359
rect 10994 -2405 11046 -2393
rect 11074 -2359 11126 -2353
rect 11074 -2393 11084 -2359
rect 11084 -2393 11118 -2359
rect 11118 -2393 11126 -2359
rect 11074 -2405 11126 -2393
rect 11154 -2359 11206 -2353
rect 11154 -2393 11164 -2359
rect 11164 -2393 11198 -2359
rect 11198 -2393 11206 -2359
rect 11154 -2405 11206 -2393
rect 11234 -2359 11286 -2353
rect 11234 -2393 11244 -2359
rect 11244 -2393 11278 -2359
rect 11278 -2393 11286 -2359
rect 11234 -2405 11286 -2393
rect 11438 -2359 11490 -2353
rect 11438 -2393 11446 -2359
rect 11446 -2393 11480 -2359
rect 11480 -2393 11490 -2359
rect 11438 -2405 11490 -2393
rect 11518 -2359 11570 -2353
rect 11518 -2393 11526 -2359
rect 11526 -2393 11560 -2359
rect 11560 -2393 11570 -2359
rect 11518 -2405 11570 -2393
rect 11598 -2359 11650 -2353
rect 11598 -2393 11606 -2359
rect 11606 -2393 11640 -2359
rect 11640 -2393 11650 -2359
rect 11598 -2405 11650 -2393
rect 11678 -2359 11730 -2353
rect 11678 -2393 11686 -2359
rect 11686 -2393 11720 -2359
rect 11720 -2393 11730 -2359
rect 11678 -2405 11730 -2393
rect 11758 -2359 11810 -2353
rect 11758 -2393 11766 -2359
rect 11766 -2393 11800 -2359
rect 11800 -2393 11810 -2359
rect 11758 -2405 11810 -2393
rect 11838 -2359 11890 -2353
rect 11838 -2393 11846 -2359
rect 11846 -2393 11880 -2359
rect 11880 -2393 11890 -2359
rect 11838 -2405 11890 -2393
rect 12170 -2356 12222 -2350
rect 12170 -2390 12178 -2356
rect 12178 -2390 12212 -2356
rect 12212 -2390 12222 -2356
rect 12170 -2402 12222 -2390
rect 12250 -2356 12302 -2350
rect 12250 -2390 12258 -2356
rect 12258 -2390 12292 -2356
rect 12292 -2390 12302 -2356
rect 12250 -2402 12302 -2390
rect 12330 -2356 12382 -2350
rect 12330 -2390 12338 -2356
rect 12338 -2390 12372 -2356
rect 12372 -2390 12382 -2356
rect 12330 -2402 12382 -2390
rect 12410 -2356 12462 -2350
rect 12410 -2390 12418 -2356
rect 12418 -2390 12452 -2356
rect 12452 -2390 12462 -2356
rect 12410 -2402 12462 -2390
rect 12490 -2356 12542 -2350
rect 12490 -2390 12498 -2356
rect 12498 -2390 12532 -2356
rect 12532 -2390 12542 -2356
rect 12490 -2402 12542 -2390
rect 12570 -2356 12622 -2350
rect 12570 -2390 12578 -2356
rect 12578 -2390 12612 -2356
rect 12612 -2390 12622 -2356
rect 12570 -2402 12622 -2390
rect 12668 -2411 12720 -2359
<< metal2 >>
rect 733 3734 807 3738
rect 733 3678 742 3734
rect 798 3729 807 3734
rect 7442 3734 7516 3738
rect 798 3725 1404 3729
rect 798 3678 838 3725
rect 733 3674 838 3678
rect 734 3669 838 3674
rect 894 3669 918 3725
rect 974 3669 998 3725
rect 1054 3669 1078 3725
rect 1134 3669 1158 3725
rect 1214 3669 1238 3725
rect 1294 3669 1404 3725
rect 734 3663 1404 3669
rect 1466 3728 6374 3732
rect 1466 3672 1570 3728
rect 1626 3672 1650 3728
rect 1706 3672 1730 3728
rect 1786 3672 1810 3728
rect 1866 3672 1890 3728
rect 1946 3672 1970 3728
rect 2026 3672 2178 3728
rect 2234 3672 2258 3728
rect 2314 3672 2338 3728
rect 2394 3672 2418 3728
rect 2474 3672 2498 3728
rect 2554 3672 2578 3728
rect 2634 3672 2782 3728
rect 2838 3672 2862 3728
rect 2918 3672 2942 3728
rect 2998 3672 3022 3728
rect 3078 3672 3102 3728
rect 3158 3672 3182 3728
rect 3238 3672 3390 3728
rect 3446 3672 3470 3728
rect 3526 3672 3550 3728
rect 3606 3672 3630 3728
rect 3686 3672 3710 3728
rect 3766 3672 3790 3728
rect 3846 3672 3994 3728
rect 4050 3672 4074 3728
rect 4130 3672 4154 3728
rect 4210 3672 4234 3728
rect 4290 3672 4314 3728
rect 4370 3672 4394 3728
rect 4450 3672 4602 3728
rect 4658 3672 4682 3728
rect 4738 3672 4762 3728
rect 4818 3672 4842 3728
rect 4898 3672 4922 3728
rect 4978 3672 5002 3728
rect 5058 3672 5206 3728
rect 5262 3672 5286 3728
rect 5342 3672 5366 3728
rect 5422 3672 5446 3728
rect 5502 3672 5526 3728
rect 5582 3672 5606 3728
rect 5662 3672 5814 3728
rect 5870 3672 5894 3728
rect 5950 3672 5974 3728
rect 6030 3672 6054 3728
rect 6110 3672 6134 3728
rect 6190 3672 6214 3728
rect 6270 3672 6374 3728
rect 1466 3666 6374 3672
rect 6542 3672 6616 3676
rect 6542 3616 6551 3672
rect 6607 3616 6616 3672
rect 6542 3612 6616 3616
rect 7019 3675 7093 3679
rect 7019 3619 7028 3675
rect 7084 3619 7093 3675
rect 7442 3678 7451 3734
rect 7507 3729 7516 3734
rect 7507 3725 8113 3729
rect 7507 3678 7547 3725
rect 7442 3674 7547 3678
rect 7443 3669 7547 3674
rect 7603 3669 7627 3725
rect 7683 3669 7707 3725
rect 7763 3669 7787 3725
rect 7843 3669 7867 3725
rect 7923 3669 7947 3725
rect 8003 3669 8113 3725
rect 7443 3663 8113 3669
rect 8175 3728 13083 3732
rect 8175 3672 8279 3728
rect 8335 3672 8359 3728
rect 8415 3672 8439 3728
rect 8495 3672 8519 3728
rect 8575 3672 8599 3728
rect 8655 3672 8679 3728
rect 8735 3672 8887 3728
rect 8943 3672 8967 3728
rect 9023 3672 9047 3728
rect 9103 3672 9127 3728
rect 9183 3672 9207 3728
rect 9263 3672 9287 3728
rect 9343 3672 9491 3728
rect 9547 3672 9571 3728
rect 9627 3672 9651 3728
rect 9707 3672 9731 3728
rect 9787 3672 9811 3728
rect 9867 3672 9891 3728
rect 9947 3672 10099 3728
rect 10155 3672 10179 3728
rect 10235 3672 10259 3728
rect 10315 3672 10339 3728
rect 10395 3672 10419 3728
rect 10475 3672 10499 3728
rect 10555 3672 10703 3728
rect 10759 3672 10783 3728
rect 10839 3672 10863 3728
rect 10919 3672 10943 3728
rect 10999 3672 11023 3728
rect 11079 3672 11103 3728
rect 11159 3672 11311 3728
rect 11367 3672 11391 3728
rect 11447 3672 11471 3728
rect 11527 3672 11551 3728
rect 11607 3672 11631 3728
rect 11687 3672 11711 3728
rect 11767 3672 11915 3728
rect 11971 3672 11995 3728
rect 12051 3672 12075 3728
rect 12131 3672 12155 3728
rect 12211 3672 12235 3728
rect 12291 3672 12315 3728
rect 12371 3672 12523 3728
rect 12579 3672 12603 3728
rect 12659 3672 12683 3728
rect 12739 3672 12763 3728
rect 12819 3672 12843 3728
rect 12899 3672 12923 3728
rect 12979 3672 13083 3728
rect 8175 3666 13083 3672
rect 13251 3672 13325 3676
rect 7019 3615 7093 3619
rect 13251 3616 13260 3672
rect 13316 3616 13325 3672
rect 13251 3612 13325 3616
rect 6547 3528 6621 3532
rect 6547 3472 6556 3528
rect 6612 3472 6621 3528
rect 13256 3528 13330 3532
rect 6547 3468 6621 3472
rect 7008 3503 7082 3507
rect 7008 3447 7017 3503
rect 7073 3447 7082 3503
rect 13256 3472 13265 3528
rect 13321 3472 13330 3528
rect 13256 3468 13330 3472
rect 7008 3443 7082 3447
rect 6548 3376 6622 3380
rect 6548 3320 6557 3376
rect 6613 3320 6622 3376
rect 6548 3316 6622 3320
rect 13257 3376 13331 3380
rect 13257 3320 13266 3376
rect 13322 3320 13331 3376
rect 13257 3316 13331 3320
rect 7008 3311 7082 3315
rect 7008 3255 7017 3311
rect 7073 3255 7082 3311
rect 7008 3251 7082 3255
rect 6548 3206 6622 3210
rect 6548 3150 6557 3206
rect 6613 3150 6622 3206
rect 6548 3146 6622 3150
rect 13257 3206 13331 3210
rect 13257 3150 13266 3206
rect 13322 3150 13331 3206
rect 13257 3146 13331 3150
rect 125 3129 181 3138
rect 125 3064 181 3073
rect 256 3128 312 3137
rect 256 3063 312 3072
rect 400 3129 456 3138
rect 400 3064 456 3073
rect 6834 3129 6890 3138
rect 6834 3064 6890 3073
rect 6965 3128 7021 3137
rect 6965 3063 7021 3072
rect 7109 3129 7165 3138
rect 7109 3064 7165 3073
rect 6547 3049 6621 3053
rect 6547 2993 6556 3049
rect 6612 2993 6621 3049
rect 6547 2989 6621 2993
rect 13256 3049 13330 3053
rect 13256 2993 13265 3049
rect 13321 2993 13330 3049
rect 13256 2989 13330 2993
rect 392 2764 400 2816
rect 452 2764 458 2816
rect 392 2763 458 2764
rect 6465 2807 6539 2811
rect 410 2687 456 2763
rect 6465 2751 6474 2807
rect 6530 2751 6539 2807
rect 7101 2764 7109 2816
rect 7161 2764 7167 2816
rect 7101 2763 7167 2764
rect 13174 2807 13248 2811
rect 6465 2747 6539 2751
rect 7119 2687 7165 2763
rect 13174 2751 13183 2807
rect 13239 2751 13248 2807
rect 13174 2747 13248 2751
rect 410 2641 649 2687
rect 7119 2641 7358 2687
rect 143 2583 199 2592
rect 143 2518 199 2527
rect 263 2583 319 2592
rect 263 2518 319 2527
rect 406 2583 462 2592
rect 406 2518 462 2527
rect 406 2238 471 2239
rect 406 2186 412 2238
rect 464 2235 471 2238
rect 603 2235 649 2641
rect 6852 2583 6908 2592
rect 1949 2548 2028 2549
rect 2176 2548 2255 2549
rect 3161 2548 3240 2549
rect 3388 2548 3467 2549
rect 4373 2548 4452 2549
rect 4600 2548 4679 2549
rect 5585 2548 5664 2549
rect 5812 2548 5891 2549
rect 1217 2545 1296 2546
rect 1214 2481 1224 2545
rect 1288 2481 1297 2545
rect 1946 2484 1956 2548
rect 2020 2484 2029 2548
rect 2175 2484 2184 2548
rect 2248 2484 2258 2548
rect 3158 2484 3168 2548
rect 3232 2484 3241 2548
rect 3387 2484 3396 2548
rect 3460 2484 3470 2548
rect 4370 2484 4380 2548
rect 4444 2484 4453 2548
rect 4599 2484 4608 2548
rect 4672 2484 4682 2548
rect 5582 2484 5592 2548
rect 5656 2484 5665 2548
rect 5811 2484 5820 2548
rect 5884 2484 5894 2548
rect 6553 2546 6627 2550
rect 6553 2490 6562 2546
rect 6618 2490 6627 2546
rect 6852 2518 6908 2527
rect 6972 2583 7028 2592
rect 6972 2518 7028 2527
rect 7115 2583 7171 2592
rect 7115 2518 7171 2527
rect 6553 2486 6627 2490
rect 1571 2282 1580 2346
rect 1644 2282 1653 2346
rect 1571 2281 1653 2282
rect 2303 2282 2312 2346
rect 2376 2282 2385 2346
rect 2303 2281 2385 2282
rect 2521 2282 2530 2346
rect 2594 2282 2603 2346
rect 2521 2281 2603 2282
rect 3515 2282 3524 2346
rect 3588 2282 3597 2346
rect 3515 2281 3597 2282
rect 3733 2282 3742 2346
rect 3806 2282 3815 2346
rect 3733 2281 3815 2282
rect 4853 2282 4862 2346
rect 4926 2282 4935 2346
rect 4853 2281 4935 2282
rect 5071 2282 5080 2346
rect 5144 2282 5153 2346
rect 5071 2281 5153 2282
rect 5805 2282 5814 2346
rect 5878 2282 5887 2346
rect 6553 2343 6627 2347
rect 6553 2287 6562 2343
rect 6618 2287 6627 2343
rect 6553 2283 6627 2287
rect 5805 2281 5887 2282
rect 7115 2238 7180 2239
rect 893 2235 900 2238
rect 464 2189 900 2235
rect 464 2186 471 2189
rect 893 2186 900 2189
rect 952 2186 958 2238
rect 7115 2186 7121 2238
rect 7173 2235 7180 2238
rect 7312 2235 7358 2641
rect 8658 2548 8737 2549
rect 8885 2548 8964 2549
rect 9870 2548 9949 2549
rect 10097 2548 10176 2549
rect 11082 2548 11161 2549
rect 11309 2548 11388 2549
rect 12294 2548 12373 2549
rect 12521 2548 12600 2549
rect 7926 2545 8005 2546
rect 7923 2481 7933 2545
rect 7997 2481 8006 2545
rect 8655 2484 8665 2548
rect 8729 2484 8738 2548
rect 8884 2484 8893 2548
rect 8957 2484 8967 2548
rect 9867 2484 9877 2548
rect 9941 2484 9950 2548
rect 10096 2484 10105 2548
rect 10169 2484 10179 2548
rect 11079 2484 11089 2548
rect 11153 2484 11162 2548
rect 11308 2484 11317 2548
rect 11381 2484 11391 2548
rect 12291 2484 12301 2548
rect 12365 2484 12374 2548
rect 12520 2484 12529 2548
rect 12593 2484 12603 2548
rect 13262 2546 13336 2550
rect 13262 2490 13271 2546
rect 13327 2490 13336 2546
rect 13262 2486 13336 2490
rect 8280 2282 8289 2346
rect 8353 2282 8362 2346
rect 8280 2281 8362 2282
rect 9012 2282 9021 2346
rect 9085 2282 9094 2346
rect 9012 2281 9094 2282
rect 9230 2282 9239 2346
rect 9303 2282 9312 2346
rect 9230 2281 9312 2282
rect 10224 2282 10233 2346
rect 10297 2282 10306 2346
rect 10224 2281 10306 2282
rect 10442 2282 10451 2346
rect 10515 2282 10524 2346
rect 10442 2281 10524 2282
rect 11562 2282 11571 2346
rect 11635 2282 11644 2346
rect 11562 2281 11644 2282
rect 11780 2282 11789 2346
rect 11853 2282 11862 2346
rect 11780 2281 11862 2282
rect 12514 2282 12523 2346
rect 12587 2282 12596 2346
rect 13262 2343 13336 2347
rect 13262 2287 13271 2343
rect 13327 2287 13336 2343
rect 13262 2283 13336 2287
rect 12514 2281 12596 2282
rect 7602 2235 7609 2238
rect 7173 2189 7609 2235
rect 7173 2186 7180 2189
rect 7602 2186 7609 2189
rect 7661 2186 7667 2238
rect 893 2185 958 2186
rect 7602 2185 7667 2186
rect 72 1701 199 1716
rect 72 1643 102 1701
rect 169 1643 199 1701
rect 72 1625 199 1643
rect 719 1156 793 1160
rect 719 1100 728 1156
rect 784 1100 793 1156
rect 719 1096 793 1100
rect 900 687 952 2185
rect 6462 2081 6536 2085
rect 6462 2025 6471 2081
rect 6527 2025 6536 2081
rect 6462 2021 6536 2025
rect 1254 1159 1586 1163
rect 1254 1103 1270 1159
rect 1326 1103 1350 1159
rect 1406 1103 1430 1159
rect 1486 1103 1510 1159
rect 1566 1103 1586 1159
rect 1254 1095 1586 1103
rect 1986 1159 2318 1163
rect 1986 1103 2002 1159
rect 2058 1103 2082 1159
rect 2138 1103 2162 1159
rect 2218 1103 2242 1159
rect 2298 1103 2318 1159
rect 1986 1095 2318 1103
rect 2588 1159 2920 1163
rect 2588 1103 2608 1159
rect 2664 1103 2688 1159
rect 2744 1103 2768 1159
rect 2824 1103 2848 1159
rect 2904 1103 2920 1159
rect 2588 1095 2920 1103
rect 3198 1159 3530 1163
rect 3198 1103 3214 1159
rect 3270 1103 3294 1159
rect 3350 1103 3374 1159
rect 3430 1103 3454 1159
rect 3510 1103 3530 1159
rect 3198 1095 3530 1103
rect 3800 1159 4132 1163
rect 3800 1103 3820 1159
rect 3876 1103 3900 1159
rect 3956 1103 3980 1159
rect 4036 1103 4060 1159
rect 4116 1103 4132 1159
rect 3800 1095 4132 1103
rect 4536 1159 4868 1163
rect 4536 1103 4552 1159
rect 4608 1103 4632 1159
rect 4688 1103 4712 1159
rect 4768 1103 4792 1159
rect 4848 1103 4868 1159
rect 4536 1095 4868 1103
rect 5138 1159 5470 1163
rect 5138 1103 5158 1159
rect 5214 1103 5238 1159
rect 5294 1103 5318 1159
rect 5374 1103 5398 1159
rect 5454 1103 5470 1159
rect 5138 1095 5470 1103
rect 5872 1159 6204 1163
rect 5872 1103 5892 1159
rect 5948 1103 5972 1159
rect 6028 1103 6052 1159
rect 6108 1103 6132 1159
rect 6188 1103 6204 1159
rect 5872 1095 6204 1103
rect 7428 1156 7502 1160
rect 7428 1100 7437 1156
rect 7493 1100 7502 1156
rect 7428 1096 7502 1100
rect 891 684 961 687
rect 891 632 900 684
rect 952 632 961 684
rect 7609 681 7661 2185
rect 13171 2081 13245 2085
rect 13171 2025 13180 2081
rect 13236 2025 13245 2081
rect 13171 2021 13245 2025
rect 7963 1159 8295 1163
rect 7963 1103 7979 1159
rect 8035 1103 8059 1159
rect 8115 1103 8139 1159
rect 8195 1103 8219 1159
rect 8275 1103 8295 1159
rect 7963 1095 8295 1103
rect 8695 1159 9027 1163
rect 8695 1103 8711 1159
rect 8767 1103 8791 1159
rect 8847 1103 8871 1159
rect 8927 1103 8951 1159
rect 9007 1103 9027 1159
rect 8695 1095 9027 1103
rect 9297 1159 9629 1163
rect 9297 1103 9317 1159
rect 9373 1103 9397 1159
rect 9453 1103 9477 1159
rect 9533 1103 9557 1159
rect 9613 1103 9629 1159
rect 9297 1095 9629 1103
rect 9907 1159 10239 1163
rect 9907 1103 9923 1159
rect 9979 1103 10003 1159
rect 10059 1103 10083 1159
rect 10139 1103 10163 1159
rect 10219 1103 10239 1159
rect 9907 1095 10239 1103
rect 10509 1159 10841 1163
rect 10509 1103 10529 1159
rect 10585 1103 10609 1159
rect 10665 1103 10689 1159
rect 10745 1103 10769 1159
rect 10825 1103 10841 1159
rect 10509 1095 10841 1103
rect 11245 1159 11577 1163
rect 11245 1103 11261 1159
rect 11317 1103 11341 1159
rect 11397 1103 11421 1159
rect 11477 1103 11501 1159
rect 11557 1103 11577 1159
rect 11245 1095 11577 1103
rect 11847 1159 12179 1163
rect 11847 1103 11867 1159
rect 11923 1103 11947 1159
rect 12003 1103 12027 1159
rect 12083 1103 12107 1159
rect 12163 1103 12179 1159
rect 11847 1095 12179 1103
rect 12581 1159 12913 1163
rect 12581 1103 12601 1159
rect 12657 1103 12681 1159
rect 12737 1103 12761 1159
rect 12817 1103 12841 1159
rect 12897 1103 12913 1159
rect 12581 1095 12913 1103
rect 12498 685 12574 686
rect 891 624 961 632
rect 5791 674 5861 681
rect 5791 622 5800 674
rect 5853 622 5861 674
rect 7602 677 7670 681
rect 7602 624 7609 677
rect 7661 624 7670 677
rect 5791 614 5861 622
rect 12498 621 12504 685
rect 12568 621 12574 685
rect 551 218 883 226
rect 551 162 567 218
rect 623 162 647 218
rect 703 162 727 218
rect 783 162 807 218
rect 863 162 883 218
rect 551 158 883 162
rect 1285 218 1617 226
rect 1285 162 1301 218
rect 1357 162 1381 218
rect 1437 162 1461 218
rect 1517 162 1541 218
rect 1597 162 1617 218
rect 1285 158 1617 162
rect 1887 218 2219 226
rect 1887 162 1907 218
rect 1963 162 1987 218
rect 2043 162 2067 218
rect 2123 162 2147 218
rect 2203 162 2219 218
rect 1887 158 2219 162
rect 2623 218 2955 226
rect 2623 162 2639 218
rect 2695 162 2719 218
rect 2775 162 2799 218
rect 2855 162 2879 218
rect 2935 162 2955 218
rect 2623 158 2955 162
rect 3225 218 3557 226
rect 3225 162 3245 218
rect 3301 162 3325 218
rect 3381 162 3405 218
rect 3461 162 3485 218
rect 3541 162 3557 218
rect 3225 158 3557 162
rect 3835 218 4167 226
rect 3835 162 3851 218
rect 3907 162 3931 218
rect 3987 162 4011 218
rect 4067 162 4091 218
rect 4147 162 4167 218
rect 3835 158 4167 162
rect 4437 218 4769 226
rect 4437 162 4457 218
rect 4513 162 4537 218
rect 4593 162 4617 218
rect 4673 162 4697 218
rect 4753 162 4769 218
rect 4437 158 4769 162
rect 5169 218 5501 226
rect 5169 162 5189 218
rect 5245 162 5269 218
rect 5325 162 5349 218
rect 5405 162 5429 218
rect 5485 162 5501 218
rect 5169 158 5501 162
rect 219 -704 293 -700
rect 219 -760 228 -704
rect 284 -760 293 -704
rect 219 -764 293 -760
rect 5799 -864 5851 614
rect 5962 221 6036 225
rect 5962 165 5971 221
rect 6027 165 6036 221
rect 5962 161 6036 165
rect 7260 218 7592 226
rect 7260 162 7276 218
rect 7332 162 7356 218
rect 7412 162 7436 218
rect 7492 162 7516 218
rect 7572 162 7592 218
rect 7260 158 7592 162
rect 7994 218 8326 226
rect 7994 162 8010 218
rect 8066 162 8090 218
rect 8146 162 8170 218
rect 8226 162 8250 218
rect 8306 162 8326 218
rect 7994 158 8326 162
rect 8596 218 8928 226
rect 8596 162 8616 218
rect 8672 162 8696 218
rect 8752 162 8776 218
rect 8832 162 8856 218
rect 8912 162 8928 218
rect 8596 158 8928 162
rect 9332 218 9664 226
rect 9332 162 9348 218
rect 9404 162 9428 218
rect 9484 162 9508 218
rect 9564 162 9588 218
rect 9644 162 9664 218
rect 9332 158 9664 162
rect 9934 218 10266 226
rect 9934 162 9954 218
rect 10010 162 10034 218
rect 10090 162 10114 218
rect 10170 162 10194 218
rect 10250 162 10266 218
rect 9934 158 10266 162
rect 10544 218 10876 226
rect 10544 162 10560 218
rect 10616 162 10640 218
rect 10696 162 10720 218
rect 10776 162 10800 218
rect 10856 162 10876 218
rect 10544 158 10876 162
rect 11146 218 11478 226
rect 11146 162 11166 218
rect 11222 162 11246 218
rect 11302 162 11326 218
rect 11382 162 11406 218
rect 11462 162 11478 218
rect 11146 158 11478 162
rect 11878 218 12210 226
rect 11878 162 11898 218
rect 11954 162 11978 218
rect 12034 162 12058 218
rect 12114 162 12138 218
rect 12194 162 12210 218
rect 11878 158 12210 162
rect 6928 -704 7002 -700
rect 6928 -760 6937 -704
rect 6993 -760 7002 -704
rect 6928 -764 7002 -760
rect 12511 -864 12563 621
rect 12671 221 12745 225
rect 12671 165 12680 221
rect 12736 165 12745 221
rect 12671 161 12745 165
rect 5797 -865 5862 -864
rect 12506 -865 12571 -864
rect 5797 -917 5803 -865
rect 5855 -868 5862 -865
rect 6284 -868 6291 -865
rect 5855 -914 6291 -868
rect 5855 -917 5862 -914
rect 868 -961 950 -960
rect 128 -966 202 -962
rect 128 -1022 137 -966
rect 193 -1022 202 -966
rect 128 -1026 202 -1022
rect 868 -1025 877 -961
rect 941 -1025 950 -961
rect 1602 -961 1684 -960
rect 1602 -1025 1611 -961
rect 1675 -1025 1684 -961
rect 1820 -961 1902 -960
rect 1820 -1025 1829 -961
rect 1893 -1025 1902 -961
rect 2940 -961 3022 -960
rect 2940 -1025 2949 -961
rect 3013 -1025 3022 -961
rect 3158 -961 3240 -960
rect 3158 -1025 3167 -961
rect 3231 -1025 3240 -961
rect 4152 -961 4234 -960
rect 4152 -1025 4161 -961
rect 4225 -1025 4234 -961
rect 4370 -961 4452 -960
rect 4370 -1025 4379 -961
rect 4443 -1025 4452 -961
rect 5102 -961 5184 -960
rect 5102 -1025 5111 -961
rect 5175 -1025 5184 -961
rect 128 -1169 202 -1165
rect 128 -1225 137 -1169
rect 193 -1225 202 -1169
rect 128 -1229 202 -1225
rect 861 -1227 871 -1163
rect 935 -1227 944 -1163
rect 1090 -1227 1099 -1163
rect 1163 -1227 1173 -1163
rect 2073 -1227 2083 -1163
rect 2147 -1227 2156 -1163
rect 2302 -1227 2311 -1163
rect 2375 -1227 2385 -1163
rect 3285 -1227 3295 -1163
rect 3359 -1227 3368 -1163
rect 3514 -1227 3523 -1163
rect 3587 -1227 3597 -1163
rect 4497 -1227 4507 -1163
rect 4571 -1227 4580 -1163
rect 4726 -1227 4735 -1163
rect 4799 -1227 4809 -1163
rect 5458 -1224 5467 -1160
rect 5531 -1224 5541 -1160
rect 5459 -1225 5538 -1224
rect 864 -1228 943 -1227
rect 1091 -1228 1170 -1227
rect 2076 -1228 2155 -1227
rect 2303 -1228 2382 -1227
rect 3288 -1228 3367 -1227
rect 3515 -1228 3594 -1227
rect 4500 -1228 4579 -1227
rect 4727 -1228 4806 -1227
rect 6106 -1320 6152 -914
rect 6284 -917 6291 -914
rect 6343 -917 6349 -865
rect 12506 -917 12512 -865
rect 12564 -868 12571 -865
rect 12993 -868 13000 -865
rect 12564 -914 13000 -868
rect 12564 -917 12571 -914
rect 6284 -918 6349 -917
rect 7577 -961 7659 -960
rect 6837 -966 6911 -962
rect 6837 -1022 6846 -966
rect 6902 -1022 6911 -966
rect 6837 -1026 6911 -1022
rect 7577 -1025 7586 -961
rect 7650 -1025 7659 -961
rect 8311 -961 8393 -960
rect 8311 -1025 8320 -961
rect 8384 -1025 8393 -961
rect 8529 -961 8611 -960
rect 8529 -1025 8538 -961
rect 8602 -1025 8611 -961
rect 9649 -961 9731 -960
rect 9649 -1025 9658 -961
rect 9722 -1025 9731 -961
rect 9867 -961 9949 -960
rect 9867 -1025 9876 -961
rect 9940 -1025 9949 -961
rect 10861 -961 10943 -960
rect 10861 -1025 10870 -961
rect 10934 -1025 10943 -961
rect 11079 -961 11161 -960
rect 11079 -1025 11088 -961
rect 11152 -1025 11161 -961
rect 11811 -961 11893 -960
rect 11811 -1025 11820 -961
rect 11884 -1025 11893 -961
rect 6837 -1169 6911 -1165
rect 6293 -1206 6349 -1197
rect 6293 -1271 6349 -1262
rect 6436 -1206 6492 -1197
rect 6436 -1271 6492 -1262
rect 6556 -1206 6612 -1197
rect 6837 -1225 6846 -1169
rect 6902 -1225 6911 -1169
rect 6837 -1229 6911 -1225
rect 7570 -1227 7580 -1163
rect 7644 -1227 7653 -1163
rect 7799 -1227 7808 -1163
rect 7872 -1227 7882 -1163
rect 8782 -1227 8792 -1163
rect 8856 -1227 8865 -1163
rect 9011 -1227 9020 -1163
rect 9084 -1227 9094 -1163
rect 9994 -1227 10004 -1163
rect 10068 -1227 10077 -1163
rect 10223 -1227 10232 -1163
rect 10296 -1227 10306 -1163
rect 11206 -1227 11216 -1163
rect 11280 -1227 11289 -1163
rect 11435 -1227 11444 -1163
rect 11508 -1227 11518 -1163
rect 12167 -1224 12176 -1160
rect 12240 -1224 12250 -1160
rect 12168 -1225 12247 -1224
rect 7573 -1228 7652 -1227
rect 7800 -1228 7879 -1227
rect 8785 -1228 8864 -1227
rect 9012 -1228 9091 -1227
rect 9997 -1228 10076 -1227
rect 10224 -1228 10303 -1227
rect 11209 -1228 11288 -1227
rect 11436 -1228 11515 -1227
rect 6556 -1271 6612 -1262
rect 12815 -1320 12861 -914
rect 12993 -917 13000 -914
rect 13052 -917 13058 -865
rect 12993 -918 13058 -917
rect 13002 -1206 13058 -1197
rect 13002 -1271 13058 -1262
rect 13145 -1206 13201 -1197
rect 13145 -1271 13201 -1262
rect 13265 -1206 13321 -1197
rect 13265 -1271 13321 -1262
rect 6106 -1366 6345 -1320
rect 12815 -1366 13054 -1320
rect 216 -1430 290 -1426
rect 216 -1486 225 -1430
rect 281 -1486 290 -1430
rect 6299 -1442 6345 -1366
rect 6925 -1430 6999 -1426
rect 216 -1490 290 -1486
rect 6297 -1443 6363 -1442
rect 6297 -1495 6303 -1443
rect 6355 -1495 6363 -1443
rect 6925 -1486 6934 -1430
rect 6990 -1486 6999 -1430
rect 13008 -1442 13054 -1366
rect 6925 -1490 6999 -1486
rect 13006 -1443 13072 -1442
rect 13006 -1495 13012 -1443
rect 13064 -1495 13072 -1443
rect 134 -1672 208 -1668
rect 134 -1728 143 -1672
rect 199 -1728 208 -1672
rect 134 -1732 208 -1728
rect 6843 -1672 6917 -1668
rect 6843 -1728 6852 -1672
rect 6908 -1728 6917 -1672
rect 6843 -1732 6917 -1728
rect 6299 -1752 6355 -1743
rect 6299 -1817 6355 -1808
rect 6443 -1751 6499 -1742
rect 6443 -1816 6499 -1807
rect 6574 -1752 6630 -1743
rect 6574 -1817 6630 -1808
rect 13008 -1752 13064 -1743
rect 13008 -1817 13064 -1808
rect 13152 -1751 13208 -1742
rect 13152 -1816 13208 -1807
rect 13283 -1752 13339 -1743
rect 13283 -1817 13339 -1808
rect 133 -1829 207 -1825
rect 133 -1885 142 -1829
rect 198 -1885 207 -1829
rect 133 -1889 207 -1885
rect 6842 -1829 6916 -1825
rect 6842 -1885 6851 -1829
rect 6907 -1885 6916 -1829
rect 6842 -1889 6916 -1885
rect 6420 -1901 6494 -1897
rect 6420 -1957 6429 -1901
rect 6485 -1957 6494 -1901
rect 6420 -1961 6494 -1957
rect 133 -1999 207 -1995
rect 133 -2055 142 -1999
rect 198 -2055 207 -1999
rect 133 -2059 207 -2055
rect 6842 -1999 6916 -1995
rect 6842 -2055 6851 -1999
rect 6907 -2055 6916 -1999
rect 6842 -2059 6916 -2055
rect 6420 -2097 6494 -2093
rect 134 -2151 208 -2147
rect 134 -2207 143 -2151
rect 199 -2207 208 -2151
rect 6420 -2153 6429 -2097
rect 6485 -2153 6494 -2097
rect 6420 -2157 6494 -2153
rect 6843 -2151 6917 -2147
rect 134 -2211 208 -2207
rect 6843 -2207 6852 -2151
rect 6908 -2207 6917 -2151
rect 6843 -2211 6917 -2207
rect 6420 -2272 6494 -2268
rect 139 -2295 213 -2291
rect 139 -2351 148 -2295
rect 204 -2351 213 -2295
rect 6420 -2328 6429 -2272
rect 6485 -2328 6494 -2272
rect 6420 -2332 6494 -2328
rect 6848 -2295 6922 -2291
rect 139 -2355 213 -2351
rect 381 -2351 5289 -2345
rect 381 -2407 485 -2351
rect 541 -2407 565 -2351
rect 621 -2407 645 -2351
rect 701 -2407 725 -2351
rect 781 -2407 805 -2351
rect 861 -2407 885 -2351
rect 941 -2407 1093 -2351
rect 1149 -2407 1173 -2351
rect 1229 -2407 1253 -2351
rect 1309 -2407 1333 -2351
rect 1389 -2407 1413 -2351
rect 1469 -2407 1493 -2351
rect 1549 -2407 1697 -2351
rect 1753 -2407 1777 -2351
rect 1833 -2407 1857 -2351
rect 1913 -2407 1937 -2351
rect 1993 -2407 2017 -2351
rect 2073 -2407 2097 -2351
rect 2153 -2407 2305 -2351
rect 2361 -2407 2385 -2351
rect 2441 -2407 2465 -2351
rect 2521 -2407 2545 -2351
rect 2601 -2407 2625 -2351
rect 2681 -2407 2705 -2351
rect 2761 -2407 2909 -2351
rect 2965 -2407 2989 -2351
rect 3045 -2407 3069 -2351
rect 3125 -2407 3149 -2351
rect 3205 -2407 3229 -2351
rect 3285 -2407 3309 -2351
rect 3365 -2407 3517 -2351
rect 3573 -2407 3597 -2351
rect 3653 -2407 3677 -2351
rect 3733 -2407 3757 -2351
rect 3813 -2407 3837 -2351
rect 3893 -2407 3917 -2351
rect 3973 -2407 4121 -2351
rect 4177 -2407 4201 -2351
rect 4257 -2407 4281 -2351
rect 4337 -2407 4361 -2351
rect 4417 -2407 4441 -2351
rect 4497 -2407 4521 -2351
rect 4577 -2407 4729 -2351
rect 4785 -2407 4809 -2351
rect 4865 -2407 4889 -2351
rect 4945 -2407 4969 -2351
rect 5025 -2407 5049 -2351
rect 5105 -2407 5129 -2351
rect 5185 -2407 5289 -2351
rect 381 -2411 5289 -2407
rect 5351 -2348 6021 -2342
rect 5351 -2404 5461 -2348
rect 5517 -2404 5541 -2348
rect 5597 -2404 5621 -2348
rect 5677 -2404 5701 -2348
rect 5757 -2404 5781 -2348
rect 5837 -2404 5861 -2348
rect 5917 -2353 6021 -2348
rect 6848 -2351 6857 -2295
rect 6913 -2351 6922 -2295
rect 5917 -2357 6022 -2353
rect 6848 -2355 6922 -2351
rect 7090 -2351 11998 -2345
rect 5917 -2404 5957 -2357
rect 5351 -2408 5957 -2404
rect 5948 -2413 5957 -2408
rect 6013 -2413 6022 -2357
rect 7090 -2407 7194 -2351
rect 7250 -2407 7274 -2351
rect 7330 -2407 7354 -2351
rect 7410 -2407 7434 -2351
rect 7490 -2407 7514 -2351
rect 7570 -2407 7594 -2351
rect 7650 -2407 7802 -2351
rect 7858 -2407 7882 -2351
rect 7938 -2407 7962 -2351
rect 8018 -2407 8042 -2351
rect 8098 -2407 8122 -2351
rect 8178 -2407 8202 -2351
rect 8258 -2407 8406 -2351
rect 8462 -2407 8486 -2351
rect 8542 -2407 8566 -2351
rect 8622 -2407 8646 -2351
rect 8702 -2407 8726 -2351
rect 8782 -2407 8806 -2351
rect 8862 -2407 9014 -2351
rect 9070 -2407 9094 -2351
rect 9150 -2407 9174 -2351
rect 9230 -2407 9254 -2351
rect 9310 -2407 9334 -2351
rect 9390 -2407 9414 -2351
rect 9470 -2407 9618 -2351
rect 9674 -2407 9698 -2351
rect 9754 -2407 9778 -2351
rect 9834 -2407 9858 -2351
rect 9914 -2407 9938 -2351
rect 9994 -2407 10018 -2351
rect 10074 -2407 10226 -2351
rect 10282 -2407 10306 -2351
rect 10362 -2407 10386 -2351
rect 10442 -2407 10466 -2351
rect 10522 -2407 10546 -2351
rect 10602 -2407 10626 -2351
rect 10682 -2407 10830 -2351
rect 10886 -2407 10910 -2351
rect 10966 -2407 10990 -2351
rect 11046 -2407 11070 -2351
rect 11126 -2407 11150 -2351
rect 11206 -2407 11230 -2351
rect 11286 -2407 11438 -2351
rect 11494 -2407 11518 -2351
rect 11574 -2407 11598 -2351
rect 11654 -2407 11678 -2351
rect 11734 -2407 11758 -2351
rect 11814 -2407 11838 -2351
rect 11894 -2407 11998 -2351
rect 7090 -2411 11998 -2407
rect 12060 -2348 12730 -2342
rect 12060 -2404 12170 -2348
rect 12226 -2404 12250 -2348
rect 12306 -2404 12330 -2348
rect 12386 -2404 12410 -2348
rect 12466 -2404 12490 -2348
rect 12546 -2404 12570 -2348
rect 12626 -2353 12730 -2348
rect 12626 -2357 12731 -2353
rect 12626 -2404 12666 -2357
rect 12060 -2408 12666 -2404
rect 5948 -2417 6022 -2413
rect 12657 -2413 12666 -2408
rect 12722 -2413 12731 -2357
rect 12657 -2417 12731 -2413
<< via2 >>
rect 742 3732 798 3734
rect 742 3680 744 3732
rect 744 3680 796 3732
rect 796 3680 798 3732
rect 742 3678 798 3680
rect 838 3723 894 3725
rect 838 3671 842 3723
rect 842 3671 894 3723
rect 838 3669 894 3671
rect 918 3723 974 3725
rect 918 3671 922 3723
rect 922 3671 974 3723
rect 918 3669 974 3671
rect 998 3723 1054 3725
rect 998 3671 1002 3723
rect 1002 3671 1054 3723
rect 998 3669 1054 3671
rect 1078 3723 1134 3725
rect 1078 3671 1082 3723
rect 1082 3671 1134 3723
rect 1078 3669 1134 3671
rect 1158 3723 1214 3725
rect 1158 3671 1162 3723
rect 1162 3671 1214 3723
rect 1158 3669 1214 3671
rect 1238 3723 1294 3725
rect 1238 3671 1242 3723
rect 1242 3671 1294 3723
rect 1238 3669 1294 3671
rect 1570 3726 1626 3728
rect 1570 3674 1574 3726
rect 1574 3674 1626 3726
rect 1570 3672 1626 3674
rect 1650 3726 1706 3728
rect 1650 3674 1654 3726
rect 1654 3674 1706 3726
rect 1650 3672 1706 3674
rect 1730 3726 1786 3728
rect 1730 3674 1734 3726
rect 1734 3674 1786 3726
rect 1730 3672 1786 3674
rect 1810 3726 1866 3728
rect 1810 3674 1814 3726
rect 1814 3674 1866 3726
rect 1810 3672 1866 3674
rect 1890 3726 1946 3728
rect 1890 3674 1894 3726
rect 1894 3674 1946 3726
rect 1890 3672 1946 3674
rect 1970 3726 2026 3728
rect 1970 3674 1974 3726
rect 1974 3674 2026 3726
rect 1970 3672 2026 3674
rect 2178 3726 2234 3728
rect 2178 3674 2230 3726
rect 2230 3674 2234 3726
rect 2178 3672 2234 3674
rect 2258 3726 2314 3728
rect 2258 3674 2310 3726
rect 2310 3674 2314 3726
rect 2258 3672 2314 3674
rect 2338 3726 2394 3728
rect 2338 3674 2390 3726
rect 2390 3674 2394 3726
rect 2338 3672 2394 3674
rect 2418 3726 2474 3728
rect 2418 3674 2470 3726
rect 2470 3674 2474 3726
rect 2418 3672 2474 3674
rect 2498 3726 2554 3728
rect 2498 3674 2550 3726
rect 2550 3674 2554 3726
rect 2498 3672 2554 3674
rect 2578 3726 2634 3728
rect 2578 3674 2630 3726
rect 2630 3674 2634 3726
rect 2578 3672 2634 3674
rect 2782 3726 2838 3728
rect 2782 3674 2786 3726
rect 2786 3674 2838 3726
rect 2782 3672 2838 3674
rect 2862 3726 2918 3728
rect 2862 3674 2866 3726
rect 2866 3674 2918 3726
rect 2862 3672 2918 3674
rect 2942 3726 2998 3728
rect 2942 3674 2946 3726
rect 2946 3674 2998 3726
rect 2942 3672 2998 3674
rect 3022 3726 3078 3728
rect 3022 3674 3026 3726
rect 3026 3674 3078 3726
rect 3022 3672 3078 3674
rect 3102 3726 3158 3728
rect 3102 3674 3106 3726
rect 3106 3674 3158 3726
rect 3102 3672 3158 3674
rect 3182 3726 3238 3728
rect 3182 3674 3186 3726
rect 3186 3674 3238 3726
rect 3182 3672 3238 3674
rect 3390 3726 3446 3728
rect 3390 3674 3442 3726
rect 3442 3674 3446 3726
rect 3390 3672 3446 3674
rect 3470 3726 3526 3728
rect 3470 3674 3522 3726
rect 3522 3674 3526 3726
rect 3470 3672 3526 3674
rect 3550 3726 3606 3728
rect 3550 3674 3602 3726
rect 3602 3674 3606 3726
rect 3550 3672 3606 3674
rect 3630 3726 3686 3728
rect 3630 3674 3682 3726
rect 3682 3674 3686 3726
rect 3630 3672 3686 3674
rect 3710 3726 3766 3728
rect 3710 3674 3762 3726
rect 3762 3674 3766 3726
rect 3710 3672 3766 3674
rect 3790 3726 3846 3728
rect 3790 3674 3842 3726
rect 3842 3674 3846 3726
rect 3790 3672 3846 3674
rect 3994 3726 4050 3728
rect 3994 3674 3998 3726
rect 3998 3674 4050 3726
rect 3994 3672 4050 3674
rect 4074 3726 4130 3728
rect 4074 3674 4078 3726
rect 4078 3674 4130 3726
rect 4074 3672 4130 3674
rect 4154 3726 4210 3728
rect 4154 3674 4158 3726
rect 4158 3674 4210 3726
rect 4154 3672 4210 3674
rect 4234 3726 4290 3728
rect 4234 3674 4238 3726
rect 4238 3674 4290 3726
rect 4234 3672 4290 3674
rect 4314 3726 4370 3728
rect 4314 3674 4318 3726
rect 4318 3674 4370 3726
rect 4314 3672 4370 3674
rect 4394 3726 4450 3728
rect 4394 3674 4398 3726
rect 4398 3674 4450 3726
rect 4394 3672 4450 3674
rect 4602 3726 4658 3728
rect 4602 3674 4654 3726
rect 4654 3674 4658 3726
rect 4602 3672 4658 3674
rect 4682 3726 4738 3728
rect 4682 3674 4734 3726
rect 4734 3674 4738 3726
rect 4682 3672 4738 3674
rect 4762 3726 4818 3728
rect 4762 3674 4814 3726
rect 4814 3674 4818 3726
rect 4762 3672 4818 3674
rect 4842 3726 4898 3728
rect 4842 3674 4894 3726
rect 4894 3674 4898 3726
rect 4842 3672 4898 3674
rect 4922 3726 4978 3728
rect 4922 3674 4974 3726
rect 4974 3674 4978 3726
rect 4922 3672 4978 3674
rect 5002 3726 5058 3728
rect 5002 3674 5054 3726
rect 5054 3674 5058 3726
rect 5002 3672 5058 3674
rect 5206 3726 5262 3728
rect 5206 3674 5210 3726
rect 5210 3674 5262 3726
rect 5206 3672 5262 3674
rect 5286 3726 5342 3728
rect 5286 3674 5290 3726
rect 5290 3674 5342 3726
rect 5286 3672 5342 3674
rect 5366 3726 5422 3728
rect 5366 3674 5370 3726
rect 5370 3674 5422 3726
rect 5366 3672 5422 3674
rect 5446 3726 5502 3728
rect 5446 3674 5450 3726
rect 5450 3674 5502 3726
rect 5446 3672 5502 3674
rect 5526 3726 5582 3728
rect 5526 3674 5530 3726
rect 5530 3674 5582 3726
rect 5526 3672 5582 3674
rect 5606 3726 5662 3728
rect 5606 3674 5610 3726
rect 5610 3674 5662 3726
rect 5606 3672 5662 3674
rect 5814 3726 5870 3728
rect 5814 3674 5866 3726
rect 5866 3674 5870 3726
rect 5814 3672 5870 3674
rect 5894 3726 5950 3728
rect 5894 3674 5946 3726
rect 5946 3674 5950 3726
rect 5894 3672 5950 3674
rect 5974 3726 6030 3728
rect 5974 3674 6026 3726
rect 6026 3674 6030 3726
rect 5974 3672 6030 3674
rect 6054 3726 6110 3728
rect 6054 3674 6106 3726
rect 6106 3674 6110 3726
rect 6054 3672 6110 3674
rect 6134 3726 6190 3728
rect 6134 3674 6186 3726
rect 6186 3674 6190 3726
rect 6134 3672 6190 3674
rect 6214 3726 6270 3728
rect 6214 3674 6266 3726
rect 6266 3674 6270 3726
rect 6214 3672 6270 3674
rect 6551 3670 6607 3672
rect 6551 3618 6553 3670
rect 6553 3618 6605 3670
rect 6605 3618 6607 3670
rect 6551 3616 6607 3618
rect 7028 3673 7084 3675
rect 7028 3621 7030 3673
rect 7030 3621 7082 3673
rect 7082 3621 7084 3673
rect 7028 3619 7084 3621
rect 7451 3732 7507 3734
rect 7451 3680 7453 3732
rect 7453 3680 7505 3732
rect 7505 3680 7507 3732
rect 7451 3678 7507 3680
rect 7547 3723 7603 3725
rect 7547 3671 7551 3723
rect 7551 3671 7603 3723
rect 7547 3669 7603 3671
rect 7627 3723 7683 3725
rect 7627 3671 7631 3723
rect 7631 3671 7683 3723
rect 7627 3669 7683 3671
rect 7707 3723 7763 3725
rect 7707 3671 7711 3723
rect 7711 3671 7763 3723
rect 7707 3669 7763 3671
rect 7787 3723 7843 3725
rect 7787 3671 7791 3723
rect 7791 3671 7843 3723
rect 7787 3669 7843 3671
rect 7867 3723 7923 3725
rect 7867 3671 7871 3723
rect 7871 3671 7923 3723
rect 7867 3669 7923 3671
rect 7947 3723 8003 3725
rect 7947 3671 7951 3723
rect 7951 3671 8003 3723
rect 7947 3669 8003 3671
rect 8279 3726 8335 3728
rect 8279 3674 8283 3726
rect 8283 3674 8335 3726
rect 8279 3672 8335 3674
rect 8359 3726 8415 3728
rect 8359 3674 8363 3726
rect 8363 3674 8415 3726
rect 8359 3672 8415 3674
rect 8439 3726 8495 3728
rect 8439 3674 8443 3726
rect 8443 3674 8495 3726
rect 8439 3672 8495 3674
rect 8519 3726 8575 3728
rect 8519 3674 8523 3726
rect 8523 3674 8575 3726
rect 8519 3672 8575 3674
rect 8599 3726 8655 3728
rect 8599 3674 8603 3726
rect 8603 3674 8655 3726
rect 8599 3672 8655 3674
rect 8679 3726 8735 3728
rect 8679 3674 8683 3726
rect 8683 3674 8735 3726
rect 8679 3672 8735 3674
rect 8887 3726 8943 3728
rect 8887 3674 8939 3726
rect 8939 3674 8943 3726
rect 8887 3672 8943 3674
rect 8967 3726 9023 3728
rect 8967 3674 9019 3726
rect 9019 3674 9023 3726
rect 8967 3672 9023 3674
rect 9047 3726 9103 3728
rect 9047 3674 9099 3726
rect 9099 3674 9103 3726
rect 9047 3672 9103 3674
rect 9127 3726 9183 3728
rect 9127 3674 9179 3726
rect 9179 3674 9183 3726
rect 9127 3672 9183 3674
rect 9207 3726 9263 3728
rect 9207 3674 9259 3726
rect 9259 3674 9263 3726
rect 9207 3672 9263 3674
rect 9287 3726 9343 3728
rect 9287 3674 9339 3726
rect 9339 3674 9343 3726
rect 9287 3672 9343 3674
rect 9491 3726 9547 3728
rect 9491 3674 9495 3726
rect 9495 3674 9547 3726
rect 9491 3672 9547 3674
rect 9571 3726 9627 3728
rect 9571 3674 9575 3726
rect 9575 3674 9627 3726
rect 9571 3672 9627 3674
rect 9651 3726 9707 3728
rect 9651 3674 9655 3726
rect 9655 3674 9707 3726
rect 9651 3672 9707 3674
rect 9731 3726 9787 3728
rect 9731 3674 9735 3726
rect 9735 3674 9787 3726
rect 9731 3672 9787 3674
rect 9811 3726 9867 3728
rect 9811 3674 9815 3726
rect 9815 3674 9867 3726
rect 9811 3672 9867 3674
rect 9891 3726 9947 3728
rect 9891 3674 9895 3726
rect 9895 3674 9947 3726
rect 9891 3672 9947 3674
rect 10099 3726 10155 3728
rect 10099 3674 10151 3726
rect 10151 3674 10155 3726
rect 10099 3672 10155 3674
rect 10179 3726 10235 3728
rect 10179 3674 10231 3726
rect 10231 3674 10235 3726
rect 10179 3672 10235 3674
rect 10259 3726 10315 3728
rect 10259 3674 10311 3726
rect 10311 3674 10315 3726
rect 10259 3672 10315 3674
rect 10339 3726 10395 3728
rect 10339 3674 10391 3726
rect 10391 3674 10395 3726
rect 10339 3672 10395 3674
rect 10419 3726 10475 3728
rect 10419 3674 10471 3726
rect 10471 3674 10475 3726
rect 10419 3672 10475 3674
rect 10499 3726 10555 3728
rect 10499 3674 10551 3726
rect 10551 3674 10555 3726
rect 10499 3672 10555 3674
rect 10703 3726 10759 3728
rect 10703 3674 10707 3726
rect 10707 3674 10759 3726
rect 10703 3672 10759 3674
rect 10783 3726 10839 3728
rect 10783 3674 10787 3726
rect 10787 3674 10839 3726
rect 10783 3672 10839 3674
rect 10863 3726 10919 3728
rect 10863 3674 10867 3726
rect 10867 3674 10919 3726
rect 10863 3672 10919 3674
rect 10943 3726 10999 3728
rect 10943 3674 10947 3726
rect 10947 3674 10999 3726
rect 10943 3672 10999 3674
rect 11023 3726 11079 3728
rect 11023 3674 11027 3726
rect 11027 3674 11079 3726
rect 11023 3672 11079 3674
rect 11103 3726 11159 3728
rect 11103 3674 11107 3726
rect 11107 3674 11159 3726
rect 11103 3672 11159 3674
rect 11311 3726 11367 3728
rect 11311 3674 11363 3726
rect 11363 3674 11367 3726
rect 11311 3672 11367 3674
rect 11391 3726 11447 3728
rect 11391 3674 11443 3726
rect 11443 3674 11447 3726
rect 11391 3672 11447 3674
rect 11471 3726 11527 3728
rect 11471 3674 11523 3726
rect 11523 3674 11527 3726
rect 11471 3672 11527 3674
rect 11551 3726 11607 3728
rect 11551 3674 11603 3726
rect 11603 3674 11607 3726
rect 11551 3672 11607 3674
rect 11631 3726 11687 3728
rect 11631 3674 11683 3726
rect 11683 3674 11687 3726
rect 11631 3672 11687 3674
rect 11711 3726 11767 3728
rect 11711 3674 11763 3726
rect 11763 3674 11767 3726
rect 11711 3672 11767 3674
rect 11915 3726 11971 3728
rect 11915 3674 11919 3726
rect 11919 3674 11971 3726
rect 11915 3672 11971 3674
rect 11995 3726 12051 3728
rect 11995 3674 11999 3726
rect 11999 3674 12051 3726
rect 11995 3672 12051 3674
rect 12075 3726 12131 3728
rect 12075 3674 12079 3726
rect 12079 3674 12131 3726
rect 12075 3672 12131 3674
rect 12155 3726 12211 3728
rect 12155 3674 12159 3726
rect 12159 3674 12211 3726
rect 12155 3672 12211 3674
rect 12235 3726 12291 3728
rect 12235 3674 12239 3726
rect 12239 3674 12291 3726
rect 12235 3672 12291 3674
rect 12315 3726 12371 3728
rect 12315 3674 12319 3726
rect 12319 3674 12371 3726
rect 12315 3672 12371 3674
rect 12523 3726 12579 3728
rect 12523 3674 12575 3726
rect 12575 3674 12579 3726
rect 12523 3672 12579 3674
rect 12603 3726 12659 3728
rect 12603 3674 12655 3726
rect 12655 3674 12659 3726
rect 12603 3672 12659 3674
rect 12683 3726 12739 3728
rect 12683 3674 12735 3726
rect 12735 3674 12739 3726
rect 12683 3672 12739 3674
rect 12763 3726 12819 3728
rect 12763 3674 12815 3726
rect 12815 3674 12819 3726
rect 12763 3672 12819 3674
rect 12843 3726 12899 3728
rect 12843 3674 12895 3726
rect 12895 3674 12899 3726
rect 12843 3672 12899 3674
rect 12923 3726 12979 3728
rect 12923 3674 12975 3726
rect 12975 3674 12979 3726
rect 12923 3672 12979 3674
rect 13260 3670 13316 3672
rect 13260 3618 13262 3670
rect 13262 3618 13314 3670
rect 13314 3618 13316 3670
rect 13260 3616 13316 3618
rect 6556 3526 6612 3528
rect 6556 3474 6558 3526
rect 6558 3474 6610 3526
rect 6610 3474 6612 3526
rect 6556 3472 6612 3474
rect 7017 3501 7073 3503
rect 7017 3449 7019 3501
rect 7019 3449 7071 3501
rect 7071 3449 7073 3501
rect 7017 3447 7073 3449
rect 13265 3526 13321 3528
rect 13265 3474 13267 3526
rect 13267 3474 13319 3526
rect 13319 3474 13321 3526
rect 13265 3472 13321 3474
rect 6557 3374 6613 3376
rect 6557 3322 6559 3374
rect 6559 3322 6611 3374
rect 6611 3322 6613 3374
rect 6557 3320 6613 3322
rect 13266 3374 13322 3376
rect 13266 3322 13268 3374
rect 13268 3322 13320 3374
rect 13320 3322 13322 3374
rect 13266 3320 13322 3322
rect 7017 3309 7073 3311
rect 7017 3257 7019 3309
rect 7019 3257 7071 3309
rect 7071 3257 7073 3309
rect 7017 3255 7073 3257
rect 6557 3204 6613 3206
rect 6557 3152 6559 3204
rect 6559 3152 6611 3204
rect 6611 3152 6613 3204
rect 6557 3150 6613 3152
rect 13266 3204 13322 3206
rect 13266 3152 13268 3204
rect 13268 3152 13320 3204
rect 13320 3152 13322 3204
rect 13266 3150 13322 3152
rect 125 3127 181 3129
rect 125 3075 127 3127
rect 127 3075 179 3127
rect 179 3075 181 3127
rect 125 3073 181 3075
rect 256 3126 312 3128
rect 256 3074 258 3126
rect 258 3074 310 3126
rect 310 3074 312 3126
rect 256 3072 312 3074
rect 400 3127 456 3129
rect 400 3075 402 3127
rect 402 3075 454 3127
rect 454 3075 456 3127
rect 400 3073 456 3075
rect 6834 3127 6890 3129
rect 6834 3075 6836 3127
rect 6836 3075 6888 3127
rect 6888 3075 6890 3127
rect 6834 3073 6890 3075
rect 6965 3126 7021 3128
rect 6965 3074 6967 3126
rect 6967 3074 7019 3126
rect 7019 3074 7021 3126
rect 6965 3072 7021 3074
rect 7109 3127 7165 3129
rect 7109 3075 7111 3127
rect 7111 3075 7163 3127
rect 7163 3075 7165 3127
rect 7109 3073 7165 3075
rect 6556 3047 6612 3049
rect 6556 2995 6558 3047
rect 6558 2995 6610 3047
rect 6610 2995 6612 3047
rect 6556 2993 6612 2995
rect 13265 3047 13321 3049
rect 13265 2995 13267 3047
rect 13267 2995 13319 3047
rect 13319 2995 13321 3047
rect 13265 2993 13321 2995
rect 6474 2805 6530 2807
rect 6474 2753 6476 2805
rect 6476 2753 6528 2805
rect 6528 2753 6530 2805
rect 6474 2751 6530 2753
rect 13183 2805 13239 2807
rect 13183 2753 13185 2805
rect 13185 2753 13237 2805
rect 13237 2753 13239 2805
rect 13183 2751 13239 2753
rect 143 2581 199 2583
rect 143 2529 145 2581
rect 145 2529 197 2581
rect 197 2529 199 2581
rect 143 2527 199 2529
rect 263 2581 319 2583
rect 263 2529 265 2581
rect 265 2529 317 2581
rect 317 2529 319 2581
rect 263 2527 319 2529
rect 406 2581 462 2583
rect 406 2529 408 2581
rect 408 2529 460 2581
rect 460 2529 462 2581
rect 406 2527 462 2529
rect 6852 2581 6908 2583
rect 1224 2481 1288 2545
rect 1956 2484 2020 2548
rect 2184 2484 2248 2548
rect 3168 2484 3232 2548
rect 3396 2484 3460 2548
rect 4380 2484 4444 2548
rect 4608 2484 4672 2548
rect 5592 2484 5656 2548
rect 5820 2484 5884 2548
rect 6562 2544 6618 2546
rect 6562 2492 6564 2544
rect 6564 2492 6616 2544
rect 6616 2492 6618 2544
rect 6562 2490 6618 2492
rect 6852 2529 6854 2581
rect 6854 2529 6906 2581
rect 6906 2529 6908 2581
rect 6852 2527 6908 2529
rect 6972 2581 7028 2583
rect 6972 2529 6974 2581
rect 6974 2529 7026 2581
rect 7026 2529 7028 2581
rect 6972 2527 7028 2529
rect 7115 2581 7171 2583
rect 7115 2529 7117 2581
rect 7117 2529 7169 2581
rect 7169 2529 7171 2581
rect 7115 2527 7171 2529
rect 1580 2282 1644 2346
rect 2312 2282 2376 2346
rect 2530 2282 2594 2346
rect 3524 2282 3588 2346
rect 3742 2282 3806 2346
rect 4862 2282 4926 2346
rect 5080 2282 5144 2346
rect 5814 2282 5878 2346
rect 6562 2341 6618 2343
rect 6562 2289 6564 2341
rect 6564 2289 6616 2341
rect 6616 2289 6618 2341
rect 6562 2287 6618 2289
rect 7933 2481 7997 2545
rect 8665 2484 8729 2548
rect 8893 2484 8957 2548
rect 9877 2484 9941 2548
rect 10105 2484 10169 2548
rect 11089 2484 11153 2548
rect 11317 2484 11381 2548
rect 12301 2484 12365 2548
rect 12529 2484 12593 2548
rect 13271 2544 13327 2546
rect 13271 2492 13273 2544
rect 13273 2492 13325 2544
rect 13325 2492 13327 2544
rect 13271 2490 13327 2492
rect 8289 2282 8353 2346
rect 9021 2282 9085 2346
rect 9239 2282 9303 2346
rect 10233 2282 10297 2346
rect 10451 2282 10515 2346
rect 11571 2282 11635 2346
rect 11789 2282 11853 2346
rect 12523 2282 12587 2346
rect 13271 2341 13327 2343
rect 13271 2289 13273 2341
rect 13273 2289 13325 2341
rect 13325 2289 13327 2341
rect 13271 2287 13327 2289
rect 102 1700 169 1701
rect 102 1644 105 1700
rect 105 1644 165 1700
rect 165 1644 169 1700
rect 102 1643 169 1644
rect 728 1154 784 1156
rect 728 1102 730 1154
rect 730 1102 782 1154
rect 782 1102 784 1154
rect 728 1100 784 1102
rect 6471 2079 6527 2081
rect 6471 2027 6473 2079
rect 6473 2027 6525 2079
rect 6525 2027 6527 2079
rect 6471 2025 6527 2027
rect 1270 1157 1326 1159
rect 1270 1105 1272 1157
rect 1272 1105 1324 1157
rect 1324 1105 1326 1157
rect 1270 1103 1326 1105
rect 1350 1157 1406 1159
rect 1350 1105 1352 1157
rect 1352 1105 1404 1157
rect 1404 1105 1406 1157
rect 1350 1103 1406 1105
rect 1430 1157 1486 1159
rect 1430 1105 1432 1157
rect 1432 1105 1484 1157
rect 1484 1105 1486 1157
rect 1430 1103 1486 1105
rect 1510 1157 1566 1159
rect 1510 1105 1512 1157
rect 1512 1105 1564 1157
rect 1564 1105 1566 1157
rect 1510 1103 1566 1105
rect 2002 1157 2058 1159
rect 2002 1105 2004 1157
rect 2004 1105 2056 1157
rect 2056 1105 2058 1157
rect 2002 1103 2058 1105
rect 2082 1157 2138 1159
rect 2082 1105 2084 1157
rect 2084 1105 2136 1157
rect 2136 1105 2138 1157
rect 2082 1103 2138 1105
rect 2162 1157 2218 1159
rect 2162 1105 2164 1157
rect 2164 1105 2216 1157
rect 2216 1105 2218 1157
rect 2162 1103 2218 1105
rect 2242 1157 2298 1159
rect 2242 1105 2244 1157
rect 2244 1105 2296 1157
rect 2296 1105 2298 1157
rect 2242 1103 2298 1105
rect 2608 1157 2664 1159
rect 2608 1105 2610 1157
rect 2610 1105 2662 1157
rect 2662 1105 2664 1157
rect 2608 1103 2664 1105
rect 2688 1157 2744 1159
rect 2688 1105 2690 1157
rect 2690 1105 2742 1157
rect 2742 1105 2744 1157
rect 2688 1103 2744 1105
rect 2768 1157 2824 1159
rect 2768 1105 2770 1157
rect 2770 1105 2822 1157
rect 2822 1105 2824 1157
rect 2768 1103 2824 1105
rect 2848 1157 2904 1159
rect 2848 1105 2850 1157
rect 2850 1105 2902 1157
rect 2902 1105 2904 1157
rect 2848 1103 2904 1105
rect 3214 1157 3270 1159
rect 3214 1105 3216 1157
rect 3216 1105 3268 1157
rect 3268 1105 3270 1157
rect 3214 1103 3270 1105
rect 3294 1157 3350 1159
rect 3294 1105 3296 1157
rect 3296 1105 3348 1157
rect 3348 1105 3350 1157
rect 3294 1103 3350 1105
rect 3374 1157 3430 1159
rect 3374 1105 3376 1157
rect 3376 1105 3428 1157
rect 3428 1105 3430 1157
rect 3374 1103 3430 1105
rect 3454 1157 3510 1159
rect 3454 1105 3456 1157
rect 3456 1105 3508 1157
rect 3508 1105 3510 1157
rect 3454 1103 3510 1105
rect 3820 1157 3876 1159
rect 3820 1105 3822 1157
rect 3822 1105 3874 1157
rect 3874 1105 3876 1157
rect 3820 1103 3876 1105
rect 3900 1157 3956 1159
rect 3900 1105 3902 1157
rect 3902 1105 3954 1157
rect 3954 1105 3956 1157
rect 3900 1103 3956 1105
rect 3980 1157 4036 1159
rect 3980 1105 3982 1157
rect 3982 1105 4034 1157
rect 4034 1105 4036 1157
rect 3980 1103 4036 1105
rect 4060 1157 4116 1159
rect 4060 1105 4062 1157
rect 4062 1105 4114 1157
rect 4114 1105 4116 1157
rect 4060 1103 4116 1105
rect 4552 1157 4608 1159
rect 4552 1105 4554 1157
rect 4554 1105 4606 1157
rect 4606 1105 4608 1157
rect 4552 1103 4608 1105
rect 4632 1157 4688 1159
rect 4632 1105 4634 1157
rect 4634 1105 4686 1157
rect 4686 1105 4688 1157
rect 4632 1103 4688 1105
rect 4712 1157 4768 1159
rect 4712 1105 4714 1157
rect 4714 1105 4766 1157
rect 4766 1105 4768 1157
rect 4712 1103 4768 1105
rect 4792 1157 4848 1159
rect 4792 1105 4794 1157
rect 4794 1105 4846 1157
rect 4846 1105 4848 1157
rect 4792 1103 4848 1105
rect 5158 1157 5214 1159
rect 5158 1105 5160 1157
rect 5160 1105 5212 1157
rect 5212 1105 5214 1157
rect 5158 1103 5214 1105
rect 5238 1157 5294 1159
rect 5238 1105 5240 1157
rect 5240 1105 5292 1157
rect 5292 1105 5294 1157
rect 5238 1103 5294 1105
rect 5318 1157 5374 1159
rect 5318 1105 5320 1157
rect 5320 1105 5372 1157
rect 5372 1105 5374 1157
rect 5318 1103 5374 1105
rect 5398 1157 5454 1159
rect 5398 1105 5400 1157
rect 5400 1105 5452 1157
rect 5452 1105 5454 1157
rect 5398 1103 5454 1105
rect 5892 1157 5948 1159
rect 5892 1105 5894 1157
rect 5894 1105 5946 1157
rect 5946 1105 5948 1157
rect 5892 1103 5948 1105
rect 5972 1157 6028 1159
rect 5972 1105 5974 1157
rect 5974 1105 6026 1157
rect 6026 1105 6028 1157
rect 5972 1103 6028 1105
rect 6052 1157 6108 1159
rect 6052 1105 6054 1157
rect 6054 1105 6106 1157
rect 6106 1105 6108 1157
rect 6052 1103 6108 1105
rect 6132 1157 6188 1159
rect 6132 1105 6134 1157
rect 6134 1105 6186 1157
rect 6186 1105 6188 1157
rect 6132 1103 6188 1105
rect 7437 1154 7493 1156
rect 7437 1102 7439 1154
rect 7439 1102 7491 1154
rect 7491 1102 7493 1154
rect 7437 1100 7493 1102
rect 13180 2079 13236 2081
rect 13180 2027 13182 2079
rect 13182 2027 13234 2079
rect 13234 2027 13236 2079
rect 13180 2025 13236 2027
rect 7979 1157 8035 1159
rect 7979 1105 7981 1157
rect 7981 1105 8033 1157
rect 8033 1105 8035 1157
rect 7979 1103 8035 1105
rect 8059 1157 8115 1159
rect 8059 1105 8061 1157
rect 8061 1105 8113 1157
rect 8113 1105 8115 1157
rect 8059 1103 8115 1105
rect 8139 1157 8195 1159
rect 8139 1105 8141 1157
rect 8141 1105 8193 1157
rect 8193 1105 8195 1157
rect 8139 1103 8195 1105
rect 8219 1157 8275 1159
rect 8219 1105 8221 1157
rect 8221 1105 8273 1157
rect 8273 1105 8275 1157
rect 8219 1103 8275 1105
rect 8711 1157 8767 1159
rect 8711 1105 8713 1157
rect 8713 1105 8765 1157
rect 8765 1105 8767 1157
rect 8711 1103 8767 1105
rect 8791 1157 8847 1159
rect 8791 1105 8793 1157
rect 8793 1105 8845 1157
rect 8845 1105 8847 1157
rect 8791 1103 8847 1105
rect 8871 1157 8927 1159
rect 8871 1105 8873 1157
rect 8873 1105 8925 1157
rect 8925 1105 8927 1157
rect 8871 1103 8927 1105
rect 8951 1157 9007 1159
rect 8951 1105 8953 1157
rect 8953 1105 9005 1157
rect 9005 1105 9007 1157
rect 8951 1103 9007 1105
rect 9317 1157 9373 1159
rect 9317 1105 9319 1157
rect 9319 1105 9371 1157
rect 9371 1105 9373 1157
rect 9317 1103 9373 1105
rect 9397 1157 9453 1159
rect 9397 1105 9399 1157
rect 9399 1105 9451 1157
rect 9451 1105 9453 1157
rect 9397 1103 9453 1105
rect 9477 1157 9533 1159
rect 9477 1105 9479 1157
rect 9479 1105 9531 1157
rect 9531 1105 9533 1157
rect 9477 1103 9533 1105
rect 9557 1157 9613 1159
rect 9557 1105 9559 1157
rect 9559 1105 9611 1157
rect 9611 1105 9613 1157
rect 9557 1103 9613 1105
rect 9923 1157 9979 1159
rect 9923 1105 9925 1157
rect 9925 1105 9977 1157
rect 9977 1105 9979 1157
rect 9923 1103 9979 1105
rect 10003 1157 10059 1159
rect 10003 1105 10005 1157
rect 10005 1105 10057 1157
rect 10057 1105 10059 1157
rect 10003 1103 10059 1105
rect 10083 1157 10139 1159
rect 10083 1105 10085 1157
rect 10085 1105 10137 1157
rect 10137 1105 10139 1157
rect 10083 1103 10139 1105
rect 10163 1157 10219 1159
rect 10163 1105 10165 1157
rect 10165 1105 10217 1157
rect 10217 1105 10219 1157
rect 10163 1103 10219 1105
rect 10529 1157 10585 1159
rect 10529 1105 10531 1157
rect 10531 1105 10583 1157
rect 10583 1105 10585 1157
rect 10529 1103 10585 1105
rect 10609 1157 10665 1159
rect 10609 1105 10611 1157
rect 10611 1105 10663 1157
rect 10663 1105 10665 1157
rect 10609 1103 10665 1105
rect 10689 1157 10745 1159
rect 10689 1105 10691 1157
rect 10691 1105 10743 1157
rect 10743 1105 10745 1157
rect 10689 1103 10745 1105
rect 10769 1157 10825 1159
rect 10769 1105 10771 1157
rect 10771 1105 10823 1157
rect 10823 1105 10825 1157
rect 10769 1103 10825 1105
rect 11261 1157 11317 1159
rect 11261 1105 11263 1157
rect 11263 1105 11315 1157
rect 11315 1105 11317 1157
rect 11261 1103 11317 1105
rect 11341 1157 11397 1159
rect 11341 1105 11343 1157
rect 11343 1105 11395 1157
rect 11395 1105 11397 1157
rect 11341 1103 11397 1105
rect 11421 1157 11477 1159
rect 11421 1105 11423 1157
rect 11423 1105 11475 1157
rect 11475 1105 11477 1157
rect 11421 1103 11477 1105
rect 11501 1157 11557 1159
rect 11501 1105 11503 1157
rect 11503 1105 11555 1157
rect 11555 1105 11557 1157
rect 11501 1103 11557 1105
rect 11867 1157 11923 1159
rect 11867 1105 11869 1157
rect 11869 1105 11921 1157
rect 11921 1105 11923 1157
rect 11867 1103 11923 1105
rect 11947 1157 12003 1159
rect 11947 1105 11949 1157
rect 11949 1105 12001 1157
rect 12001 1105 12003 1157
rect 11947 1103 12003 1105
rect 12027 1157 12083 1159
rect 12027 1105 12029 1157
rect 12029 1105 12081 1157
rect 12081 1105 12083 1157
rect 12027 1103 12083 1105
rect 12107 1157 12163 1159
rect 12107 1105 12109 1157
rect 12109 1105 12161 1157
rect 12161 1105 12163 1157
rect 12107 1103 12163 1105
rect 12601 1157 12657 1159
rect 12601 1105 12603 1157
rect 12603 1105 12655 1157
rect 12655 1105 12657 1157
rect 12601 1103 12657 1105
rect 12681 1157 12737 1159
rect 12681 1105 12683 1157
rect 12683 1105 12735 1157
rect 12735 1105 12737 1157
rect 12681 1103 12737 1105
rect 12761 1157 12817 1159
rect 12761 1105 12763 1157
rect 12763 1105 12815 1157
rect 12815 1105 12817 1157
rect 12761 1103 12817 1105
rect 12841 1157 12897 1159
rect 12841 1105 12843 1157
rect 12843 1105 12895 1157
rect 12895 1105 12897 1157
rect 12841 1103 12897 1105
rect 567 216 623 218
rect 567 164 569 216
rect 569 164 621 216
rect 621 164 623 216
rect 567 162 623 164
rect 647 216 703 218
rect 647 164 649 216
rect 649 164 701 216
rect 701 164 703 216
rect 647 162 703 164
rect 727 216 783 218
rect 727 164 729 216
rect 729 164 781 216
rect 781 164 783 216
rect 727 162 783 164
rect 807 216 863 218
rect 807 164 809 216
rect 809 164 861 216
rect 861 164 863 216
rect 807 162 863 164
rect 1301 216 1357 218
rect 1301 164 1303 216
rect 1303 164 1355 216
rect 1355 164 1357 216
rect 1301 162 1357 164
rect 1381 216 1437 218
rect 1381 164 1383 216
rect 1383 164 1435 216
rect 1435 164 1437 216
rect 1381 162 1437 164
rect 1461 216 1517 218
rect 1461 164 1463 216
rect 1463 164 1515 216
rect 1515 164 1517 216
rect 1461 162 1517 164
rect 1541 216 1597 218
rect 1541 164 1543 216
rect 1543 164 1595 216
rect 1595 164 1597 216
rect 1541 162 1597 164
rect 1907 216 1963 218
rect 1907 164 1909 216
rect 1909 164 1961 216
rect 1961 164 1963 216
rect 1907 162 1963 164
rect 1987 216 2043 218
rect 1987 164 1989 216
rect 1989 164 2041 216
rect 2041 164 2043 216
rect 1987 162 2043 164
rect 2067 216 2123 218
rect 2067 164 2069 216
rect 2069 164 2121 216
rect 2121 164 2123 216
rect 2067 162 2123 164
rect 2147 216 2203 218
rect 2147 164 2149 216
rect 2149 164 2201 216
rect 2201 164 2203 216
rect 2147 162 2203 164
rect 2639 216 2695 218
rect 2639 164 2641 216
rect 2641 164 2693 216
rect 2693 164 2695 216
rect 2639 162 2695 164
rect 2719 216 2775 218
rect 2719 164 2721 216
rect 2721 164 2773 216
rect 2773 164 2775 216
rect 2719 162 2775 164
rect 2799 216 2855 218
rect 2799 164 2801 216
rect 2801 164 2853 216
rect 2853 164 2855 216
rect 2799 162 2855 164
rect 2879 216 2935 218
rect 2879 164 2881 216
rect 2881 164 2933 216
rect 2933 164 2935 216
rect 2879 162 2935 164
rect 3245 216 3301 218
rect 3245 164 3247 216
rect 3247 164 3299 216
rect 3299 164 3301 216
rect 3245 162 3301 164
rect 3325 216 3381 218
rect 3325 164 3327 216
rect 3327 164 3379 216
rect 3379 164 3381 216
rect 3325 162 3381 164
rect 3405 216 3461 218
rect 3405 164 3407 216
rect 3407 164 3459 216
rect 3459 164 3461 216
rect 3405 162 3461 164
rect 3485 216 3541 218
rect 3485 164 3487 216
rect 3487 164 3539 216
rect 3539 164 3541 216
rect 3485 162 3541 164
rect 3851 216 3907 218
rect 3851 164 3853 216
rect 3853 164 3905 216
rect 3905 164 3907 216
rect 3851 162 3907 164
rect 3931 216 3987 218
rect 3931 164 3933 216
rect 3933 164 3985 216
rect 3985 164 3987 216
rect 3931 162 3987 164
rect 4011 216 4067 218
rect 4011 164 4013 216
rect 4013 164 4065 216
rect 4065 164 4067 216
rect 4011 162 4067 164
rect 4091 216 4147 218
rect 4091 164 4093 216
rect 4093 164 4145 216
rect 4145 164 4147 216
rect 4091 162 4147 164
rect 4457 216 4513 218
rect 4457 164 4459 216
rect 4459 164 4511 216
rect 4511 164 4513 216
rect 4457 162 4513 164
rect 4537 216 4593 218
rect 4537 164 4539 216
rect 4539 164 4591 216
rect 4591 164 4593 216
rect 4537 162 4593 164
rect 4617 216 4673 218
rect 4617 164 4619 216
rect 4619 164 4671 216
rect 4671 164 4673 216
rect 4617 162 4673 164
rect 4697 216 4753 218
rect 4697 164 4699 216
rect 4699 164 4751 216
rect 4751 164 4753 216
rect 4697 162 4753 164
rect 5189 216 5245 218
rect 5189 164 5191 216
rect 5191 164 5243 216
rect 5243 164 5245 216
rect 5189 162 5245 164
rect 5269 216 5325 218
rect 5269 164 5271 216
rect 5271 164 5323 216
rect 5323 164 5325 216
rect 5269 162 5325 164
rect 5349 216 5405 218
rect 5349 164 5351 216
rect 5351 164 5403 216
rect 5403 164 5405 216
rect 5349 162 5405 164
rect 5429 216 5485 218
rect 5429 164 5431 216
rect 5431 164 5483 216
rect 5483 164 5485 216
rect 5429 162 5485 164
rect 228 -706 284 -704
rect 228 -758 230 -706
rect 230 -758 282 -706
rect 282 -758 284 -706
rect 228 -760 284 -758
rect 5971 219 6027 221
rect 5971 167 5973 219
rect 5973 167 6025 219
rect 6025 167 6027 219
rect 5971 165 6027 167
rect 7276 216 7332 218
rect 7276 164 7278 216
rect 7278 164 7330 216
rect 7330 164 7332 216
rect 7276 162 7332 164
rect 7356 216 7412 218
rect 7356 164 7358 216
rect 7358 164 7410 216
rect 7410 164 7412 216
rect 7356 162 7412 164
rect 7436 216 7492 218
rect 7436 164 7438 216
rect 7438 164 7490 216
rect 7490 164 7492 216
rect 7436 162 7492 164
rect 7516 216 7572 218
rect 7516 164 7518 216
rect 7518 164 7570 216
rect 7570 164 7572 216
rect 7516 162 7572 164
rect 8010 216 8066 218
rect 8010 164 8012 216
rect 8012 164 8064 216
rect 8064 164 8066 216
rect 8010 162 8066 164
rect 8090 216 8146 218
rect 8090 164 8092 216
rect 8092 164 8144 216
rect 8144 164 8146 216
rect 8090 162 8146 164
rect 8170 216 8226 218
rect 8170 164 8172 216
rect 8172 164 8224 216
rect 8224 164 8226 216
rect 8170 162 8226 164
rect 8250 216 8306 218
rect 8250 164 8252 216
rect 8252 164 8304 216
rect 8304 164 8306 216
rect 8250 162 8306 164
rect 8616 216 8672 218
rect 8616 164 8618 216
rect 8618 164 8670 216
rect 8670 164 8672 216
rect 8616 162 8672 164
rect 8696 216 8752 218
rect 8696 164 8698 216
rect 8698 164 8750 216
rect 8750 164 8752 216
rect 8696 162 8752 164
rect 8776 216 8832 218
rect 8776 164 8778 216
rect 8778 164 8830 216
rect 8830 164 8832 216
rect 8776 162 8832 164
rect 8856 216 8912 218
rect 8856 164 8858 216
rect 8858 164 8910 216
rect 8910 164 8912 216
rect 8856 162 8912 164
rect 9348 216 9404 218
rect 9348 164 9350 216
rect 9350 164 9402 216
rect 9402 164 9404 216
rect 9348 162 9404 164
rect 9428 216 9484 218
rect 9428 164 9430 216
rect 9430 164 9482 216
rect 9482 164 9484 216
rect 9428 162 9484 164
rect 9508 216 9564 218
rect 9508 164 9510 216
rect 9510 164 9562 216
rect 9562 164 9564 216
rect 9508 162 9564 164
rect 9588 216 9644 218
rect 9588 164 9590 216
rect 9590 164 9642 216
rect 9642 164 9644 216
rect 9588 162 9644 164
rect 9954 216 10010 218
rect 9954 164 9956 216
rect 9956 164 10008 216
rect 10008 164 10010 216
rect 9954 162 10010 164
rect 10034 216 10090 218
rect 10034 164 10036 216
rect 10036 164 10088 216
rect 10088 164 10090 216
rect 10034 162 10090 164
rect 10114 216 10170 218
rect 10114 164 10116 216
rect 10116 164 10168 216
rect 10168 164 10170 216
rect 10114 162 10170 164
rect 10194 216 10250 218
rect 10194 164 10196 216
rect 10196 164 10248 216
rect 10248 164 10250 216
rect 10194 162 10250 164
rect 10560 216 10616 218
rect 10560 164 10562 216
rect 10562 164 10614 216
rect 10614 164 10616 216
rect 10560 162 10616 164
rect 10640 216 10696 218
rect 10640 164 10642 216
rect 10642 164 10694 216
rect 10694 164 10696 216
rect 10640 162 10696 164
rect 10720 216 10776 218
rect 10720 164 10722 216
rect 10722 164 10774 216
rect 10774 164 10776 216
rect 10720 162 10776 164
rect 10800 216 10856 218
rect 10800 164 10802 216
rect 10802 164 10854 216
rect 10854 164 10856 216
rect 10800 162 10856 164
rect 11166 216 11222 218
rect 11166 164 11168 216
rect 11168 164 11220 216
rect 11220 164 11222 216
rect 11166 162 11222 164
rect 11246 216 11302 218
rect 11246 164 11248 216
rect 11248 164 11300 216
rect 11300 164 11302 216
rect 11246 162 11302 164
rect 11326 216 11382 218
rect 11326 164 11328 216
rect 11328 164 11380 216
rect 11380 164 11382 216
rect 11326 162 11382 164
rect 11406 216 11462 218
rect 11406 164 11408 216
rect 11408 164 11460 216
rect 11460 164 11462 216
rect 11406 162 11462 164
rect 11898 216 11954 218
rect 11898 164 11900 216
rect 11900 164 11952 216
rect 11952 164 11954 216
rect 11898 162 11954 164
rect 11978 216 12034 218
rect 11978 164 11980 216
rect 11980 164 12032 216
rect 12032 164 12034 216
rect 11978 162 12034 164
rect 12058 216 12114 218
rect 12058 164 12060 216
rect 12060 164 12112 216
rect 12112 164 12114 216
rect 12058 162 12114 164
rect 12138 216 12194 218
rect 12138 164 12140 216
rect 12140 164 12192 216
rect 12192 164 12194 216
rect 12138 162 12194 164
rect 6937 -706 6993 -704
rect 6937 -758 6939 -706
rect 6939 -758 6991 -706
rect 6991 -758 6993 -706
rect 6937 -760 6993 -758
rect 12680 219 12736 221
rect 12680 167 12682 219
rect 12682 167 12734 219
rect 12734 167 12736 219
rect 12680 165 12736 167
rect 137 -968 193 -966
rect 137 -1020 139 -968
rect 139 -1020 191 -968
rect 191 -1020 193 -968
rect 137 -1022 193 -1020
rect 877 -1025 941 -961
rect 1611 -1025 1675 -961
rect 1829 -1025 1893 -961
rect 2949 -1025 3013 -961
rect 3167 -1025 3231 -961
rect 4161 -1025 4225 -961
rect 4379 -1025 4443 -961
rect 5111 -1025 5175 -961
rect 137 -1171 193 -1169
rect 137 -1223 139 -1171
rect 139 -1223 191 -1171
rect 191 -1223 193 -1171
rect 137 -1225 193 -1223
rect 871 -1227 935 -1163
rect 1099 -1227 1163 -1163
rect 2083 -1227 2147 -1163
rect 2311 -1227 2375 -1163
rect 3295 -1227 3359 -1163
rect 3523 -1227 3587 -1163
rect 4507 -1227 4571 -1163
rect 4735 -1227 4799 -1163
rect 5467 -1224 5531 -1160
rect 6846 -968 6902 -966
rect 6846 -1020 6848 -968
rect 6848 -1020 6900 -968
rect 6900 -1020 6902 -968
rect 6846 -1022 6902 -1020
rect 7586 -1025 7650 -961
rect 8320 -1025 8384 -961
rect 8538 -1025 8602 -961
rect 9658 -1025 9722 -961
rect 9876 -1025 9940 -961
rect 10870 -1025 10934 -961
rect 11088 -1025 11152 -961
rect 11820 -1025 11884 -961
rect 6293 -1208 6349 -1206
rect 6293 -1260 6295 -1208
rect 6295 -1260 6347 -1208
rect 6347 -1260 6349 -1208
rect 6293 -1262 6349 -1260
rect 6436 -1208 6492 -1206
rect 6436 -1260 6438 -1208
rect 6438 -1260 6490 -1208
rect 6490 -1260 6492 -1208
rect 6436 -1262 6492 -1260
rect 6556 -1208 6612 -1206
rect 6556 -1260 6558 -1208
rect 6558 -1260 6610 -1208
rect 6610 -1260 6612 -1208
rect 6846 -1171 6902 -1169
rect 6846 -1223 6848 -1171
rect 6848 -1223 6900 -1171
rect 6900 -1223 6902 -1171
rect 6846 -1225 6902 -1223
rect 7580 -1227 7644 -1163
rect 7808 -1227 7872 -1163
rect 8792 -1227 8856 -1163
rect 9020 -1227 9084 -1163
rect 10004 -1227 10068 -1163
rect 10232 -1227 10296 -1163
rect 11216 -1227 11280 -1163
rect 11444 -1227 11508 -1163
rect 12176 -1224 12240 -1160
rect 6556 -1262 6612 -1260
rect 13002 -1208 13058 -1206
rect 13002 -1260 13004 -1208
rect 13004 -1260 13056 -1208
rect 13056 -1260 13058 -1208
rect 13002 -1262 13058 -1260
rect 13145 -1208 13201 -1206
rect 13145 -1260 13147 -1208
rect 13147 -1260 13199 -1208
rect 13199 -1260 13201 -1208
rect 13145 -1262 13201 -1260
rect 13265 -1208 13321 -1206
rect 13265 -1260 13267 -1208
rect 13267 -1260 13319 -1208
rect 13319 -1260 13321 -1208
rect 13265 -1262 13321 -1260
rect 225 -1432 281 -1430
rect 225 -1484 227 -1432
rect 227 -1484 279 -1432
rect 279 -1484 281 -1432
rect 225 -1486 281 -1484
rect 6934 -1432 6990 -1430
rect 6934 -1484 6936 -1432
rect 6936 -1484 6988 -1432
rect 6988 -1484 6990 -1432
rect 6934 -1486 6990 -1484
rect 143 -1674 199 -1672
rect 143 -1726 145 -1674
rect 145 -1726 197 -1674
rect 197 -1726 199 -1674
rect 143 -1728 199 -1726
rect 6852 -1674 6908 -1672
rect 6852 -1726 6854 -1674
rect 6854 -1726 6906 -1674
rect 6906 -1726 6908 -1674
rect 6852 -1728 6908 -1726
rect 6299 -1754 6355 -1752
rect 6299 -1806 6301 -1754
rect 6301 -1806 6353 -1754
rect 6353 -1806 6355 -1754
rect 6299 -1808 6355 -1806
rect 6443 -1753 6499 -1751
rect 6443 -1805 6445 -1753
rect 6445 -1805 6497 -1753
rect 6497 -1805 6499 -1753
rect 6443 -1807 6499 -1805
rect 6574 -1754 6630 -1752
rect 6574 -1806 6576 -1754
rect 6576 -1806 6628 -1754
rect 6628 -1806 6630 -1754
rect 6574 -1808 6630 -1806
rect 13008 -1754 13064 -1752
rect 13008 -1806 13010 -1754
rect 13010 -1806 13062 -1754
rect 13062 -1806 13064 -1754
rect 13008 -1808 13064 -1806
rect 13152 -1753 13208 -1751
rect 13152 -1805 13154 -1753
rect 13154 -1805 13206 -1753
rect 13206 -1805 13208 -1753
rect 13152 -1807 13208 -1805
rect 13283 -1754 13339 -1752
rect 13283 -1806 13285 -1754
rect 13285 -1806 13337 -1754
rect 13337 -1806 13339 -1754
rect 13283 -1808 13339 -1806
rect 142 -1831 198 -1829
rect 142 -1883 144 -1831
rect 144 -1883 196 -1831
rect 196 -1883 198 -1831
rect 142 -1885 198 -1883
rect 6851 -1831 6907 -1829
rect 6851 -1883 6853 -1831
rect 6853 -1883 6905 -1831
rect 6905 -1883 6907 -1831
rect 6851 -1885 6907 -1883
rect 6429 -1903 6485 -1901
rect 6429 -1955 6431 -1903
rect 6431 -1955 6483 -1903
rect 6483 -1955 6485 -1903
rect 6429 -1957 6485 -1955
rect 142 -2001 198 -1999
rect 142 -2053 144 -2001
rect 144 -2053 196 -2001
rect 196 -2053 198 -2001
rect 142 -2055 198 -2053
rect 6851 -2001 6907 -1999
rect 6851 -2053 6853 -2001
rect 6853 -2053 6905 -2001
rect 6905 -2053 6907 -2001
rect 6851 -2055 6907 -2053
rect 143 -2153 199 -2151
rect 143 -2205 145 -2153
rect 145 -2205 197 -2153
rect 197 -2205 199 -2153
rect 143 -2207 199 -2205
rect 6429 -2099 6485 -2097
rect 6429 -2151 6431 -2099
rect 6431 -2151 6483 -2099
rect 6483 -2151 6485 -2099
rect 6429 -2153 6485 -2151
rect 6852 -2153 6908 -2151
rect 6852 -2205 6854 -2153
rect 6854 -2205 6906 -2153
rect 6906 -2205 6908 -2153
rect 6852 -2207 6908 -2205
rect 148 -2297 204 -2295
rect 148 -2349 150 -2297
rect 150 -2349 202 -2297
rect 202 -2349 204 -2297
rect 148 -2351 204 -2349
rect 6429 -2274 6485 -2272
rect 6429 -2326 6431 -2274
rect 6431 -2326 6483 -2274
rect 6483 -2326 6485 -2274
rect 6429 -2328 6485 -2326
rect 485 -2353 541 -2351
rect 485 -2405 489 -2353
rect 489 -2405 541 -2353
rect 485 -2407 541 -2405
rect 565 -2353 621 -2351
rect 565 -2405 569 -2353
rect 569 -2405 621 -2353
rect 565 -2407 621 -2405
rect 645 -2353 701 -2351
rect 645 -2405 649 -2353
rect 649 -2405 701 -2353
rect 645 -2407 701 -2405
rect 725 -2353 781 -2351
rect 725 -2405 729 -2353
rect 729 -2405 781 -2353
rect 725 -2407 781 -2405
rect 805 -2353 861 -2351
rect 805 -2405 809 -2353
rect 809 -2405 861 -2353
rect 805 -2407 861 -2405
rect 885 -2353 941 -2351
rect 885 -2405 889 -2353
rect 889 -2405 941 -2353
rect 885 -2407 941 -2405
rect 1093 -2353 1149 -2351
rect 1093 -2405 1145 -2353
rect 1145 -2405 1149 -2353
rect 1093 -2407 1149 -2405
rect 1173 -2353 1229 -2351
rect 1173 -2405 1225 -2353
rect 1225 -2405 1229 -2353
rect 1173 -2407 1229 -2405
rect 1253 -2353 1309 -2351
rect 1253 -2405 1305 -2353
rect 1305 -2405 1309 -2353
rect 1253 -2407 1309 -2405
rect 1333 -2353 1389 -2351
rect 1333 -2405 1385 -2353
rect 1385 -2405 1389 -2353
rect 1333 -2407 1389 -2405
rect 1413 -2353 1469 -2351
rect 1413 -2405 1465 -2353
rect 1465 -2405 1469 -2353
rect 1413 -2407 1469 -2405
rect 1493 -2353 1549 -2351
rect 1493 -2405 1545 -2353
rect 1545 -2405 1549 -2353
rect 1493 -2407 1549 -2405
rect 1697 -2353 1753 -2351
rect 1697 -2405 1701 -2353
rect 1701 -2405 1753 -2353
rect 1697 -2407 1753 -2405
rect 1777 -2353 1833 -2351
rect 1777 -2405 1781 -2353
rect 1781 -2405 1833 -2353
rect 1777 -2407 1833 -2405
rect 1857 -2353 1913 -2351
rect 1857 -2405 1861 -2353
rect 1861 -2405 1913 -2353
rect 1857 -2407 1913 -2405
rect 1937 -2353 1993 -2351
rect 1937 -2405 1941 -2353
rect 1941 -2405 1993 -2353
rect 1937 -2407 1993 -2405
rect 2017 -2353 2073 -2351
rect 2017 -2405 2021 -2353
rect 2021 -2405 2073 -2353
rect 2017 -2407 2073 -2405
rect 2097 -2353 2153 -2351
rect 2097 -2405 2101 -2353
rect 2101 -2405 2153 -2353
rect 2097 -2407 2153 -2405
rect 2305 -2353 2361 -2351
rect 2305 -2405 2357 -2353
rect 2357 -2405 2361 -2353
rect 2305 -2407 2361 -2405
rect 2385 -2353 2441 -2351
rect 2385 -2405 2437 -2353
rect 2437 -2405 2441 -2353
rect 2385 -2407 2441 -2405
rect 2465 -2353 2521 -2351
rect 2465 -2405 2517 -2353
rect 2517 -2405 2521 -2353
rect 2465 -2407 2521 -2405
rect 2545 -2353 2601 -2351
rect 2545 -2405 2597 -2353
rect 2597 -2405 2601 -2353
rect 2545 -2407 2601 -2405
rect 2625 -2353 2681 -2351
rect 2625 -2405 2677 -2353
rect 2677 -2405 2681 -2353
rect 2625 -2407 2681 -2405
rect 2705 -2353 2761 -2351
rect 2705 -2405 2757 -2353
rect 2757 -2405 2761 -2353
rect 2705 -2407 2761 -2405
rect 2909 -2353 2965 -2351
rect 2909 -2405 2913 -2353
rect 2913 -2405 2965 -2353
rect 2909 -2407 2965 -2405
rect 2989 -2353 3045 -2351
rect 2989 -2405 2993 -2353
rect 2993 -2405 3045 -2353
rect 2989 -2407 3045 -2405
rect 3069 -2353 3125 -2351
rect 3069 -2405 3073 -2353
rect 3073 -2405 3125 -2353
rect 3069 -2407 3125 -2405
rect 3149 -2353 3205 -2351
rect 3149 -2405 3153 -2353
rect 3153 -2405 3205 -2353
rect 3149 -2407 3205 -2405
rect 3229 -2353 3285 -2351
rect 3229 -2405 3233 -2353
rect 3233 -2405 3285 -2353
rect 3229 -2407 3285 -2405
rect 3309 -2353 3365 -2351
rect 3309 -2405 3313 -2353
rect 3313 -2405 3365 -2353
rect 3309 -2407 3365 -2405
rect 3517 -2353 3573 -2351
rect 3517 -2405 3569 -2353
rect 3569 -2405 3573 -2353
rect 3517 -2407 3573 -2405
rect 3597 -2353 3653 -2351
rect 3597 -2405 3649 -2353
rect 3649 -2405 3653 -2353
rect 3597 -2407 3653 -2405
rect 3677 -2353 3733 -2351
rect 3677 -2405 3729 -2353
rect 3729 -2405 3733 -2353
rect 3677 -2407 3733 -2405
rect 3757 -2353 3813 -2351
rect 3757 -2405 3809 -2353
rect 3809 -2405 3813 -2353
rect 3757 -2407 3813 -2405
rect 3837 -2353 3893 -2351
rect 3837 -2405 3889 -2353
rect 3889 -2405 3893 -2353
rect 3837 -2407 3893 -2405
rect 3917 -2353 3973 -2351
rect 3917 -2405 3969 -2353
rect 3969 -2405 3973 -2353
rect 3917 -2407 3973 -2405
rect 4121 -2353 4177 -2351
rect 4121 -2405 4125 -2353
rect 4125 -2405 4177 -2353
rect 4121 -2407 4177 -2405
rect 4201 -2353 4257 -2351
rect 4201 -2405 4205 -2353
rect 4205 -2405 4257 -2353
rect 4201 -2407 4257 -2405
rect 4281 -2353 4337 -2351
rect 4281 -2405 4285 -2353
rect 4285 -2405 4337 -2353
rect 4281 -2407 4337 -2405
rect 4361 -2353 4417 -2351
rect 4361 -2405 4365 -2353
rect 4365 -2405 4417 -2353
rect 4361 -2407 4417 -2405
rect 4441 -2353 4497 -2351
rect 4441 -2405 4445 -2353
rect 4445 -2405 4497 -2353
rect 4441 -2407 4497 -2405
rect 4521 -2353 4577 -2351
rect 4521 -2405 4525 -2353
rect 4525 -2405 4577 -2353
rect 4521 -2407 4577 -2405
rect 4729 -2353 4785 -2351
rect 4729 -2405 4781 -2353
rect 4781 -2405 4785 -2353
rect 4729 -2407 4785 -2405
rect 4809 -2353 4865 -2351
rect 4809 -2405 4861 -2353
rect 4861 -2405 4865 -2353
rect 4809 -2407 4865 -2405
rect 4889 -2353 4945 -2351
rect 4889 -2405 4941 -2353
rect 4941 -2405 4945 -2353
rect 4889 -2407 4945 -2405
rect 4969 -2353 5025 -2351
rect 4969 -2405 5021 -2353
rect 5021 -2405 5025 -2353
rect 4969 -2407 5025 -2405
rect 5049 -2353 5105 -2351
rect 5049 -2405 5101 -2353
rect 5101 -2405 5105 -2353
rect 5049 -2407 5105 -2405
rect 5129 -2353 5185 -2351
rect 5129 -2405 5181 -2353
rect 5181 -2405 5185 -2353
rect 5129 -2407 5185 -2405
rect 5461 -2350 5517 -2348
rect 5461 -2402 5513 -2350
rect 5513 -2402 5517 -2350
rect 5461 -2404 5517 -2402
rect 5541 -2350 5597 -2348
rect 5541 -2402 5593 -2350
rect 5593 -2402 5597 -2350
rect 5541 -2404 5597 -2402
rect 5621 -2350 5677 -2348
rect 5621 -2402 5673 -2350
rect 5673 -2402 5677 -2350
rect 5621 -2404 5677 -2402
rect 5701 -2350 5757 -2348
rect 5701 -2402 5753 -2350
rect 5753 -2402 5757 -2350
rect 5701 -2404 5757 -2402
rect 5781 -2350 5837 -2348
rect 5781 -2402 5833 -2350
rect 5833 -2402 5837 -2350
rect 5781 -2404 5837 -2402
rect 5861 -2350 5917 -2348
rect 5861 -2402 5913 -2350
rect 5913 -2402 5917 -2350
rect 6857 -2297 6913 -2295
rect 6857 -2349 6859 -2297
rect 6859 -2349 6911 -2297
rect 6911 -2349 6913 -2297
rect 6857 -2351 6913 -2349
rect 5861 -2404 5917 -2402
rect 5957 -2359 6013 -2357
rect 5957 -2411 5959 -2359
rect 5959 -2411 6011 -2359
rect 6011 -2411 6013 -2359
rect 5957 -2413 6013 -2411
rect 7194 -2353 7250 -2351
rect 7194 -2405 7198 -2353
rect 7198 -2405 7250 -2353
rect 7194 -2407 7250 -2405
rect 7274 -2353 7330 -2351
rect 7274 -2405 7278 -2353
rect 7278 -2405 7330 -2353
rect 7274 -2407 7330 -2405
rect 7354 -2353 7410 -2351
rect 7354 -2405 7358 -2353
rect 7358 -2405 7410 -2353
rect 7354 -2407 7410 -2405
rect 7434 -2353 7490 -2351
rect 7434 -2405 7438 -2353
rect 7438 -2405 7490 -2353
rect 7434 -2407 7490 -2405
rect 7514 -2353 7570 -2351
rect 7514 -2405 7518 -2353
rect 7518 -2405 7570 -2353
rect 7514 -2407 7570 -2405
rect 7594 -2353 7650 -2351
rect 7594 -2405 7598 -2353
rect 7598 -2405 7650 -2353
rect 7594 -2407 7650 -2405
rect 7802 -2353 7858 -2351
rect 7802 -2405 7854 -2353
rect 7854 -2405 7858 -2353
rect 7802 -2407 7858 -2405
rect 7882 -2353 7938 -2351
rect 7882 -2405 7934 -2353
rect 7934 -2405 7938 -2353
rect 7882 -2407 7938 -2405
rect 7962 -2353 8018 -2351
rect 7962 -2405 8014 -2353
rect 8014 -2405 8018 -2353
rect 7962 -2407 8018 -2405
rect 8042 -2353 8098 -2351
rect 8042 -2405 8094 -2353
rect 8094 -2405 8098 -2353
rect 8042 -2407 8098 -2405
rect 8122 -2353 8178 -2351
rect 8122 -2405 8174 -2353
rect 8174 -2405 8178 -2353
rect 8122 -2407 8178 -2405
rect 8202 -2353 8258 -2351
rect 8202 -2405 8254 -2353
rect 8254 -2405 8258 -2353
rect 8202 -2407 8258 -2405
rect 8406 -2353 8462 -2351
rect 8406 -2405 8410 -2353
rect 8410 -2405 8462 -2353
rect 8406 -2407 8462 -2405
rect 8486 -2353 8542 -2351
rect 8486 -2405 8490 -2353
rect 8490 -2405 8542 -2353
rect 8486 -2407 8542 -2405
rect 8566 -2353 8622 -2351
rect 8566 -2405 8570 -2353
rect 8570 -2405 8622 -2353
rect 8566 -2407 8622 -2405
rect 8646 -2353 8702 -2351
rect 8646 -2405 8650 -2353
rect 8650 -2405 8702 -2353
rect 8646 -2407 8702 -2405
rect 8726 -2353 8782 -2351
rect 8726 -2405 8730 -2353
rect 8730 -2405 8782 -2353
rect 8726 -2407 8782 -2405
rect 8806 -2353 8862 -2351
rect 8806 -2405 8810 -2353
rect 8810 -2405 8862 -2353
rect 8806 -2407 8862 -2405
rect 9014 -2353 9070 -2351
rect 9014 -2405 9066 -2353
rect 9066 -2405 9070 -2353
rect 9014 -2407 9070 -2405
rect 9094 -2353 9150 -2351
rect 9094 -2405 9146 -2353
rect 9146 -2405 9150 -2353
rect 9094 -2407 9150 -2405
rect 9174 -2353 9230 -2351
rect 9174 -2405 9226 -2353
rect 9226 -2405 9230 -2353
rect 9174 -2407 9230 -2405
rect 9254 -2353 9310 -2351
rect 9254 -2405 9306 -2353
rect 9306 -2405 9310 -2353
rect 9254 -2407 9310 -2405
rect 9334 -2353 9390 -2351
rect 9334 -2405 9386 -2353
rect 9386 -2405 9390 -2353
rect 9334 -2407 9390 -2405
rect 9414 -2353 9470 -2351
rect 9414 -2405 9466 -2353
rect 9466 -2405 9470 -2353
rect 9414 -2407 9470 -2405
rect 9618 -2353 9674 -2351
rect 9618 -2405 9622 -2353
rect 9622 -2405 9674 -2353
rect 9618 -2407 9674 -2405
rect 9698 -2353 9754 -2351
rect 9698 -2405 9702 -2353
rect 9702 -2405 9754 -2353
rect 9698 -2407 9754 -2405
rect 9778 -2353 9834 -2351
rect 9778 -2405 9782 -2353
rect 9782 -2405 9834 -2353
rect 9778 -2407 9834 -2405
rect 9858 -2353 9914 -2351
rect 9858 -2405 9862 -2353
rect 9862 -2405 9914 -2353
rect 9858 -2407 9914 -2405
rect 9938 -2353 9994 -2351
rect 9938 -2405 9942 -2353
rect 9942 -2405 9994 -2353
rect 9938 -2407 9994 -2405
rect 10018 -2353 10074 -2351
rect 10018 -2405 10022 -2353
rect 10022 -2405 10074 -2353
rect 10018 -2407 10074 -2405
rect 10226 -2353 10282 -2351
rect 10226 -2405 10278 -2353
rect 10278 -2405 10282 -2353
rect 10226 -2407 10282 -2405
rect 10306 -2353 10362 -2351
rect 10306 -2405 10358 -2353
rect 10358 -2405 10362 -2353
rect 10306 -2407 10362 -2405
rect 10386 -2353 10442 -2351
rect 10386 -2405 10438 -2353
rect 10438 -2405 10442 -2353
rect 10386 -2407 10442 -2405
rect 10466 -2353 10522 -2351
rect 10466 -2405 10518 -2353
rect 10518 -2405 10522 -2353
rect 10466 -2407 10522 -2405
rect 10546 -2353 10602 -2351
rect 10546 -2405 10598 -2353
rect 10598 -2405 10602 -2353
rect 10546 -2407 10602 -2405
rect 10626 -2353 10682 -2351
rect 10626 -2405 10678 -2353
rect 10678 -2405 10682 -2353
rect 10626 -2407 10682 -2405
rect 10830 -2353 10886 -2351
rect 10830 -2405 10834 -2353
rect 10834 -2405 10886 -2353
rect 10830 -2407 10886 -2405
rect 10910 -2353 10966 -2351
rect 10910 -2405 10914 -2353
rect 10914 -2405 10966 -2353
rect 10910 -2407 10966 -2405
rect 10990 -2353 11046 -2351
rect 10990 -2405 10994 -2353
rect 10994 -2405 11046 -2353
rect 10990 -2407 11046 -2405
rect 11070 -2353 11126 -2351
rect 11070 -2405 11074 -2353
rect 11074 -2405 11126 -2353
rect 11070 -2407 11126 -2405
rect 11150 -2353 11206 -2351
rect 11150 -2405 11154 -2353
rect 11154 -2405 11206 -2353
rect 11150 -2407 11206 -2405
rect 11230 -2353 11286 -2351
rect 11230 -2405 11234 -2353
rect 11234 -2405 11286 -2353
rect 11230 -2407 11286 -2405
rect 11438 -2353 11494 -2351
rect 11438 -2405 11490 -2353
rect 11490 -2405 11494 -2353
rect 11438 -2407 11494 -2405
rect 11518 -2353 11574 -2351
rect 11518 -2405 11570 -2353
rect 11570 -2405 11574 -2353
rect 11518 -2407 11574 -2405
rect 11598 -2353 11654 -2351
rect 11598 -2405 11650 -2353
rect 11650 -2405 11654 -2353
rect 11598 -2407 11654 -2405
rect 11678 -2353 11734 -2351
rect 11678 -2405 11730 -2353
rect 11730 -2405 11734 -2353
rect 11678 -2407 11734 -2405
rect 11758 -2353 11814 -2351
rect 11758 -2405 11810 -2353
rect 11810 -2405 11814 -2353
rect 11758 -2407 11814 -2405
rect 11838 -2353 11894 -2351
rect 11838 -2405 11890 -2353
rect 11890 -2405 11894 -2353
rect 11838 -2407 11894 -2405
rect 12170 -2350 12226 -2348
rect 12170 -2402 12222 -2350
rect 12222 -2402 12226 -2350
rect 12170 -2404 12226 -2402
rect 12250 -2350 12306 -2348
rect 12250 -2402 12302 -2350
rect 12302 -2402 12306 -2350
rect 12250 -2404 12306 -2402
rect 12330 -2350 12386 -2348
rect 12330 -2402 12382 -2350
rect 12382 -2402 12386 -2350
rect 12330 -2404 12386 -2402
rect 12410 -2350 12466 -2348
rect 12410 -2402 12462 -2350
rect 12462 -2402 12466 -2350
rect 12410 -2404 12466 -2402
rect 12490 -2350 12546 -2348
rect 12490 -2402 12542 -2350
rect 12542 -2402 12546 -2350
rect 12490 -2404 12546 -2402
rect 12570 -2350 12626 -2348
rect 12570 -2402 12622 -2350
rect 12622 -2402 12626 -2350
rect 12570 -2404 12626 -2402
rect 12666 -2359 12722 -2357
rect 12666 -2411 12668 -2359
rect 12668 -2411 12720 -2359
rect 12720 -2411 12722 -2359
rect 12666 -2413 12722 -2411
<< metal3 >>
rect 707 3738 833 3748
rect 707 3674 738 3738
rect 802 3730 833 3738
rect 7416 3738 7542 3748
rect 1463 3731 6377 3733
rect 802 3728 1403 3730
rect 802 3674 835 3728
rect 707 3665 835 3674
rect 731 3664 835 3665
rect 899 3664 915 3728
rect 979 3664 995 3728
rect 1059 3664 1075 3728
rect 1139 3664 1155 3728
rect 1219 3664 1235 3728
rect 1299 3664 1403 3728
rect 1463 3667 1567 3731
rect 1631 3667 1647 3731
rect 1711 3667 1727 3731
rect 1791 3667 1807 3731
rect 1871 3667 1887 3731
rect 1951 3667 1967 3731
rect 2031 3667 2173 3731
rect 2237 3667 2253 3731
rect 2317 3667 2333 3731
rect 2397 3667 2413 3731
rect 2477 3667 2493 3731
rect 2557 3667 2573 3731
rect 2637 3667 2779 3731
rect 2843 3667 2859 3731
rect 2923 3667 2939 3731
rect 3003 3667 3019 3731
rect 3083 3667 3099 3731
rect 3163 3667 3179 3731
rect 3243 3667 3385 3731
rect 3449 3667 3465 3731
rect 3529 3667 3545 3731
rect 3609 3667 3625 3731
rect 3689 3667 3705 3731
rect 3769 3667 3785 3731
rect 3849 3667 3991 3731
rect 4055 3667 4071 3731
rect 4135 3667 4151 3731
rect 4215 3667 4231 3731
rect 4295 3667 4311 3731
rect 4375 3667 4391 3731
rect 4455 3667 4597 3731
rect 4661 3667 4677 3731
rect 4741 3667 4757 3731
rect 4821 3667 4837 3731
rect 4901 3667 4917 3731
rect 4981 3667 4997 3731
rect 5061 3667 5203 3731
rect 5267 3667 5283 3731
rect 5347 3667 5363 3731
rect 5427 3667 5443 3731
rect 5507 3667 5523 3731
rect 5587 3667 5603 3731
rect 5667 3667 5809 3731
rect 5873 3667 5889 3731
rect 5953 3667 5969 3731
rect 6033 3667 6049 3731
rect 6113 3667 6129 3731
rect 6193 3667 6209 3731
rect 6273 3667 6377 3731
rect 1463 3665 6377 3667
rect 6516 3676 6642 3686
rect 731 3662 1403 3664
rect 731 3508 797 3598
rect 731 3444 732 3508
rect 796 3444 797 3508
rect 731 3428 797 3444
rect 731 3364 732 3428
rect 796 3364 797 3428
rect 731 3348 797 3364
rect 731 3284 732 3348
rect 796 3284 797 3348
rect 731 3268 797 3284
rect 731 3204 732 3268
rect 796 3204 797 3268
rect 731 3188 797 3204
rect 106 3147 224 3148
rect 355 3147 499 3148
rect 106 3133 499 3147
rect 106 3069 121 3133
rect 185 3132 396 3133
rect 185 3069 252 3132
rect 106 3068 252 3069
rect 316 3069 396 3132
rect 460 3069 499 3133
rect 316 3068 499 3069
rect 106 3052 499 3068
rect 731 3124 732 3188
rect 796 3124 797 3188
rect 731 3108 797 3124
rect 211 3051 355 3052
rect 731 3044 732 3108
rect 796 3044 797 3108
rect 731 3028 797 3044
rect 731 2964 732 3028
rect 796 2964 797 3028
rect 731 2948 797 2964
rect 731 2884 732 2948
rect 796 2884 797 2948
rect 731 2868 797 2884
rect 731 2804 732 2868
rect 796 2804 797 2868
rect 731 2788 797 2804
rect 731 2724 732 2788
rect 796 2724 797 2788
rect 246 2602 338 2603
rect 132 2587 505 2602
rect 132 2523 139 2587
rect 203 2523 259 2587
rect 323 2523 402 2587
rect 466 2523 505 2587
rect 132 2506 505 2523
rect 731 2570 797 2724
rect 857 2570 917 3602
rect 977 2632 1037 3662
rect 1097 2570 1157 3602
rect 1217 2632 1277 3662
rect 1337 3508 1403 3598
rect 1337 3444 1338 3508
rect 1402 3444 1403 3508
rect 1337 3428 1403 3444
rect 1337 3364 1338 3428
rect 1402 3364 1403 3428
rect 1337 3348 1403 3364
rect 1337 3284 1338 3348
rect 1402 3284 1403 3348
rect 1337 3268 1403 3284
rect 1337 3204 1338 3268
rect 1402 3204 1403 3268
rect 1337 3188 1403 3204
rect 1337 3124 1338 3188
rect 1402 3124 1403 3188
rect 1337 3108 1403 3124
rect 1337 3044 1338 3108
rect 1402 3044 1403 3108
rect 1337 3028 1403 3044
rect 1337 2964 1338 3028
rect 1402 2964 1403 3028
rect 1337 2948 1403 2964
rect 1337 2884 1338 2948
rect 1402 2884 1403 2948
rect 1337 2868 1403 2884
rect 1337 2804 1338 2868
rect 1402 2804 1403 2868
rect 1337 2788 1403 2804
rect 1337 2724 1338 2788
rect 1402 2724 1403 2788
rect 1337 2570 1403 2724
rect 731 2568 1403 2570
rect 731 2504 835 2568
rect 899 2504 915 2568
rect 979 2504 995 2568
rect 1059 2504 1075 2568
rect 1139 2504 1155 2568
rect 1219 2545 1235 2568
rect 1219 2504 1224 2545
rect 1299 2504 1403 2568
rect 1463 3511 1529 3601
rect 1463 3447 1464 3511
rect 1528 3447 1529 3511
rect 1463 3431 1529 3447
rect 1463 3367 1464 3431
rect 1528 3367 1529 3431
rect 1463 3351 1529 3367
rect 1463 3287 1464 3351
rect 1528 3287 1529 3351
rect 1463 3271 1529 3287
rect 1463 3207 1464 3271
rect 1528 3207 1529 3271
rect 1463 3191 1529 3207
rect 1463 3127 1464 3191
rect 1528 3127 1529 3191
rect 1463 3111 1529 3127
rect 1463 3047 1464 3111
rect 1528 3047 1529 3111
rect 1463 3031 1529 3047
rect 1463 2967 1464 3031
rect 1528 2967 1529 3031
rect 1463 2951 1529 2967
rect 1463 2887 1464 2951
rect 1528 2887 1529 2951
rect 1463 2871 1529 2887
rect 1463 2807 1464 2871
rect 1528 2807 1529 2871
rect 1463 2791 1529 2807
rect 1463 2727 1464 2791
rect 1528 2727 1529 2791
rect 1463 2573 1529 2727
rect 1589 2573 1649 3605
rect 1709 2635 1769 3665
rect 1829 2573 1889 3605
rect 1949 2635 2009 3665
rect 2069 3511 2135 3601
rect 2069 3447 2070 3511
rect 2134 3447 2135 3511
rect 2069 3431 2135 3447
rect 2069 3367 2070 3431
rect 2134 3367 2135 3431
rect 2069 3351 2135 3367
rect 2069 3287 2070 3351
rect 2134 3287 2135 3351
rect 2069 3271 2135 3287
rect 2069 3207 2070 3271
rect 2134 3207 2135 3271
rect 2069 3191 2135 3207
rect 2069 3127 2070 3191
rect 2134 3127 2135 3191
rect 2069 3111 2135 3127
rect 2069 3047 2070 3111
rect 2134 3047 2135 3111
rect 2069 3031 2135 3047
rect 2069 2967 2070 3031
rect 2134 2967 2135 3031
rect 2069 2951 2135 2967
rect 2069 2887 2070 2951
rect 2134 2887 2135 2951
rect 2069 2871 2135 2887
rect 2069 2807 2070 2871
rect 2134 2807 2135 2871
rect 2069 2791 2135 2807
rect 2069 2727 2070 2791
rect 2134 2727 2135 2791
rect 2069 2573 2135 2727
rect 2195 2635 2255 3665
rect 2315 2573 2375 3605
rect 2435 2635 2495 3665
rect 2555 2573 2615 3605
rect 2675 3511 2741 3601
rect 2675 3447 2676 3511
rect 2740 3447 2741 3511
rect 2675 3431 2741 3447
rect 2675 3367 2676 3431
rect 2740 3367 2741 3431
rect 2675 3351 2741 3367
rect 2675 3287 2676 3351
rect 2740 3287 2741 3351
rect 2675 3271 2741 3287
rect 2675 3207 2676 3271
rect 2740 3207 2741 3271
rect 2675 3191 2741 3207
rect 2675 3127 2676 3191
rect 2740 3127 2741 3191
rect 2675 3111 2741 3127
rect 2675 3047 2676 3111
rect 2740 3047 2741 3111
rect 2675 3031 2741 3047
rect 2675 2967 2676 3031
rect 2740 2967 2741 3031
rect 2675 2951 2741 2967
rect 2675 2887 2676 2951
rect 2740 2887 2741 2951
rect 2675 2871 2741 2887
rect 2675 2807 2676 2871
rect 2740 2807 2741 2871
rect 2675 2791 2741 2807
rect 2675 2727 2676 2791
rect 2740 2727 2741 2791
rect 2675 2573 2741 2727
rect 2801 2573 2861 3605
rect 2921 2635 2981 3665
rect 3041 2573 3101 3605
rect 3161 2635 3221 3665
rect 3281 3511 3347 3601
rect 3281 3447 3282 3511
rect 3346 3447 3347 3511
rect 3281 3431 3347 3447
rect 3281 3367 3282 3431
rect 3346 3367 3347 3431
rect 3281 3351 3347 3367
rect 3281 3287 3282 3351
rect 3346 3287 3347 3351
rect 3281 3271 3347 3287
rect 3281 3207 3282 3271
rect 3346 3207 3347 3271
rect 3281 3191 3347 3207
rect 3281 3127 3282 3191
rect 3346 3127 3347 3191
rect 3281 3111 3347 3127
rect 3281 3047 3282 3111
rect 3346 3047 3347 3111
rect 3281 3031 3347 3047
rect 3281 2967 3282 3031
rect 3346 2967 3347 3031
rect 3281 2951 3347 2967
rect 3281 2887 3282 2951
rect 3346 2887 3347 2951
rect 3281 2871 3347 2887
rect 3281 2807 3282 2871
rect 3346 2807 3347 2871
rect 3281 2791 3347 2807
rect 3281 2727 3282 2791
rect 3346 2727 3347 2791
rect 3281 2573 3347 2727
rect 3407 2635 3467 3665
rect 3527 2573 3587 3605
rect 3647 2635 3707 3665
rect 3767 2573 3827 3605
rect 3887 3511 3953 3601
rect 3887 3447 3888 3511
rect 3952 3447 3953 3511
rect 3887 3431 3953 3447
rect 3887 3367 3888 3431
rect 3952 3367 3953 3431
rect 3887 3351 3953 3367
rect 3887 3287 3888 3351
rect 3952 3287 3953 3351
rect 3887 3271 3953 3287
rect 3887 3207 3888 3271
rect 3952 3207 3953 3271
rect 3887 3191 3953 3207
rect 3887 3127 3888 3191
rect 3952 3127 3953 3191
rect 3887 3111 3953 3127
rect 3887 3047 3888 3111
rect 3952 3047 3953 3111
rect 3887 3031 3953 3047
rect 3887 2967 3888 3031
rect 3952 2967 3953 3031
rect 3887 2951 3953 2967
rect 3887 2887 3888 2951
rect 3952 2887 3953 2951
rect 3887 2871 3953 2887
rect 3887 2807 3888 2871
rect 3952 2807 3953 2871
rect 3887 2791 3953 2807
rect 3887 2727 3888 2791
rect 3952 2727 3953 2791
rect 3887 2573 3953 2727
rect 4013 2573 4073 3605
rect 4133 2635 4193 3665
rect 4253 2573 4313 3605
rect 4373 2635 4433 3665
rect 4493 3511 4559 3601
rect 4493 3447 4494 3511
rect 4558 3447 4559 3511
rect 4493 3431 4559 3447
rect 4493 3367 4494 3431
rect 4558 3367 4559 3431
rect 4493 3351 4559 3367
rect 4493 3287 4494 3351
rect 4558 3287 4559 3351
rect 4493 3271 4559 3287
rect 4493 3207 4494 3271
rect 4558 3207 4559 3271
rect 4493 3191 4559 3207
rect 4493 3127 4494 3191
rect 4558 3127 4559 3191
rect 4493 3111 4559 3127
rect 4493 3047 4494 3111
rect 4558 3047 4559 3111
rect 4493 3031 4559 3047
rect 4493 2967 4494 3031
rect 4558 2967 4559 3031
rect 4493 2951 4559 2967
rect 4493 2887 4494 2951
rect 4558 2887 4559 2951
rect 4493 2871 4559 2887
rect 4493 2807 4494 2871
rect 4558 2807 4559 2871
rect 4493 2791 4559 2807
rect 4493 2727 4494 2791
rect 4558 2727 4559 2791
rect 4493 2573 4559 2727
rect 4619 2635 4679 3665
rect 4739 2573 4799 3605
rect 4859 2635 4919 3665
rect 4979 2573 5039 3605
rect 5099 3511 5165 3601
rect 5099 3447 5100 3511
rect 5164 3447 5165 3511
rect 5099 3431 5165 3447
rect 5099 3367 5100 3431
rect 5164 3367 5165 3431
rect 5099 3351 5165 3367
rect 5099 3287 5100 3351
rect 5164 3287 5165 3351
rect 5099 3271 5165 3287
rect 5099 3207 5100 3271
rect 5164 3207 5165 3271
rect 5099 3191 5165 3207
rect 5099 3127 5100 3191
rect 5164 3127 5165 3191
rect 5099 3111 5165 3127
rect 5099 3047 5100 3111
rect 5164 3047 5165 3111
rect 5099 3031 5165 3047
rect 5099 2967 5100 3031
rect 5164 2967 5165 3031
rect 5099 2951 5165 2967
rect 5099 2887 5100 2951
rect 5164 2887 5165 2951
rect 5099 2871 5165 2887
rect 5099 2807 5100 2871
rect 5164 2807 5165 2871
rect 5099 2791 5165 2807
rect 5099 2727 5100 2791
rect 5164 2727 5165 2791
rect 5099 2573 5165 2727
rect 5225 2573 5285 3605
rect 5345 2635 5405 3665
rect 5465 2573 5525 3605
rect 5585 2635 5645 3665
rect 5705 3511 5771 3601
rect 5705 3447 5706 3511
rect 5770 3447 5771 3511
rect 5705 3431 5771 3447
rect 5705 3367 5706 3431
rect 5770 3367 5771 3431
rect 5705 3351 5771 3367
rect 5705 3287 5706 3351
rect 5770 3287 5771 3351
rect 5705 3271 5771 3287
rect 5705 3207 5706 3271
rect 5770 3207 5771 3271
rect 5705 3191 5771 3207
rect 5705 3127 5706 3191
rect 5770 3127 5771 3191
rect 5705 3111 5771 3127
rect 5705 3047 5706 3111
rect 5770 3047 5771 3111
rect 5705 3031 5771 3047
rect 5705 2967 5706 3031
rect 5770 2967 5771 3031
rect 5705 2951 5771 2967
rect 5705 2887 5706 2951
rect 5770 2887 5771 2951
rect 5705 2871 5771 2887
rect 5705 2807 5706 2871
rect 5770 2807 5771 2871
rect 5705 2791 5771 2807
rect 5705 2727 5706 2791
rect 5770 2727 5771 2791
rect 5705 2573 5771 2727
rect 5831 2635 5891 3665
rect 5951 2573 6011 3605
rect 6071 2635 6131 3665
rect 6516 3612 6547 3676
rect 6611 3612 6642 3676
rect 6191 2573 6251 3605
rect 6516 3602 6642 3612
rect 6993 3679 7119 3689
rect 6993 3615 7024 3679
rect 7088 3615 7119 3679
rect 7416 3674 7447 3738
rect 7511 3730 7542 3738
rect 8172 3731 13086 3733
rect 7511 3728 8112 3730
rect 7511 3674 7544 3728
rect 7416 3665 7544 3674
rect 7440 3664 7544 3665
rect 7608 3664 7624 3728
rect 7688 3664 7704 3728
rect 7768 3664 7784 3728
rect 7848 3664 7864 3728
rect 7928 3664 7944 3728
rect 8008 3664 8112 3728
rect 8172 3667 8276 3731
rect 8340 3667 8356 3731
rect 8420 3667 8436 3731
rect 8500 3667 8516 3731
rect 8580 3667 8596 3731
rect 8660 3667 8676 3731
rect 8740 3667 8882 3731
rect 8946 3667 8962 3731
rect 9026 3667 9042 3731
rect 9106 3667 9122 3731
rect 9186 3667 9202 3731
rect 9266 3667 9282 3731
rect 9346 3667 9488 3731
rect 9552 3667 9568 3731
rect 9632 3667 9648 3731
rect 9712 3667 9728 3731
rect 9792 3667 9808 3731
rect 9872 3667 9888 3731
rect 9952 3667 10094 3731
rect 10158 3667 10174 3731
rect 10238 3667 10254 3731
rect 10318 3667 10334 3731
rect 10398 3667 10414 3731
rect 10478 3667 10494 3731
rect 10558 3667 10700 3731
rect 10764 3667 10780 3731
rect 10844 3667 10860 3731
rect 10924 3667 10940 3731
rect 11004 3667 11020 3731
rect 11084 3667 11100 3731
rect 11164 3667 11306 3731
rect 11370 3667 11386 3731
rect 11450 3667 11466 3731
rect 11530 3667 11546 3731
rect 11610 3667 11626 3731
rect 11690 3667 11706 3731
rect 11770 3667 11912 3731
rect 11976 3667 11992 3731
rect 12056 3667 12072 3731
rect 12136 3667 12152 3731
rect 12216 3667 12232 3731
rect 12296 3667 12312 3731
rect 12376 3667 12518 3731
rect 12582 3667 12598 3731
rect 12662 3667 12678 3731
rect 12742 3667 12758 3731
rect 12822 3667 12838 3731
rect 12902 3667 12918 3731
rect 12982 3667 13086 3731
rect 8172 3665 13086 3667
rect 13225 3676 13351 3686
rect 7440 3662 8112 3664
rect 6993 3605 7119 3615
rect 6311 3511 6377 3601
rect 6311 3447 6312 3511
rect 6376 3447 6377 3511
rect 6521 3532 6647 3542
rect 6521 3468 6552 3532
rect 6616 3468 6647 3532
rect 6521 3458 6647 3468
rect 6982 3507 7108 3517
rect 6311 3431 6377 3447
rect 6982 3443 7013 3507
rect 7077 3443 7108 3507
rect 6982 3433 7108 3443
rect 7440 3508 7506 3598
rect 7440 3444 7441 3508
rect 7505 3444 7506 3508
rect 6311 3367 6312 3431
rect 6376 3367 6377 3431
rect 7440 3428 7506 3444
rect 6311 3351 6377 3367
rect 6311 3287 6312 3351
rect 6376 3287 6377 3351
rect 6522 3380 6648 3390
rect 6522 3316 6553 3380
rect 6617 3316 6648 3380
rect 7440 3364 7441 3428
rect 7505 3364 7506 3428
rect 7440 3348 7506 3364
rect 6522 3306 6648 3316
rect 6982 3315 7108 3325
rect 6311 3271 6377 3287
rect 6311 3207 6312 3271
rect 6376 3207 6377 3271
rect 6982 3251 7013 3315
rect 7077 3251 7108 3315
rect 6982 3241 7108 3251
rect 7440 3284 7441 3348
rect 7505 3284 7506 3348
rect 7440 3268 7506 3284
rect 6311 3191 6377 3207
rect 6311 3127 6312 3191
rect 6376 3127 6377 3191
rect 6522 3210 6648 3220
rect 6522 3146 6553 3210
rect 6617 3146 6648 3210
rect 7440 3204 7441 3268
rect 7505 3204 7506 3268
rect 7440 3188 7506 3204
rect 6522 3136 6648 3146
rect 6815 3147 6933 3148
rect 7064 3147 7208 3148
rect 6311 3111 6377 3127
rect 6311 3047 6312 3111
rect 6376 3047 6377 3111
rect 6815 3133 7208 3147
rect 6815 3069 6830 3133
rect 6894 3132 7105 3133
rect 6894 3069 6961 3132
rect 6815 3068 6961 3069
rect 7025 3069 7105 3132
rect 7169 3069 7208 3133
rect 7025 3068 7208 3069
rect 6311 3031 6377 3047
rect 6311 2967 6312 3031
rect 6376 2967 6377 3031
rect 6521 3053 6647 3063
rect 6521 2989 6552 3053
rect 6616 2989 6647 3053
rect 6815 3052 7208 3068
rect 7440 3124 7441 3188
rect 7505 3124 7506 3188
rect 7440 3108 7506 3124
rect 6920 3051 7064 3052
rect 6521 2979 6647 2989
rect 7440 3044 7441 3108
rect 7505 3044 7506 3108
rect 7440 3028 7506 3044
rect 6311 2951 6377 2967
rect 6311 2887 6312 2951
rect 6376 2887 6377 2951
rect 6311 2871 6377 2887
rect 6311 2807 6312 2871
rect 6376 2807 6377 2871
rect 7440 2964 7441 3028
rect 7505 2964 7506 3028
rect 7440 2948 7506 2964
rect 7440 2884 7441 2948
rect 7505 2884 7506 2948
rect 7440 2868 7506 2884
rect 6311 2791 6377 2807
rect 6311 2727 6312 2791
rect 6376 2727 6377 2791
rect 6439 2811 6565 2821
rect 6439 2747 6470 2811
rect 6534 2747 6565 2811
rect 6439 2737 6565 2747
rect 7440 2804 7441 2868
rect 7505 2804 7506 2868
rect 7440 2788 7506 2804
rect 6311 2573 6377 2727
rect 7440 2724 7441 2788
rect 7505 2724 7506 2788
rect 6955 2602 7047 2603
rect 1463 2571 6377 2573
rect 1463 2507 1567 2571
rect 1631 2507 1647 2571
rect 1711 2507 1727 2571
rect 1791 2507 1807 2571
rect 1871 2507 1887 2571
rect 1951 2548 1967 2571
rect 1951 2507 1956 2548
rect 2031 2507 2173 2571
rect 2237 2548 2253 2571
rect 2248 2507 2253 2548
rect 2317 2507 2333 2571
rect 2397 2507 2413 2571
rect 2477 2507 2493 2571
rect 2557 2507 2573 2571
rect 2637 2507 2779 2571
rect 2843 2507 2859 2571
rect 2923 2507 2939 2571
rect 3003 2507 3019 2571
rect 3083 2507 3099 2571
rect 3163 2548 3179 2571
rect 3163 2507 3168 2548
rect 3243 2507 3385 2571
rect 3449 2548 3465 2571
rect 3460 2507 3465 2548
rect 3529 2507 3545 2571
rect 3609 2507 3625 2571
rect 3689 2507 3705 2571
rect 3769 2507 3785 2571
rect 3849 2507 3991 2571
rect 4055 2507 4071 2571
rect 4135 2507 4151 2571
rect 4215 2507 4231 2571
rect 4295 2507 4311 2571
rect 4375 2548 4391 2571
rect 4375 2507 4380 2548
rect 4455 2507 4597 2571
rect 4661 2548 4677 2571
rect 4672 2507 4677 2548
rect 4741 2507 4757 2571
rect 4821 2507 4837 2571
rect 4901 2507 4917 2571
rect 4981 2507 4997 2571
rect 5061 2507 5203 2571
rect 5267 2507 5283 2571
rect 5347 2507 5363 2571
rect 5427 2507 5443 2571
rect 5507 2507 5523 2571
rect 5587 2548 5603 2571
rect 5587 2507 5592 2548
rect 5667 2507 5809 2571
rect 5873 2548 5889 2571
rect 5884 2507 5889 2548
rect 5953 2507 5969 2571
rect 6033 2507 6049 2571
rect 6113 2507 6129 2571
rect 6193 2507 6209 2571
rect 6273 2507 6377 2571
rect 6841 2587 7214 2602
rect 1463 2505 1956 2507
rect 731 2502 1224 2504
rect 1214 2481 1224 2502
rect 1288 2502 1403 2504
rect 1288 2481 1297 2502
rect 1214 2476 1297 2481
rect 1946 2484 1956 2505
rect 2020 2505 2184 2507
rect 2020 2484 2029 2505
rect 1946 2479 2029 2484
rect 2175 2484 2184 2505
rect 2248 2505 3168 2507
rect 2248 2484 2258 2505
rect 2175 2479 2258 2484
rect 3158 2484 3168 2505
rect 3232 2505 3396 2507
rect 3232 2484 3241 2505
rect 3158 2479 3241 2484
rect 3387 2484 3396 2505
rect 3460 2505 4380 2507
rect 3460 2484 3470 2505
rect 3387 2479 3470 2484
rect 4370 2484 4380 2505
rect 4444 2505 4608 2507
rect 4444 2484 4453 2505
rect 4370 2479 4453 2484
rect 4599 2484 4608 2505
rect 4672 2505 5592 2507
rect 4672 2484 4682 2505
rect 4599 2479 4682 2484
rect 5582 2484 5592 2505
rect 5656 2505 5820 2507
rect 5656 2484 5665 2505
rect 5582 2479 5665 2484
rect 5811 2484 5820 2505
rect 5884 2505 6377 2507
rect 6527 2550 6653 2560
rect 5884 2484 5894 2505
rect 5811 2479 5894 2484
rect 6527 2486 6558 2550
rect 6622 2486 6653 2550
rect 6841 2523 6848 2587
rect 6912 2523 6968 2587
rect 7032 2523 7111 2587
rect 7175 2523 7214 2587
rect 6841 2506 7214 2523
rect 7440 2570 7506 2724
rect 7566 2570 7626 3602
rect 7686 2632 7746 3662
rect 7806 2570 7866 3602
rect 7926 2632 7986 3662
rect 8046 3508 8112 3598
rect 8046 3444 8047 3508
rect 8111 3444 8112 3508
rect 8046 3428 8112 3444
rect 8046 3364 8047 3428
rect 8111 3364 8112 3428
rect 8046 3348 8112 3364
rect 8046 3284 8047 3348
rect 8111 3284 8112 3348
rect 8046 3268 8112 3284
rect 8046 3204 8047 3268
rect 8111 3204 8112 3268
rect 8046 3188 8112 3204
rect 8046 3124 8047 3188
rect 8111 3124 8112 3188
rect 8046 3108 8112 3124
rect 8046 3044 8047 3108
rect 8111 3044 8112 3108
rect 8046 3028 8112 3044
rect 8046 2964 8047 3028
rect 8111 2964 8112 3028
rect 8046 2948 8112 2964
rect 8046 2884 8047 2948
rect 8111 2884 8112 2948
rect 8046 2868 8112 2884
rect 8046 2804 8047 2868
rect 8111 2804 8112 2868
rect 8046 2788 8112 2804
rect 8046 2724 8047 2788
rect 8111 2724 8112 2788
rect 8046 2570 8112 2724
rect 7440 2568 8112 2570
rect 7440 2504 7544 2568
rect 7608 2504 7624 2568
rect 7688 2504 7704 2568
rect 7768 2504 7784 2568
rect 7848 2504 7864 2568
rect 7928 2545 7944 2568
rect 7928 2504 7933 2545
rect 8008 2504 8112 2568
rect 8172 3511 8238 3601
rect 8172 3447 8173 3511
rect 8237 3447 8238 3511
rect 8172 3431 8238 3447
rect 8172 3367 8173 3431
rect 8237 3367 8238 3431
rect 8172 3351 8238 3367
rect 8172 3287 8173 3351
rect 8237 3287 8238 3351
rect 8172 3271 8238 3287
rect 8172 3207 8173 3271
rect 8237 3207 8238 3271
rect 8172 3191 8238 3207
rect 8172 3127 8173 3191
rect 8237 3127 8238 3191
rect 8172 3111 8238 3127
rect 8172 3047 8173 3111
rect 8237 3047 8238 3111
rect 8172 3031 8238 3047
rect 8172 2967 8173 3031
rect 8237 2967 8238 3031
rect 8172 2951 8238 2967
rect 8172 2887 8173 2951
rect 8237 2887 8238 2951
rect 8172 2871 8238 2887
rect 8172 2807 8173 2871
rect 8237 2807 8238 2871
rect 8172 2791 8238 2807
rect 8172 2727 8173 2791
rect 8237 2727 8238 2791
rect 8172 2573 8238 2727
rect 8298 2573 8358 3605
rect 8418 2635 8478 3665
rect 8538 2573 8598 3605
rect 8658 2635 8718 3665
rect 8778 3511 8844 3601
rect 8778 3447 8779 3511
rect 8843 3447 8844 3511
rect 8778 3431 8844 3447
rect 8778 3367 8779 3431
rect 8843 3367 8844 3431
rect 8778 3351 8844 3367
rect 8778 3287 8779 3351
rect 8843 3287 8844 3351
rect 8778 3271 8844 3287
rect 8778 3207 8779 3271
rect 8843 3207 8844 3271
rect 8778 3191 8844 3207
rect 8778 3127 8779 3191
rect 8843 3127 8844 3191
rect 8778 3111 8844 3127
rect 8778 3047 8779 3111
rect 8843 3047 8844 3111
rect 8778 3031 8844 3047
rect 8778 2967 8779 3031
rect 8843 2967 8844 3031
rect 8778 2951 8844 2967
rect 8778 2887 8779 2951
rect 8843 2887 8844 2951
rect 8778 2871 8844 2887
rect 8778 2807 8779 2871
rect 8843 2807 8844 2871
rect 8778 2791 8844 2807
rect 8778 2727 8779 2791
rect 8843 2727 8844 2791
rect 8778 2573 8844 2727
rect 8904 2635 8964 3665
rect 9024 2573 9084 3605
rect 9144 2635 9204 3665
rect 9264 2573 9324 3605
rect 9384 3511 9450 3601
rect 9384 3447 9385 3511
rect 9449 3447 9450 3511
rect 9384 3431 9450 3447
rect 9384 3367 9385 3431
rect 9449 3367 9450 3431
rect 9384 3351 9450 3367
rect 9384 3287 9385 3351
rect 9449 3287 9450 3351
rect 9384 3271 9450 3287
rect 9384 3207 9385 3271
rect 9449 3207 9450 3271
rect 9384 3191 9450 3207
rect 9384 3127 9385 3191
rect 9449 3127 9450 3191
rect 9384 3111 9450 3127
rect 9384 3047 9385 3111
rect 9449 3047 9450 3111
rect 9384 3031 9450 3047
rect 9384 2967 9385 3031
rect 9449 2967 9450 3031
rect 9384 2951 9450 2967
rect 9384 2887 9385 2951
rect 9449 2887 9450 2951
rect 9384 2871 9450 2887
rect 9384 2807 9385 2871
rect 9449 2807 9450 2871
rect 9384 2791 9450 2807
rect 9384 2727 9385 2791
rect 9449 2727 9450 2791
rect 9384 2573 9450 2727
rect 9510 2573 9570 3605
rect 9630 2635 9690 3665
rect 9750 2573 9810 3605
rect 9870 2635 9930 3665
rect 9990 3511 10056 3601
rect 9990 3447 9991 3511
rect 10055 3447 10056 3511
rect 9990 3431 10056 3447
rect 9990 3367 9991 3431
rect 10055 3367 10056 3431
rect 9990 3351 10056 3367
rect 9990 3287 9991 3351
rect 10055 3287 10056 3351
rect 9990 3271 10056 3287
rect 9990 3207 9991 3271
rect 10055 3207 10056 3271
rect 9990 3191 10056 3207
rect 9990 3127 9991 3191
rect 10055 3127 10056 3191
rect 9990 3111 10056 3127
rect 9990 3047 9991 3111
rect 10055 3047 10056 3111
rect 9990 3031 10056 3047
rect 9990 2967 9991 3031
rect 10055 2967 10056 3031
rect 9990 2951 10056 2967
rect 9990 2887 9991 2951
rect 10055 2887 10056 2951
rect 9990 2871 10056 2887
rect 9990 2807 9991 2871
rect 10055 2807 10056 2871
rect 9990 2791 10056 2807
rect 9990 2727 9991 2791
rect 10055 2727 10056 2791
rect 9990 2573 10056 2727
rect 10116 2635 10176 3665
rect 10236 2573 10296 3605
rect 10356 2635 10416 3665
rect 10476 2573 10536 3605
rect 10596 3511 10662 3601
rect 10596 3447 10597 3511
rect 10661 3447 10662 3511
rect 10596 3431 10662 3447
rect 10596 3367 10597 3431
rect 10661 3367 10662 3431
rect 10596 3351 10662 3367
rect 10596 3287 10597 3351
rect 10661 3287 10662 3351
rect 10596 3271 10662 3287
rect 10596 3207 10597 3271
rect 10661 3207 10662 3271
rect 10596 3191 10662 3207
rect 10596 3127 10597 3191
rect 10661 3127 10662 3191
rect 10596 3111 10662 3127
rect 10596 3047 10597 3111
rect 10661 3047 10662 3111
rect 10596 3031 10662 3047
rect 10596 2967 10597 3031
rect 10661 2967 10662 3031
rect 10596 2951 10662 2967
rect 10596 2887 10597 2951
rect 10661 2887 10662 2951
rect 10596 2871 10662 2887
rect 10596 2807 10597 2871
rect 10661 2807 10662 2871
rect 10596 2791 10662 2807
rect 10596 2727 10597 2791
rect 10661 2727 10662 2791
rect 10596 2573 10662 2727
rect 10722 2573 10782 3605
rect 10842 2635 10902 3665
rect 10962 2573 11022 3605
rect 11082 2635 11142 3665
rect 11202 3511 11268 3601
rect 11202 3447 11203 3511
rect 11267 3447 11268 3511
rect 11202 3431 11268 3447
rect 11202 3367 11203 3431
rect 11267 3367 11268 3431
rect 11202 3351 11268 3367
rect 11202 3287 11203 3351
rect 11267 3287 11268 3351
rect 11202 3271 11268 3287
rect 11202 3207 11203 3271
rect 11267 3207 11268 3271
rect 11202 3191 11268 3207
rect 11202 3127 11203 3191
rect 11267 3127 11268 3191
rect 11202 3111 11268 3127
rect 11202 3047 11203 3111
rect 11267 3047 11268 3111
rect 11202 3031 11268 3047
rect 11202 2967 11203 3031
rect 11267 2967 11268 3031
rect 11202 2951 11268 2967
rect 11202 2887 11203 2951
rect 11267 2887 11268 2951
rect 11202 2871 11268 2887
rect 11202 2807 11203 2871
rect 11267 2807 11268 2871
rect 11202 2791 11268 2807
rect 11202 2727 11203 2791
rect 11267 2727 11268 2791
rect 11202 2573 11268 2727
rect 11328 2635 11388 3665
rect 11448 2573 11508 3605
rect 11568 2635 11628 3665
rect 11688 2573 11748 3605
rect 11808 3511 11874 3601
rect 11808 3447 11809 3511
rect 11873 3447 11874 3511
rect 11808 3431 11874 3447
rect 11808 3367 11809 3431
rect 11873 3367 11874 3431
rect 11808 3351 11874 3367
rect 11808 3287 11809 3351
rect 11873 3287 11874 3351
rect 11808 3271 11874 3287
rect 11808 3207 11809 3271
rect 11873 3207 11874 3271
rect 11808 3191 11874 3207
rect 11808 3127 11809 3191
rect 11873 3127 11874 3191
rect 11808 3111 11874 3127
rect 11808 3047 11809 3111
rect 11873 3047 11874 3111
rect 11808 3031 11874 3047
rect 11808 2967 11809 3031
rect 11873 2967 11874 3031
rect 11808 2951 11874 2967
rect 11808 2887 11809 2951
rect 11873 2887 11874 2951
rect 11808 2871 11874 2887
rect 11808 2807 11809 2871
rect 11873 2807 11874 2871
rect 11808 2791 11874 2807
rect 11808 2727 11809 2791
rect 11873 2727 11874 2791
rect 11808 2573 11874 2727
rect 11934 2573 11994 3605
rect 12054 2635 12114 3665
rect 12174 2573 12234 3605
rect 12294 2635 12354 3665
rect 12414 3511 12480 3601
rect 12414 3447 12415 3511
rect 12479 3447 12480 3511
rect 12414 3431 12480 3447
rect 12414 3367 12415 3431
rect 12479 3367 12480 3431
rect 12414 3351 12480 3367
rect 12414 3287 12415 3351
rect 12479 3287 12480 3351
rect 12414 3271 12480 3287
rect 12414 3207 12415 3271
rect 12479 3207 12480 3271
rect 12414 3191 12480 3207
rect 12414 3127 12415 3191
rect 12479 3127 12480 3191
rect 12414 3111 12480 3127
rect 12414 3047 12415 3111
rect 12479 3047 12480 3111
rect 12414 3031 12480 3047
rect 12414 2967 12415 3031
rect 12479 2967 12480 3031
rect 12414 2951 12480 2967
rect 12414 2887 12415 2951
rect 12479 2887 12480 2951
rect 12414 2871 12480 2887
rect 12414 2807 12415 2871
rect 12479 2807 12480 2871
rect 12414 2791 12480 2807
rect 12414 2727 12415 2791
rect 12479 2727 12480 2791
rect 12414 2573 12480 2727
rect 12540 2635 12600 3665
rect 12660 2573 12720 3605
rect 12780 2635 12840 3665
rect 13225 3612 13256 3676
rect 13320 3612 13351 3676
rect 12900 2573 12960 3605
rect 13225 3602 13351 3612
rect 13020 3511 13086 3601
rect 13020 3447 13021 3511
rect 13085 3447 13086 3511
rect 13230 3532 13356 3542
rect 13230 3468 13261 3532
rect 13325 3468 13356 3532
rect 13230 3458 13356 3468
rect 13020 3431 13086 3447
rect 13020 3367 13021 3431
rect 13085 3367 13086 3431
rect 13020 3351 13086 3367
rect 13020 3287 13021 3351
rect 13085 3287 13086 3351
rect 13231 3380 13357 3390
rect 13231 3316 13262 3380
rect 13326 3316 13357 3380
rect 13231 3306 13357 3316
rect 13020 3271 13086 3287
rect 13020 3207 13021 3271
rect 13085 3207 13086 3271
rect 13020 3191 13086 3207
rect 13020 3127 13021 3191
rect 13085 3127 13086 3191
rect 13231 3210 13357 3220
rect 13231 3146 13262 3210
rect 13326 3146 13357 3210
rect 13231 3136 13357 3146
rect 13020 3111 13086 3127
rect 13020 3047 13021 3111
rect 13085 3047 13086 3111
rect 13020 3031 13086 3047
rect 13020 2967 13021 3031
rect 13085 2967 13086 3031
rect 13230 3053 13356 3063
rect 13230 2989 13261 3053
rect 13325 2989 13356 3053
rect 13230 2979 13356 2989
rect 13020 2951 13086 2967
rect 13020 2887 13021 2951
rect 13085 2887 13086 2951
rect 13020 2871 13086 2887
rect 13020 2807 13021 2871
rect 13085 2807 13086 2871
rect 13020 2791 13086 2807
rect 13020 2727 13021 2791
rect 13085 2727 13086 2791
rect 13148 2811 13274 2821
rect 13148 2747 13179 2811
rect 13243 2747 13274 2811
rect 13148 2737 13274 2747
rect 13020 2573 13086 2727
rect 8172 2571 13086 2573
rect 8172 2507 8276 2571
rect 8340 2507 8356 2571
rect 8420 2507 8436 2571
rect 8500 2507 8516 2571
rect 8580 2507 8596 2571
rect 8660 2548 8676 2571
rect 8660 2507 8665 2548
rect 8740 2507 8882 2571
rect 8946 2548 8962 2571
rect 8957 2507 8962 2548
rect 9026 2507 9042 2571
rect 9106 2507 9122 2571
rect 9186 2507 9202 2571
rect 9266 2507 9282 2571
rect 9346 2507 9488 2571
rect 9552 2507 9568 2571
rect 9632 2507 9648 2571
rect 9712 2507 9728 2571
rect 9792 2507 9808 2571
rect 9872 2548 9888 2571
rect 9872 2507 9877 2548
rect 9952 2507 10094 2571
rect 10158 2548 10174 2571
rect 10169 2507 10174 2548
rect 10238 2507 10254 2571
rect 10318 2507 10334 2571
rect 10398 2507 10414 2571
rect 10478 2507 10494 2571
rect 10558 2507 10700 2571
rect 10764 2507 10780 2571
rect 10844 2507 10860 2571
rect 10924 2507 10940 2571
rect 11004 2507 11020 2571
rect 11084 2548 11100 2571
rect 11084 2507 11089 2548
rect 11164 2507 11306 2571
rect 11370 2548 11386 2571
rect 11381 2507 11386 2548
rect 11450 2507 11466 2571
rect 11530 2507 11546 2571
rect 11610 2507 11626 2571
rect 11690 2507 11706 2571
rect 11770 2507 11912 2571
rect 11976 2507 11992 2571
rect 12056 2507 12072 2571
rect 12136 2507 12152 2571
rect 12216 2507 12232 2571
rect 12296 2548 12312 2571
rect 12296 2507 12301 2548
rect 12376 2507 12518 2571
rect 12582 2548 12598 2571
rect 12593 2507 12598 2548
rect 12662 2507 12678 2571
rect 12742 2507 12758 2571
rect 12822 2507 12838 2571
rect 12902 2507 12918 2571
rect 12982 2507 13086 2571
rect 8172 2505 8665 2507
rect 7440 2502 7933 2504
rect 6527 2476 6653 2486
rect 7923 2481 7933 2502
rect 7997 2502 8112 2504
rect 7997 2481 8006 2502
rect 7923 2476 8006 2481
rect 8655 2484 8665 2505
rect 8729 2505 8893 2507
rect 8729 2484 8738 2505
rect 8655 2479 8738 2484
rect 8884 2484 8893 2505
rect 8957 2505 9877 2507
rect 8957 2484 8967 2505
rect 8884 2479 8967 2484
rect 9867 2484 9877 2505
rect 9941 2505 10105 2507
rect 9941 2484 9950 2505
rect 9867 2479 9950 2484
rect 10096 2484 10105 2505
rect 10169 2505 11089 2507
rect 10169 2484 10179 2505
rect 10096 2479 10179 2484
rect 11079 2484 11089 2505
rect 11153 2505 11317 2507
rect 11153 2484 11162 2505
rect 11079 2479 11162 2484
rect 11308 2484 11317 2505
rect 11381 2505 12301 2507
rect 11381 2484 11391 2505
rect 11308 2479 11391 2484
rect 12291 2484 12301 2505
rect 12365 2505 12529 2507
rect 12365 2484 12374 2505
rect 12291 2479 12374 2484
rect 12520 2484 12529 2505
rect 12593 2505 13086 2507
rect 13236 2550 13362 2560
rect 12593 2484 12603 2505
rect 12520 2479 12603 2484
rect 13236 2486 13267 2550
rect 13331 2486 13362 2550
rect 13236 2476 13362 2486
rect 1571 2346 1653 2352
rect 1571 2325 1580 2346
rect 1082 2323 1580 2325
rect 1644 2325 1653 2346
rect 2303 2346 2385 2352
rect 2303 2325 2312 2346
rect 1644 2323 1754 2325
rect 1082 2259 1186 2323
rect 1250 2259 1266 2323
rect 1330 2259 1346 2323
rect 1410 2259 1426 2323
rect 1490 2259 1506 2323
rect 1570 2282 1580 2323
rect 1570 2259 1586 2282
rect 1650 2259 1754 2323
rect 1082 2257 1754 2259
rect 1082 2103 1148 2257
rect 1082 2039 1083 2103
rect 1147 2039 1148 2103
rect 1082 2023 1148 2039
rect 1082 1959 1083 2023
rect 1147 1959 1148 2023
rect 1082 1943 1148 1959
rect 1082 1879 1083 1943
rect 1147 1879 1148 1943
rect 1082 1863 1148 1879
rect 1082 1799 1083 1863
rect 1147 1799 1148 1863
rect 1082 1783 1148 1799
rect 49 1707 213 1734
rect 49 1701 106 1707
rect 49 1643 102 1701
rect 171 1643 213 1707
rect 49 1612 213 1643
rect 1082 1719 1083 1783
rect 1147 1719 1148 1783
rect 1082 1703 1148 1719
rect 1082 1639 1083 1703
rect 1147 1639 1148 1703
rect 1082 1623 1148 1639
rect 1082 1559 1083 1623
rect 1147 1559 1148 1623
rect 1082 1543 1148 1559
rect 1082 1479 1083 1543
rect 1147 1479 1148 1543
rect 1082 1463 1148 1479
rect 1082 1399 1083 1463
rect 1147 1399 1148 1463
rect 1082 1383 1148 1399
rect 1082 1319 1083 1383
rect 1147 1319 1148 1383
rect 1082 1229 1148 1319
rect 1208 1225 1268 2257
rect 694 1160 819 1170
rect 1328 1165 1388 2195
rect 1448 1225 1508 2257
rect 1568 1165 1628 2195
rect 1688 2103 1754 2257
rect 1688 2039 1689 2103
rect 1753 2039 1754 2103
rect 1688 2023 1754 2039
rect 1688 1959 1689 2023
rect 1753 1959 1754 2023
rect 1688 1943 1754 1959
rect 1688 1879 1689 1943
rect 1753 1879 1754 1943
rect 1688 1863 1754 1879
rect 1688 1799 1689 1863
rect 1753 1799 1754 1863
rect 1688 1783 1754 1799
rect 1688 1719 1689 1783
rect 1753 1719 1754 1783
rect 1688 1703 1754 1719
rect 1688 1639 1689 1703
rect 1753 1639 1754 1703
rect 1688 1623 1754 1639
rect 1688 1559 1689 1623
rect 1753 1559 1754 1623
rect 1688 1543 1754 1559
rect 1688 1479 1689 1543
rect 1753 1479 1754 1543
rect 1688 1463 1754 1479
rect 1688 1399 1689 1463
rect 1753 1399 1754 1463
rect 1688 1383 1754 1399
rect 1688 1319 1689 1383
rect 1753 1319 1754 1383
rect 1688 1229 1754 1319
rect 1814 2323 2312 2325
rect 2376 2325 2385 2346
rect 2521 2346 2603 2352
rect 2521 2325 2530 2346
rect 2376 2323 2530 2325
rect 2594 2325 2603 2346
rect 3515 2346 3597 2352
rect 3515 2325 3524 2346
rect 2594 2323 3524 2325
rect 3588 2325 3597 2346
rect 3733 2346 3815 2352
rect 3733 2325 3742 2346
rect 3588 2323 3742 2325
rect 3806 2325 3815 2346
rect 4853 2346 4935 2352
rect 4853 2325 4862 2346
rect 3806 2323 4304 2325
rect 1814 2259 1918 2323
rect 1982 2259 1998 2323
rect 2062 2259 2078 2323
rect 2142 2259 2158 2323
rect 2222 2259 2238 2323
rect 2302 2282 2312 2323
rect 2302 2259 2318 2282
rect 2382 2259 2524 2323
rect 2594 2282 2604 2323
rect 2588 2259 2604 2282
rect 2668 2259 2684 2323
rect 2748 2259 2764 2323
rect 2828 2259 2844 2323
rect 2908 2259 2924 2323
rect 2988 2259 3130 2323
rect 3194 2259 3210 2323
rect 3274 2259 3290 2323
rect 3354 2259 3370 2323
rect 3434 2259 3450 2323
rect 3514 2282 3524 2323
rect 3514 2259 3530 2282
rect 3594 2259 3736 2323
rect 3806 2282 3816 2323
rect 3800 2259 3816 2282
rect 3880 2259 3896 2323
rect 3960 2259 3976 2323
rect 4040 2259 4056 2323
rect 4120 2259 4136 2323
rect 4200 2259 4304 2323
rect 1814 2257 4304 2259
rect 1814 2103 1880 2257
rect 1814 2039 1815 2103
rect 1879 2039 1880 2103
rect 1814 2023 1880 2039
rect 1814 1959 1815 2023
rect 1879 1959 1880 2023
rect 1814 1943 1880 1959
rect 1814 1879 1815 1943
rect 1879 1879 1880 1943
rect 1814 1863 1880 1879
rect 1814 1799 1815 1863
rect 1879 1799 1880 1863
rect 1814 1783 1880 1799
rect 1814 1719 1815 1783
rect 1879 1719 1880 1783
rect 1814 1703 1880 1719
rect 1814 1639 1815 1703
rect 1879 1639 1880 1703
rect 1814 1623 1880 1639
rect 1814 1559 1815 1623
rect 1879 1559 1880 1623
rect 1814 1543 1880 1559
rect 1814 1479 1815 1543
rect 1879 1479 1880 1543
rect 1814 1463 1880 1479
rect 1814 1399 1815 1463
rect 1879 1399 1880 1463
rect 1814 1383 1880 1399
rect 1814 1319 1815 1383
rect 1879 1319 1880 1383
rect 1814 1229 1880 1319
rect 1940 1225 2000 2257
rect 2060 1165 2120 2195
rect 2180 1225 2240 2257
rect 2300 1165 2360 2195
rect 2420 2103 2486 2257
rect 2420 2039 2421 2103
rect 2485 2039 2486 2103
rect 2420 2023 2486 2039
rect 2420 1959 2421 2023
rect 2485 1959 2486 2023
rect 2420 1943 2486 1959
rect 2420 1879 2421 1943
rect 2485 1879 2486 1943
rect 2420 1863 2486 1879
rect 2420 1799 2421 1863
rect 2485 1799 2486 1863
rect 2420 1783 2486 1799
rect 2420 1719 2421 1783
rect 2485 1719 2486 1783
rect 2420 1703 2486 1719
rect 2420 1639 2421 1703
rect 2485 1639 2486 1703
rect 2420 1623 2486 1639
rect 2420 1559 2421 1623
rect 2485 1559 2486 1623
rect 2420 1543 2486 1559
rect 2420 1479 2421 1543
rect 2485 1479 2486 1543
rect 2420 1463 2486 1479
rect 2420 1399 2421 1463
rect 2485 1399 2486 1463
rect 2420 1383 2486 1399
rect 2420 1319 2421 1383
rect 2485 1319 2486 1383
rect 2420 1229 2486 1319
rect 2546 1165 2606 2195
rect 2666 1225 2726 2257
rect 2786 1165 2846 2195
rect 2906 1225 2966 2257
rect 3026 2103 3092 2257
rect 3026 2039 3027 2103
rect 3091 2039 3092 2103
rect 3026 2023 3092 2039
rect 3026 1959 3027 2023
rect 3091 1959 3092 2023
rect 3026 1943 3092 1959
rect 3026 1879 3027 1943
rect 3091 1879 3092 1943
rect 3026 1863 3092 1879
rect 3026 1799 3027 1863
rect 3091 1799 3092 1863
rect 3026 1783 3092 1799
rect 3026 1719 3027 1783
rect 3091 1719 3092 1783
rect 3026 1703 3092 1719
rect 3026 1639 3027 1703
rect 3091 1639 3092 1703
rect 3026 1623 3092 1639
rect 3026 1559 3027 1623
rect 3091 1559 3092 1623
rect 3026 1543 3092 1559
rect 3026 1479 3027 1543
rect 3091 1479 3092 1543
rect 3026 1463 3092 1479
rect 3026 1399 3027 1463
rect 3091 1399 3092 1463
rect 3026 1383 3092 1399
rect 3026 1319 3027 1383
rect 3091 1319 3092 1383
rect 3026 1229 3092 1319
rect 3152 1225 3212 2257
rect 3272 1165 3332 2195
rect 3392 1225 3452 2257
rect 3512 1165 3572 2195
rect 3632 2103 3698 2257
rect 3632 2039 3633 2103
rect 3697 2039 3698 2103
rect 3632 2023 3698 2039
rect 3632 1959 3633 2023
rect 3697 1959 3698 2023
rect 3632 1943 3698 1959
rect 3632 1879 3633 1943
rect 3697 1879 3698 1943
rect 3632 1863 3698 1879
rect 3632 1799 3633 1863
rect 3697 1799 3698 1863
rect 3632 1783 3698 1799
rect 3632 1719 3633 1783
rect 3697 1719 3698 1783
rect 3632 1703 3698 1719
rect 3632 1639 3633 1703
rect 3697 1639 3698 1703
rect 3632 1623 3698 1639
rect 3632 1559 3633 1623
rect 3697 1559 3698 1623
rect 3632 1543 3698 1559
rect 3632 1479 3633 1543
rect 3697 1479 3698 1543
rect 3632 1463 3698 1479
rect 3632 1399 3633 1463
rect 3697 1399 3698 1463
rect 3632 1383 3698 1399
rect 3632 1319 3633 1383
rect 3697 1319 3698 1383
rect 3632 1229 3698 1319
rect 3758 1165 3818 2195
rect 3878 1225 3938 2257
rect 3998 1165 4058 2195
rect 4118 1225 4178 2257
rect 4238 2103 4304 2257
rect 4238 2039 4239 2103
rect 4303 2039 4304 2103
rect 4238 2023 4304 2039
rect 4238 1959 4239 2023
rect 4303 1959 4304 2023
rect 4238 1943 4304 1959
rect 4238 1879 4239 1943
rect 4303 1879 4304 1943
rect 4238 1863 4304 1879
rect 4238 1799 4239 1863
rect 4303 1799 4304 1863
rect 4238 1783 4304 1799
rect 4238 1719 4239 1783
rect 4303 1719 4304 1783
rect 4238 1703 4304 1719
rect 4238 1639 4239 1703
rect 4303 1639 4304 1703
rect 4238 1623 4304 1639
rect 4238 1559 4239 1623
rect 4303 1559 4304 1623
rect 4238 1543 4304 1559
rect 4238 1479 4239 1543
rect 4303 1479 4304 1543
rect 4238 1463 4304 1479
rect 4238 1399 4239 1463
rect 4303 1399 4304 1463
rect 4238 1383 4304 1399
rect 4238 1319 4239 1383
rect 4303 1319 4304 1383
rect 4238 1229 4304 1319
rect 4364 2323 4862 2325
rect 4926 2325 4935 2346
rect 5071 2346 5153 2352
rect 5071 2325 5080 2346
rect 4926 2323 5080 2325
rect 5144 2325 5153 2346
rect 5805 2346 5887 2352
rect 5805 2325 5814 2346
rect 5144 2323 5642 2325
rect 4364 2259 4468 2323
rect 4532 2259 4548 2323
rect 4612 2259 4628 2323
rect 4692 2259 4708 2323
rect 4772 2259 4788 2323
rect 4852 2282 4862 2323
rect 4852 2259 4868 2282
rect 4932 2259 5074 2323
rect 5144 2282 5154 2323
rect 5138 2259 5154 2282
rect 5218 2259 5234 2323
rect 5298 2259 5314 2323
rect 5378 2259 5394 2323
rect 5458 2259 5474 2323
rect 5538 2259 5642 2323
rect 4364 2257 5642 2259
rect 4364 2103 4430 2257
rect 4364 2039 4365 2103
rect 4429 2039 4430 2103
rect 4364 2023 4430 2039
rect 4364 1959 4365 2023
rect 4429 1959 4430 2023
rect 4364 1943 4430 1959
rect 4364 1879 4365 1943
rect 4429 1879 4430 1943
rect 4364 1863 4430 1879
rect 4364 1799 4365 1863
rect 4429 1799 4430 1863
rect 4364 1783 4430 1799
rect 4364 1719 4365 1783
rect 4429 1719 4430 1783
rect 4364 1703 4430 1719
rect 4364 1639 4365 1703
rect 4429 1639 4430 1703
rect 4364 1623 4430 1639
rect 4364 1559 4365 1623
rect 4429 1559 4430 1623
rect 4364 1543 4430 1559
rect 4364 1479 4365 1543
rect 4429 1479 4430 1543
rect 4364 1463 4430 1479
rect 4364 1399 4365 1463
rect 4429 1399 4430 1463
rect 4364 1383 4430 1399
rect 4364 1319 4365 1383
rect 4429 1319 4430 1383
rect 4364 1229 4430 1319
rect 4490 1225 4550 2257
rect 4610 1165 4670 2195
rect 4730 1225 4790 2257
rect 4850 1165 4910 2195
rect 4970 2103 5036 2257
rect 4970 2039 4971 2103
rect 5035 2039 5036 2103
rect 4970 2023 5036 2039
rect 4970 1959 4971 2023
rect 5035 1959 5036 2023
rect 4970 1943 5036 1959
rect 4970 1879 4971 1943
rect 5035 1879 5036 1943
rect 4970 1863 5036 1879
rect 4970 1799 4971 1863
rect 5035 1799 5036 1863
rect 4970 1783 5036 1799
rect 4970 1719 4971 1783
rect 5035 1719 5036 1783
rect 4970 1703 5036 1719
rect 4970 1639 4971 1703
rect 5035 1639 5036 1703
rect 4970 1623 5036 1639
rect 4970 1559 4971 1623
rect 5035 1559 5036 1623
rect 4970 1543 5036 1559
rect 4970 1479 4971 1543
rect 5035 1479 5036 1543
rect 4970 1463 5036 1479
rect 4970 1399 4971 1463
rect 5035 1399 5036 1463
rect 4970 1383 5036 1399
rect 4970 1319 4971 1383
rect 5035 1319 5036 1383
rect 4970 1229 5036 1319
rect 5096 1165 5156 2195
rect 5216 1225 5276 2257
rect 5336 1165 5396 2195
rect 5456 1225 5516 2257
rect 5576 2103 5642 2257
rect 5576 2039 5577 2103
rect 5641 2039 5642 2103
rect 5576 2023 5642 2039
rect 5576 1959 5577 2023
rect 5641 1959 5642 2023
rect 5576 1943 5642 1959
rect 5576 1879 5577 1943
rect 5641 1879 5642 1943
rect 5576 1863 5642 1879
rect 5576 1799 5577 1863
rect 5641 1799 5642 1863
rect 5576 1783 5642 1799
rect 5576 1719 5577 1783
rect 5641 1719 5642 1783
rect 5576 1703 5642 1719
rect 5576 1639 5577 1703
rect 5641 1639 5642 1703
rect 5576 1623 5642 1639
rect 5576 1559 5577 1623
rect 5641 1559 5642 1623
rect 5576 1543 5642 1559
rect 5576 1479 5577 1543
rect 5641 1479 5642 1543
rect 5576 1463 5642 1479
rect 5576 1399 5577 1463
rect 5641 1399 5642 1463
rect 5576 1383 5642 1399
rect 5576 1319 5577 1383
rect 5641 1319 5642 1383
rect 5576 1229 5642 1319
rect 5704 2323 5814 2325
rect 5878 2325 5887 2346
rect 6527 2347 6653 2357
rect 5878 2323 6376 2325
rect 5704 2259 5808 2323
rect 5878 2282 5888 2323
rect 5872 2259 5888 2282
rect 5952 2259 5968 2323
rect 6032 2259 6048 2323
rect 6112 2259 6128 2323
rect 6192 2259 6208 2323
rect 6272 2259 6376 2323
rect 6527 2283 6558 2347
rect 6622 2283 6653 2347
rect 8280 2346 8362 2352
rect 8280 2325 8289 2346
rect 6527 2273 6653 2283
rect 7791 2323 8289 2325
rect 8353 2325 8362 2346
rect 9012 2346 9094 2352
rect 9012 2325 9021 2346
rect 8353 2323 8463 2325
rect 6553 2272 6627 2273
rect 5704 2257 6376 2259
rect 5704 2103 5770 2257
rect 5704 2039 5705 2103
rect 5769 2039 5770 2103
rect 5704 2023 5770 2039
rect 5704 1959 5705 2023
rect 5769 1959 5770 2023
rect 5704 1943 5770 1959
rect 5704 1879 5705 1943
rect 5769 1879 5770 1943
rect 5704 1863 5770 1879
rect 5704 1799 5705 1863
rect 5769 1799 5770 1863
rect 5704 1783 5770 1799
rect 5704 1719 5705 1783
rect 5769 1719 5770 1783
rect 5704 1703 5770 1719
rect 5704 1639 5705 1703
rect 5769 1639 5770 1703
rect 5704 1623 5770 1639
rect 5704 1559 5705 1623
rect 5769 1559 5770 1623
rect 5704 1543 5770 1559
rect 5704 1479 5705 1543
rect 5769 1479 5770 1543
rect 5704 1463 5770 1479
rect 5704 1399 5705 1463
rect 5769 1399 5770 1463
rect 5704 1383 5770 1399
rect 5704 1319 5705 1383
rect 5769 1319 5770 1383
rect 5704 1229 5770 1319
rect 5830 1165 5890 2195
rect 5950 1225 6010 2257
rect 6070 1165 6130 2195
rect 6190 1225 6250 2257
rect 6310 2103 6376 2257
rect 6310 2039 6311 2103
rect 6375 2039 6376 2103
rect 7791 2259 7895 2323
rect 7959 2259 7975 2323
rect 8039 2259 8055 2323
rect 8119 2259 8135 2323
rect 8199 2259 8215 2323
rect 8279 2282 8289 2323
rect 8279 2259 8295 2282
rect 8359 2259 8463 2323
rect 7791 2257 8463 2259
rect 7791 2103 7857 2257
rect 6310 2023 6376 2039
rect 6310 1959 6311 2023
rect 6375 1959 6376 2023
rect 6437 2085 6562 2095
rect 6437 2021 6467 2085
rect 6531 2021 6562 2085
rect 6437 2011 6562 2021
rect 7791 2039 7792 2103
rect 7856 2039 7857 2103
rect 7791 2023 7857 2039
rect 6310 1943 6376 1959
rect 6310 1879 6311 1943
rect 6375 1879 6376 1943
rect 6310 1863 6376 1879
rect 6310 1799 6311 1863
rect 6375 1799 6376 1863
rect 6310 1783 6376 1799
rect 6310 1719 6311 1783
rect 6375 1719 6376 1783
rect 6310 1703 6376 1719
rect 6310 1639 6311 1703
rect 6375 1639 6376 1703
rect 6310 1623 6376 1639
rect 6310 1559 6311 1623
rect 6375 1559 6376 1623
rect 6310 1543 6376 1559
rect 6310 1479 6311 1543
rect 6375 1479 6376 1543
rect 6310 1463 6376 1479
rect 6310 1399 6311 1463
rect 6375 1399 6376 1463
rect 6310 1383 6376 1399
rect 6310 1319 6311 1383
rect 6375 1319 6376 1383
rect 6310 1229 6376 1319
rect 7791 1959 7792 2023
rect 7856 1959 7857 2023
rect 7791 1943 7857 1959
rect 7791 1879 7792 1943
rect 7856 1879 7857 1943
rect 7791 1863 7857 1879
rect 7791 1799 7792 1863
rect 7856 1799 7857 1863
rect 7791 1783 7857 1799
rect 7791 1719 7792 1783
rect 7856 1719 7857 1783
rect 7791 1703 7857 1719
rect 7791 1639 7792 1703
rect 7856 1639 7857 1703
rect 7791 1623 7857 1639
rect 7791 1559 7792 1623
rect 7856 1559 7857 1623
rect 7791 1543 7857 1559
rect 7791 1479 7792 1543
rect 7856 1479 7857 1543
rect 7791 1463 7857 1479
rect 7791 1399 7792 1463
rect 7856 1399 7857 1463
rect 7791 1383 7857 1399
rect 7791 1319 7792 1383
rect 7856 1319 7857 1383
rect 7791 1229 7857 1319
rect 7917 1225 7977 2257
rect 694 1096 724 1160
rect 788 1096 819 1160
rect 1082 1163 1754 1165
rect 1082 1099 1266 1163
rect 1330 1099 1346 1163
rect 1410 1099 1426 1163
rect 1490 1099 1506 1163
rect 1570 1099 1754 1163
rect 1082 1097 1754 1099
rect 1814 1163 4304 1165
rect 1814 1099 1998 1163
rect 2062 1099 2078 1163
rect 2142 1099 2158 1163
rect 2222 1099 2238 1163
rect 2302 1099 2604 1163
rect 2668 1099 2684 1163
rect 2748 1099 2764 1163
rect 2828 1099 2844 1163
rect 2908 1099 3210 1163
rect 3274 1099 3290 1163
rect 3354 1099 3370 1163
rect 3434 1099 3450 1163
rect 3514 1099 3816 1163
rect 3880 1099 3896 1163
rect 3960 1099 3976 1163
rect 4040 1099 4056 1163
rect 4120 1099 4304 1163
rect 1814 1097 4304 1099
rect 4364 1163 5642 1165
rect 4364 1099 4548 1163
rect 4612 1099 4628 1163
rect 4692 1099 4708 1163
rect 4772 1099 4788 1163
rect 4852 1099 5154 1163
rect 5218 1099 5234 1163
rect 5298 1099 5314 1163
rect 5378 1099 5394 1163
rect 5458 1099 5642 1163
rect 4364 1097 5642 1099
rect 5704 1163 6376 1165
rect 5704 1099 5888 1163
rect 5952 1099 5968 1163
rect 6032 1099 6048 1163
rect 6112 1099 6128 1163
rect 6192 1099 6376 1163
rect 5704 1097 6376 1099
rect 7403 1160 7528 1170
rect 8037 1165 8097 2195
rect 8157 1225 8217 2257
rect 8277 1165 8337 2195
rect 8397 2103 8463 2257
rect 8397 2039 8398 2103
rect 8462 2039 8463 2103
rect 8397 2023 8463 2039
rect 8397 1959 8398 2023
rect 8462 1959 8463 2023
rect 8397 1943 8463 1959
rect 8397 1879 8398 1943
rect 8462 1879 8463 1943
rect 8397 1863 8463 1879
rect 8397 1799 8398 1863
rect 8462 1799 8463 1863
rect 8397 1783 8463 1799
rect 8397 1719 8398 1783
rect 8462 1719 8463 1783
rect 8397 1703 8463 1719
rect 8397 1639 8398 1703
rect 8462 1639 8463 1703
rect 8397 1623 8463 1639
rect 8397 1559 8398 1623
rect 8462 1559 8463 1623
rect 8397 1543 8463 1559
rect 8397 1479 8398 1543
rect 8462 1479 8463 1543
rect 8397 1463 8463 1479
rect 8397 1399 8398 1463
rect 8462 1399 8463 1463
rect 8397 1383 8463 1399
rect 8397 1319 8398 1383
rect 8462 1319 8463 1383
rect 8397 1229 8463 1319
rect 8523 2323 9021 2325
rect 9085 2325 9094 2346
rect 9230 2346 9312 2352
rect 9230 2325 9239 2346
rect 9085 2323 9239 2325
rect 9303 2325 9312 2346
rect 10224 2346 10306 2352
rect 10224 2325 10233 2346
rect 9303 2323 10233 2325
rect 10297 2325 10306 2346
rect 10442 2346 10524 2352
rect 10442 2325 10451 2346
rect 10297 2323 10451 2325
rect 10515 2325 10524 2346
rect 11562 2346 11644 2352
rect 11562 2325 11571 2346
rect 10515 2323 11013 2325
rect 8523 2259 8627 2323
rect 8691 2259 8707 2323
rect 8771 2259 8787 2323
rect 8851 2259 8867 2323
rect 8931 2259 8947 2323
rect 9011 2282 9021 2323
rect 9011 2259 9027 2282
rect 9091 2259 9233 2323
rect 9303 2282 9313 2323
rect 9297 2259 9313 2282
rect 9377 2259 9393 2323
rect 9457 2259 9473 2323
rect 9537 2259 9553 2323
rect 9617 2259 9633 2323
rect 9697 2259 9839 2323
rect 9903 2259 9919 2323
rect 9983 2259 9999 2323
rect 10063 2259 10079 2323
rect 10143 2259 10159 2323
rect 10223 2282 10233 2323
rect 10223 2259 10239 2282
rect 10303 2259 10445 2323
rect 10515 2282 10525 2323
rect 10509 2259 10525 2282
rect 10589 2259 10605 2323
rect 10669 2259 10685 2323
rect 10749 2259 10765 2323
rect 10829 2259 10845 2323
rect 10909 2259 11013 2323
rect 8523 2257 11013 2259
rect 8523 2103 8589 2257
rect 8523 2039 8524 2103
rect 8588 2039 8589 2103
rect 8523 2023 8589 2039
rect 8523 1959 8524 2023
rect 8588 1959 8589 2023
rect 8523 1943 8589 1959
rect 8523 1879 8524 1943
rect 8588 1879 8589 1943
rect 8523 1863 8589 1879
rect 8523 1799 8524 1863
rect 8588 1799 8589 1863
rect 8523 1783 8589 1799
rect 8523 1719 8524 1783
rect 8588 1719 8589 1783
rect 8523 1703 8589 1719
rect 8523 1639 8524 1703
rect 8588 1639 8589 1703
rect 8523 1623 8589 1639
rect 8523 1559 8524 1623
rect 8588 1559 8589 1623
rect 8523 1543 8589 1559
rect 8523 1479 8524 1543
rect 8588 1479 8589 1543
rect 8523 1463 8589 1479
rect 8523 1399 8524 1463
rect 8588 1399 8589 1463
rect 8523 1383 8589 1399
rect 8523 1319 8524 1383
rect 8588 1319 8589 1383
rect 8523 1229 8589 1319
rect 8649 1225 8709 2257
rect 8769 1165 8829 2195
rect 8889 1225 8949 2257
rect 9009 1165 9069 2195
rect 9129 2103 9195 2257
rect 9129 2039 9130 2103
rect 9194 2039 9195 2103
rect 9129 2023 9195 2039
rect 9129 1959 9130 2023
rect 9194 1959 9195 2023
rect 9129 1943 9195 1959
rect 9129 1879 9130 1943
rect 9194 1879 9195 1943
rect 9129 1863 9195 1879
rect 9129 1799 9130 1863
rect 9194 1799 9195 1863
rect 9129 1783 9195 1799
rect 9129 1719 9130 1783
rect 9194 1719 9195 1783
rect 9129 1703 9195 1719
rect 9129 1639 9130 1703
rect 9194 1639 9195 1703
rect 9129 1623 9195 1639
rect 9129 1559 9130 1623
rect 9194 1559 9195 1623
rect 9129 1543 9195 1559
rect 9129 1479 9130 1543
rect 9194 1479 9195 1543
rect 9129 1463 9195 1479
rect 9129 1399 9130 1463
rect 9194 1399 9195 1463
rect 9129 1383 9195 1399
rect 9129 1319 9130 1383
rect 9194 1319 9195 1383
rect 9129 1229 9195 1319
rect 9255 1165 9315 2195
rect 9375 1225 9435 2257
rect 9495 1165 9555 2195
rect 9615 1225 9675 2257
rect 9735 2103 9801 2257
rect 9735 2039 9736 2103
rect 9800 2039 9801 2103
rect 9735 2023 9801 2039
rect 9735 1959 9736 2023
rect 9800 1959 9801 2023
rect 9735 1943 9801 1959
rect 9735 1879 9736 1943
rect 9800 1879 9801 1943
rect 9735 1863 9801 1879
rect 9735 1799 9736 1863
rect 9800 1799 9801 1863
rect 9735 1783 9801 1799
rect 9735 1719 9736 1783
rect 9800 1719 9801 1783
rect 9735 1703 9801 1719
rect 9735 1639 9736 1703
rect 9800 1639 9801 1703
rect 9735 1623 9801 1639
rect 9735 1559 9736 1623
rect 9800 1559 9801 1623
rect 9735 1543 9801 1559
rect 9735 1479 9736 1543
rect 9800 1479 9801 1543
rect 9735 1463 9801 1479
rect 9735 1399 9736 1463
rect 9800 1399 9801 1463
rect 9735 1383 9801 1399
rect 9735 1319 9736 1383
rect 9800 1319 9801 1383
rect 9735 1229 9801 1319
rect 9861 1225 9921 2257
rect 9981 1165 10041 2195
rect 10101 1225 10161 2257
rect 10221 1165 10281 2195
rect 10341 2103 10407 2257
rect 10341 2039 10342 2103
rect 10406 2039 10407 2103
rect 10341 2023 10407 2039
rect 10341 1959 10342 2023
rect 10406 1959 10407 2023
rect 10341 1943 10407 1959
rect 10341 1879 10342 1943
rect 10406 1879 10407 1943
rect 10341 1863 10407 1879
rect 10341 1799 10342 1863
rect 10406 1799 10407 1863
rect 10341 1783 10407 1799
rect 10341 1719 10342 1783
rect 10406 1719 10407 1783
rect 10341 1703 10407 1719
rect 10341 1639 10342 1703
rect 10406 1639 10407 1703
rect 10341 1623 10407 1639
rect 10341 1559 10342 1623
rect 10406 1559 10407 1623
rect 10341 1543 10407 1559
rect 10341 1479 10342 1543
rect 10406 1479 10407 1543
rect 10341 1463 10407 1479
rect 10341 1399 10342 1463
rect 10406 1399 10407 1463
rect 10341 1383 10407 1399
rect 10341 1319 10342 1383
rect 10406 1319 10407 1383
rect 10341 1229 10407 1319
rect 10467 1165 10527 2195
rect 10587 1225 10647 2257
rect 10707 1165 10767 2195
rect 10827 1225 10887 2257
rect 10947 2103 11013 2257
rect 10947 2039 10948 2103
rect 11012 2039 11013 2103
rect 10947 2023 11013 2039
rect 10947 1959 10948 2023
rect 11012 1959 11013 2023
rect 10947 1943 11013 1959
rect 10947 1879 10948 1943
rect 11012 1879 11013 1943
rect 10947 1863 11013 1879
rect 10947 1799 10948 1863
rect 11012 1799 11013 1863
rect 10947 1783 11013 1799
rect 10947 1719 10948 1783
rect 11012 1719 11013 1783
rect 10947 1703 11013 1719
rect 10947 1639 10948 1703
rect 11012 1639 11013 1703
rect 10947 1623 11013 1639
rect 10947 1559 10948 1623
rect 11012 1559 11013 1623
rect 10947 1543 11013 1559
rect 10947 1479 10948 1543
rect 11012 1479 11013 1543
rect 10947 1463 11013 1479
rect 10947 1399 10948 1463
rect 11012 1399 11013 1463
rect 10947 1383 11013 1399
rect 10947 1319 10948 1383
rect 11012 1319 11013 1383
rect 10947 1229 11013 1319
rect 11073 2323 11571 2325
rect 11635 2325 11644 2346
rect 11780 2346 11862 2352
rect 11780 2325 11789 2346
rect 11635 2323 11789 2325
rect 11853 2325 11862 2346
rect 12514 2346 12596 2352
rect 12514 2325 12523 2346
rect 11853 2323 12351 2325
rect 11073 2259 11177 2323
rect 11241 2259 11257 2323
rect 11321 2259 11337 2323
rect 11401 2259 11417 2323
rect 11481 2259 11497 2323
rect 11561 2282 11571 2323
rect 11561 2259 11577 2282
rect 11641 2259 11783 2323
rect 11853 2282 11863 2323
rect 11847 2259 11863 2282
rect 11927 2259 11943 2323
rect 12007 2259 12023 2323
rect 12087 2259 12103 2323
rect 12167 2259 12183 2323
rect 12247 2259 12351 2323
rect 11073 2257 12351 2259
rect 11073 2103 11139 2257
rect 11073 2039 11074 2103
rect 11138 2039 11139 2103
rect 11073 2023 11139 2039
rect 11073 1959 11074 2023
rect 11138 1959 11139 2023
rect 11073 1943 11139 1959
rect 11073 1879 11074 1943
rect 11138 1879 11139 1943
rect 11073 1863 11139 1879
rect 11073 1799 11074 1863
rect 11138 1799 11139 1863
rect 11073 1783 11139 1799
rect 11073 1719 11074 1783
rect 11138 1719 11139 1783
rect 11073 1703 11139 1719
rect 11073 1639 11074 1703
rect 11138 1639 11139 1703
rect 11073 1623 11139 1639
rect 11073 1559 11074 1623
rect 11138 1559 11139 1623
rect 11073 1543 11139 1559
rect 11073 1479 11074 1543
rect 11138 1479 11139 1543
rect 11073 1463 11139 1479
rect 11073 1399 11074 1463
rect 11138 1399 11139 1463
rect 11073 1383 11139 1399
rect 11073 1319 11074 1383
rect 11138 1319 11139 1383
rect 11073 1229 11139 1319
rect 11199 1225 11259 2257
rect 11319 1165 11379 2195
rect 11439 1225 11499 2257
rect 11559 1165 11619 2195
rect 11679 2103 11745 2257
rect 11679 2039 11680 2103
rect 11744 2039 11745 2103
rect 11679 2023 11745 2039
rect 11679 1959 11680 2023
rect 11744 1959 11745 2023
rect 11679 1943 11745 1959
rect 11679 1879 11680 1943
rect 11744 1879 11745 1943
rect 11679 1863 11745 1879
rect 11679 1799 11680 1863
rect 11744 1799 11745 1863
rect 11679 1783 11745 1799
rect 11679 1719 11680 1783
rect 11744 1719 11745 1783
rect 11679 1703 11745 1719
rect 11679 1639 11680 1703
rect 11744 1639 11745 1703
rect 11679 1623 11745 1639
rect 11679 1559 11680 1623
rect 11744 1559 11745 1623
rect 11679 1543 11745 1559
rect 11679 1479 11680 1543
rect 11744 1479 11745 1543
rect 11679 1463 11745 1479
rect 11679 1399 11680 1463
rect 11744 1399 11745 1463
rect 11679 1383 11745 1399
rect 11679 1319 11680 1383
rect 11744 1319 11745 1383
rect 11679 1229 11745 1319
rect 11805 1165 11865 2195
rect 11925 1225 11985 2257
rect 12045 1165 12105 2195
rect 12165 1225 12225 2257
rect 12285 2103 12351 2257
rect 12285 2039 12286 2103
rect 12350 2039 12351 2103
rect 12285 2023 12351 2039
rect 12285 1959 12286 2023
rect 12350 1959 12351 2023
rect 12285 1943 12351 1959
rect 12285 1879 12286 1943
rect 12350 1879 12351 1943
rect 12285 1863 12351 1879
rect 12285 1799 12286 1863
rect 12350 1799 12351 1863
rect 12285 1783 12351 1799
rect 12285 1719 12286 1783
rect 12350 1719 12351 1783
rect 12285 1703 12351 1719
rect 12285 1639 12286 1703
rect 12350 1639 12351 1703
rect 12285 1623 12351 1639
rect 12285 1559 12286 1623
rect 12350 1559 12351 1623
rect 12285 1543 12351 1559
rect 12285 1479 12286 1543
rect 12350 1479 12351 1543
rect 12285 1463 12351 1479
rect 12285 1399 12286 1463
rect 12350 1399 12351 1463
rect 12285 1383 12351 1399
rect 12285 1319 12286 1383
rect 12350 1319 12351 1383
rect 12285 1229 12351 1319
rect 12413 2323 12523 2325
rect 12587 2325 12596 2346
rect 13236 2347 13362 2357
rect 12587 2323 13085 2325
rect 12413 2259 12517 2323
rect 12587 2282 12597 2323
rect 12581 2259 12597 2282
rect 12661 2259 12677 2323
rect 12741 2259 12757 2323
rect 12821 2259 12837 2323
rect 12901 2259 12917 2323
rect 12981 2259 13085 2323
rect 13236 2283 13267 2347
rect 13331 2283 13362 2347
rect 13236 2273 13362 2283
rect 13262 2272 13336 2273
rect 12413 2257 13085 2259
rect 12413 2103 12479 2257
rect 12413 2039 12414 2103
rect 12478 2039 12479 2103
rect 12413 2023 12479 2039
rect 12413 1959 12414 2023
rect 12478 1959 12479 2023
rect 12413 1943 12479 1959
rect 12413 1879 12414 1943
rect 12478 1879 12479 1943
rect 12413 1863 12479 1879
rect 12413 1799 12414 1863
rect 12478 1799 12479 1863
rect 12413 1783 12479 1799
rect 12413 1719 12414 1783
rect 12478 1719 12479 1783
rect 12413 1703 12479 1719
rect 12413 1639 12414 1703
rect 12478 1639 12479 1703
rect 12413 1623 12479 1639
rect 12413 1559 12414 1623
rect 12478 1559 12479 1623
rect 12413 1543 12479 1559
rect 12413 1479 12414 1543
rect 12478 1479 12479 1543
rect 12413 1463 12479 1479
rect 12413 1399 12414 1463
rect 12478 1399 12479 1463
rect 12413 1383 12479 1399
rect 12413 1319 12414 1383
rect 12478 1319 12479 1383
rect 12413 1229 12479 1319
rect 12539 1165 12599 2195
rect 12659 1225 12719 2257
rect 12779 1165 12839 2195
rect 12899 1225 12959 2257
rect 13019 2103 13085 2257
rect 13019 2039 13020 2103
rect 13084 2039 13085 2103
rect 13019 2023 13085 2039
rect 13019 1959 13020 2023
rect 13084 1959 13085 2023
rect 13146 2085 13271 2095
rect 13146 2021 13176 2085
rect 13240 2021 13271 2085
rect 13146 2011 13271 2021
rect 13019 1943 13085 1959
rect 13019 1879 13020 1943
rect 13084 1879 13085 1943
rect 13019 1863 13085 1879
rect 13019 1799 13020 1863
rect 13084 1799 13085 1863
rect 13019 1783 13085 1799
rect 13019 1719 13020 1783
rect 13084 1719 13085 1783
rect 13019 1703 13085 1719
rect 13019 1639 13020 1703
rect 13084 1639 13085 1703
rect 13019 1623 13085 1639
rect 13019 1559 13020 1623
rect 13084 1559 13085 1623
rect 13019 1543 13085 1559
rect 13019 1479 13020 1543
rect 13084 1479 13085 1543
rect 13019 1463 13085 1479
rect 13019 1399 13020 1463
rect 13084 1399 13085 1463
rect 13019 1383 13085 1399
rect 13019 1319 13020 1383
rect 13084 1319 13085 1383
rect 13019 1229 13085 1319
rect 694 1086 819 1096
rect 7403 1096 7433 1160
rect 7497 1096 7528 1160
rect 7791 1163 8463 1165
rect 7791 1099 7975 1163
rect 8039 1099 8055 1163
rect 8119 1099 8135 1163
rect 8199 1099 8215 1163
rect 8279 1099 8463 1163
rect 7791 1097 8463 1099
rect 8523 1163 11013 1165
rect 8523 1099 8707 1163
rect 8771 1099 8787 1163
rect 8851 1099 8867 1163
rect 8931 1099 8947 1163
rect 9011 1099 9313 1163
rect 9377 1099 9393 1163
rect 9457 1099 9473 1163
rect 9537 1099 9553 1163
rect 9617 1099 9919 1163
rect 9983 1099 9999 1163
rect 10063 1099 10079 1163
rect 10143 1099 10159 1163
rect 10223 1099 10525 1163
rect 10589 1099 10605 1163
rect 10669 1099 10685 1163
rect 10749 1099 10765 1163
rect 10829 1099 11013 1163
rect 8523 1097 11013 1099
rect 11073 1163 12351 1165
rect 11073 1099 11257 1163
rect 11321 1099 11337 1163
rect 11401 1099 11417 1163
rect 11481 1099 11497 1163
rect 11561 1099 11863 1163
rect 11927 1099 11943 1163
rect 12007 1099 12023 1163
rect 12087 1099 12103 1163
rect 12167 1099 12351 1163
rect 11073 1097 12351 1099
rect 12413 1163 13085 1165
rect 12413 1099 12597 1163
rect 12661 1099 12677 1163
rect 12741 1099 12757 1163
rect 12821 1099 12837 1163
rect 12901 1099 13085 1163
rect 12413 1097 13085 1099
rect 7403 1086 7528 1096
rect 5936 225 6061 235
rect 379 222 1051 224
rect 379 158 563 222
rect 627 158 643 222
rect 707 158 723 222
rect 787 158 803 222
rect 867 158 1051 222
rect 379 156 1051 158
rect 1113 222 2391 224
rect 1113 158 1297 222
rect 1361 158 1377 222
rect 1441 158 1457 222
rect 1521 158 1537 222
rect 1601 158 1903 222
rect 1967 158 1983 222
rect 2047 158 2063 222
rect 2127 158 2143 222
rect 2207 158 2391 222
rect 1113 156 2391 158
rect 2451 222 4941 224
rect 2451 158 2635 222
rect 2699 158 2715 222
rect 2779 158 2795 222
rect 2859 158 2875 222
rect 2939 158 3241 222
rect 3305 158 3321 222
rect 3385 158 3401 222
rect 3465 158 3481 222
rect 3545 158 3847 222
rect 3911 158 3927 222
rect 3991 158 4007 222
rect 4071 158 4087 222
rect 4151 158 4453 222
rect 4517 158 4533 222
rect 4597 158 4613 222
rect 4677 158 4693 222
rect 4757 158 4941 222
rect 2451 156 4941 158
rect 5001 222 5673 224
rect 5001 158 5185 222
rect 5249 158 5265 222
rect 5329 158 5345 222
rect 5409 158 5425 222
rect 5489 158 5673 222
rect 5001 156 5673 158
rect 5936 161 5967 225
rect 6031 161 6061 225
rect 12645 225 12770 235
rect 379 2 445 92
rect 379 -62 380 2
rect 444 -62 445 2
rect 379 -78 445 -62
rect 379 -142 380 -78
rect 444 -142 445 -78
rect 379 -158 445 -142
rect 379 -222 380 -158
rect 444 -222 445 -158
rect 379 -238 445 -222
rect 379 -302 380 -238
rect 444 -302 445 -238
rect 379 -318 445 -302
rect 379 -382 380 -318
rect 444 -382 445 -318
rect 379 -398 445 -382
rect 379 -462 380 -398
rect 444 -462 445 -398
rect 379 -478 445 -462
rect 379 -542 380 -478
rect 444 -542 445 -478
rect 379 -558 445 -542
rect 379 -622 380 -558
rect 444 -622 445 -558
rect 379 -638 445 -622
rect 193 -700 318 -690
rect 193 -764 224 -700
rect 288 -764 318 -700
rect 193 -774 318 -764
rect 379 -702 380 -638
rect 444 -702 445 -638
rect 379 -718 445 -702
rect 379 -782 380 -718
rect 444 -782 445 -718
rect 379 -936 445 -782
rect 505 -936 565 96
rect 625 -874 685 156
rect 745 -936 805 96
rect 865 -874 925 156
rect 985 2 1051 92
rect 985 -62 986 2
rect 1050 -62 1051 2
rect 985 -78 1051 -62
rect 985 -142 986 -78
rect 1050 -142 1051 -78
rect 985 -158 1051 -142
rect 985 -222 986 -158
rect 1050 -222 1051 -158
rect 985 -238 1051 -222
rect 985 -302 986 -238
rect 1050 -302 1051 -238
rect 985 -318 1051 -302
rect 985 -382 986 -318
rect 1050 -382 1051 -318
rect 985 -398 1051 -382
rect 985 -462 986 -398
rect 1050 -462 1051 -398
rect 985 -478 1051 -462
rect 985 -542 986 -478
rect 1050 -542 1051 -478
rect 985 -558 1051 -542
rect 985 -622 986 -558
rect 1050 -622 1051 -558
rect 985 -638 1051 -622
rect 985 -702 986 -638
rect 1050 -702 1051 -638
rect 985 -718 1051 -702
rect 985 -782 986 -718
rect 1050 -782 1051 -718
rect 985 -936 1051 -782
rect 379 -938 1051 -936
rect 128 -952 202 -951
rect 102 -962 228 -952
rect 102 -1026 133 -962
rect 197 -1026 228 -962
rect 379 -1002 483 -938
rect 547 -1002 563 -938
rect 627 -1002 643 -938
rect 707 -1002 723 -938
rect 787 -1002 803 -938
rect 867 -961 883 -938
rect 867 -1002 877 -961
rect 947 -1002 1051 -938
rect 379 -1004 877 -1002
rect 102 -1036 228 -1026
rect 868 -1025 877 -1004
rect 941 -1004 1051 -1002
rect 1113 2 1179 92
rect 1113 -62 1114 2
rect 1178 -62 1179 2
rect 1113 -78 1179 -62
rect 1113 -142 1114 -78
rect 1178 -142 1179 -78
rect 1113 -158 1179 -142
rect 1113 -222 1114 -158
rect 1178 -222 1179 -158
rect 1113 -238 1179 -222
rect 1113 -302 1114 -238
rect 1178 -302 1179 -238
rect 1113 -318 1179 -302
rect 1113 -382 1114 -318
rect 1178 -382 1179 -318
rect 1113 -398 1179 -382
rect 1113 -462 1114 -398
rect 1178 -462 1179 -398
rect 1113 -478 1179 -462
rect 1113 -542 1114 -478
rect 1178 -542 1179 -478
rect 1113 -558 1179 -542
rect 1113 -622 1114 -558
rect 1178 -622 1179 -558
rect 1113 -638 1179 -622
rect 1113 -702 1114 -638
rect 1178 -702 1179 -638
rect 1113 -718 1179 -702
rect 1113 -782 1114 -718
rect 1178 -782 1179 -718
rect 1113 -936 1179 -782
rect 1239 -936 1299 96
rect 1359 -874 1419 156
rect 1479 -936 1539 96
rect 1599 -874 1659 156
rect 1719 2 1785 92
rect 1719 -62 1720 2
rect 1784 -62 1785 2
rect 1719 -78 1785 -62
rect 1719 -142 1720 -78
rect 1784 -142 1785 -78
rect 1719 -158 1785 -142
rect 1719 -222 1720 -158
rect 1784 -222 1785 -158
rect 1719 -238 1785 -222
rect 1719 -302 1720 -238
rect 1784 -302 1785 -238
rect 1719 -318 1785 -302
rect 1719 -382 1720 -318
rect 1784 -382 1785 -318
rect 1719 -398 1785 -382
rect 1719 -462 1720 -398
rect 1784 -462 1785 -398
rect 1719 -478 1785 -462
rect 1719 -542 1720 -478
rect 1784 -542 1785 -478
rect 1719 -558 1785 -542
rect 1719 -622 1720 -558
rect 1784 -622 1785 -558
rect 1719 -638 1785 -622
rect 1719 -702 1720 -638
rect 1784 -702 1785 -638
rect 1719 -718 1785 -702
rect 1719 -782 1720 -718
rect 1784 -782 1785 -718
rect 1719 -936 1785 -782
rect 1845 -874 1905 156
rect 1965 -936 2025 96
rect 2085 -874 2145 156
rect 2205 -936 2265 96
rect 2325 2 2391 92
rect 2325 -62 2326 2
rect 2390 -62 2391 2
rect 2325 -78 2391 -62
rect 2325 -142 2326 -78
rect 2390 -142 2391 -78
rect 2325 -158 2391 -142
rect 2325 -222 2326 -158
rect 2390 -222 2391 -158
rect 2325 -238 2391 -222
rect 2325 -302 2326 -238
rect 2390 -302 2391 -238
rect 2325 -318 2391 -302
rect 2325 -382 2326 -318
rect 2390 -382 2391 -318
rect 2325 -398 2391 -382
rect 2325 -462 2326 -398
rect 2390 -462 2391 -398
rect 2325 -478 2391 -462
rect 2325 -542 2326 -478
rect 2390 -542 2391 -478
rect 2325 -558 2391 -542
rect 2325 -622 2326 -558
rect 2390 -622 2391 -558
rect 2325 -638 2391 -622
rect 2325 -702 2326 -638
rect 2390 -702 2391 -638
rect 2325 -718 2391 -702
rect 2325 -782 2326 -718
rect 2390 -782 2391 -718
rect 2325 -936 2391 -782
rect 1113 -938 2391 -936
rect 1113 -1002 1217 -938
rect 1281 -1002 1297 -938
rect 1361 -1002 1377 -938
rect 1441 -1002 1457 -938
rect 1521 -1002 1537 -938
rect 1601 -961 1617 -938
rect 1601 -1002 1611 -961
rect 1681 -1002 1823 -938
rect 1887 -961 1903 -938
rect 1893 -1002 1903 -961
rect 1967 -1002 1983 -938
rect 2047 -1002 2063 -938
rect 2127 -1002 2143 -938
rect 2207 -1002 2223 -938
rect 2287 -1002 2391 -938
rect 1113 -1004 1611 -1002
rect 941 -1025 950 -1004
rect 868 -1031 950 -1025
rect 1602 -1025 1611 -1004
rect 1675 -1004 1829 -1002
rect 1675 -1025 1684 -1004
rect 1602 -1031 1684 -1025
rect 1820 -1025 1829 -1004
rect 1893 -1004 2391 -1002
rect 2451 2 2517 92
rect 2451 -62 2452 2
rect 2516 -62 2517 2
rect 2451 -78 2517 -62
rect 2451 -142 2452 -78
rect 2516 -142 2517 -78
rect 2451 -158 2517 -142
rect 2451 -222 2452 -158
rect 2516 -222 2517 -158
rect 2451 -238 2517 -222
rect 2451 -302 2452 -238
rect 2516 -302 2517 -238
rect 2451 -318 2517 -302
rect 2451 -382 2452 -318
rect 2516 -382 2517 -318
rect 2451 -398 2517 -382
rect 2451 -462 2452 -398
rect 2516 -462 2517 -398
rect 2451 -478 2517 -462
rect 2451 -542 2452 -478
rect 2516 -542 2517 -478
rect 2451 -558 2517 -542
rect 2451 -622 2452 -558
rect 2516 -622 2517 -558
rect 2451 -638 2517 -622
rect 2451 -702 2452 -638
rect 2516 -702 2517 -638
rect 2451 -718 2517 -702
rect 2451 -782 2452 -718
rect 2516 -782 2517 -718
rect 2451 -936 2517 -782
rect 2577 -936 2637 96
rect 2697 -874 2757 156
rect 2817 -936 2877 96
rect 2937 -874 2997 156
rect 3057 2 3123 92
rect 3057 -62 3058 2
rect 3122 -62 3123 2
rect 3057 -78 3123 -62
rect 3057 -142 3058 -78
rect 3122 -142 3123 -78
rect 3057 -158 3123 -142
rect 3057 -222 3058 -158
rect 3122 -222 3123 -158
rect 3057 -238 3123 -222
rect 3057 -302 3058 -238
rect 3122 -302 3123 -238
rect 3057 -318 3123 -302
rect 3057 -382 3058 -318
rect 3122 -382 3123 -318
rect 3057 -398 3123 -382
rect 3057 -462 3058 -398
rect 3122 -462 3123 -398
rect 3057 -478 3123 -462
rect 3057 -542 3058 -478
rect 3122 -542 3123 -478
rect 3057 -558 3123 -542
rect 3057 -622 3058 -558
rect 3122 -622 3123 -558
rect 3057 -638 3123 -622
rect 3057 -702 3058 -638
rect 3122 -702 3123 -638
rect 3057 -718 3123 -702
rect 3057 -782 3058 -718
rect 3122 -782 3123 -718
rect 3057 -936 3123 -782
rect 3183 -874 3243 156
rect 3303 -936 3363 96
rect 3423 -874 3483 156
rect 3543 -936 3603 96
rect 3663 2 3729 92
rect 3663 -62 3664 2
rect 3728 -62 3729 2
rect 3663 -78 3729 -62
rect 3663 -142 3664 -78
rect 3728 -142 3729 -78
rect 3663 -158 3729 -142
rect 3663 -222 3664 -158
rect 3728 -222 3729 -158
rect 3663 -238 3729 -222
rect 3663 -302 3664 -238
rect 3728 -302 3729 -238
rect 3663 -318 3729 -302
rect 3663 -382 3664 -318
rect 3728 -382 3729 -318
rect 3663 -398 3729 -382
rect 3663 -462 3664 -398
rect 3728 -462 3729 -398
rect 3663 -478 3729 -462
rect 3663 -542 3664 -478
rect 3728 -542 3729 -478
rect 3663 -558 3729 -542
rect 3663 -622 3664 -558
rect 3728 -622 3729 -558
rect 3663 -638 3729 -622
rect 3663 -702 3664 -638
rect 3728 -702 3729 -638
rect 3663 -718 3729 -702
rect 3663 -782 3664 -718
rect 3728 -782 3729 -718
rect 3663 -936 3729 -782
rect 3789 -936 3849 96
rect 3909 -874 3969 156
rect 4029 -936 4089 96
rect 4149 -874 4209 156
rect 4269 2 4335 92
rect 4269 -62 4270 2
rect 4334 -62 4335 2
rect 4269 -78 4335 -62
rect 4269 -142 4270 -78
rect 4334 -142 4335 -78
rect 4269 -158 4335 -142
rect 4269 -222 4270 -158
rect 4334 -222 4335 -158
rect 4269 -238 4335 -222
rect 4269 -302 4270 -238
rect 4334 -302 4335 -238
rect 4269 -318 4335 -302
rect 4269 -382 4270 -318
rect 4334 -382 4335 -318
rect 4269 -398 4335 -382
rect 4269 -462 4270 -398
rect 4334 -462 4335 -398
rect 4269 -478 4335 -462
rect 4269 -542 4270 -478
rect 4334 -542 4335 -478
rect 4269 -558 4335 -542
rect 4269 -622 4270 -558
rect 4334 -622 4335 -558
rect 4269 -638 4335 -622
rect 4269 -702 4270 -638
rect 4334 -702 4335 -638
rect 4269 -718 4335 -702
rect 4269 -782 4270 -718
rect 4334 -782 4335 -718
rect 4269 -936 4335 -782
rect 4395 -874 4455 156
rect 4515 -936 4575 96
rect 4635 -874 4695 156
rect 4755 -936 4815 96
rect 4875 2 4941 92
rect 4875 -62 4876 2
rect 4940 -62 4941 2
rect 4875 -78 4941 -62
rect 4875 -142 4876 -78
rect 4940 -142 4941 -78
rect 4875 -158 4941 -142
rect 4875 -222 4876 -158
rect 4940 -222 4941 -158
rect 4875 -238 4941 -222
rect 4875 -302 4876 -238
rect 4940 -302 4941 -238
rect 4875 -318 4941 -302
rect 4875 -382 4876 -318
rect 4940 -382 4941 -318
rect 4875 -398 4941 -382
rect 4875 -462 4876 -398
rect 4940 -462 4941 -398
rect 4875 -478 4941 -462
rect 4875 -542 4876 -478
rect 4940 -542 4941 -478
rect 4875 -558 4941 -542
rect 4875 -622 4876 -558
rect 4940 -622 4941 -558
rect 4875 -638 4941 -622
rect 4875 -702 4876 -638
rect 4940 -702 4941 -638
rect 4875 -718 4941 -702
rect 4875 -782 4876 -718
rect 4940 -782 4941 -718
rect 4875 -936 4941 -782
rect 2451 -938 4941 -936
rect 2451 -1002 2555 -938
rect 2619 -1002 2635 -938
rect 2699 -1002 2715 -938
rect 2779 -1002 2795 -938
rect 2859 -1002 2875 -938
rect 2939 -961 2955 -938
rect 2939 -1002 2949 -961
rect 3019 -1002 3161 -938
rect 3225 -961 3241 -938
rect 3231 -1002 3241 -961
rect 3305 -1002 3321 -938
rect 3385 -1002 3401 -938
rect 3465 -1002 3481 -938
rect 3545 -1002 3561 -938
rect 3625 -1002 3767 -938
rect 3831 -1002 3847 -938
rect 3911 -1002 3927 -938
rect 3991 -1002 4007 -938
rect 4071 -1002 4087 -938
rect 4151 -961 4167 -938
rect 4151 -1002 4161 -961
rect 4231 -1002 4373 -938
rect 4437 -961 4453 -938
rect 4443 -1002 4453 -961
rect 4517 -1002 4533 -938
rect 4597 -1002 4613 -938
rect 4677 -1002 4693 -938
rect 4757 -1002 4773 -938
rect 4837 -1002 4941 -938
rect 2451 -1004 2949 -1002
rect 1893 -1025 1902 -1004
rect 1820 -1031 1902 -1025
rect 2940 -1025 2949 -1004
rect 3013 -1004 3167 -1002
rect 3013 -1025 3022 -1004
rect 2940 -1031 3022 -1025
rect 3158 -1025 3167 -1004
rect 3231 -1004 4161 -1002
rect 3231 -1025 3240 -1004
rect 3158 -1031 3240 -1025
rect 4152 -1025 4161 -1004
rect 4225 -1004 4379 -1002
rect 4225 -1025 4234 -1004
rect 4152 -1031 4234 -1025
rect 4370 -1025 4379 -1004
rect 4443 -1004 4941 -1002
rect 5001 2 5067 92
rect 5001 -62 5002 2
rect 5066 -62 5067 2
rect 5001 -78 5067 -62
rect 5001 -142 5002 -78
rect 5066 -142 5067 -78
rect 5001 -158 5067 -142
rect 5001 -222 5002 -158
rect 5066 -222 5067 -158
rect 5001 -238 5067 -222
rect 5001 -302 5002 -238
rect 5066 -302 5067 -238
rect 5001 -318 5067 -302
rect 5001 -382 5002 -318
rect 5066 -382 5067 -318
rect 5001 -398 5067 -382
rect 5001 -462 5002 -398
rect 5066 -462 5067 -398
rect 5001 -478 5067 -462
rect 5001 -542 5002 -478
rect 5066 -542 5067 -478
rect 5001 -558 5067 -542
rect 5001 -622 5002 -558
rect 5066 -622 5067 -558
rect 5001 -638 5067 -622
rect 5001 -702 5002 -638
rect 5066 -702 5067 -638
rect 5001 -718 5067 -702
rect 5001 -782 5002 -718
rect 5066 -782 5067 -718
rect 5001 -936 5067 -782
rect 5127 -874 5187 156
rect 5247 -936 5307 96
rect 5367 -874 5427 156
rect 5936 151 6061 161
rect 7088 222 7760 224
rect 7088 158 7272 222
rect 7336 158 7352 222
rect 7416 158 7432 222
rect 7496 158 7512 222
rect 7576 158 7760 222
rect 7088 156 7760 158
rect 7822 222 9100 224
rect 7822 158 8006 222
rect 8070 158 8086 222
rect 8150 158 8166 222
rect 8230 158 8246 222
rect 8310 158 8612 222
rect 8676 158 8692 222
rect 8756 158 8772 222
rect 8836 158 8852 222
rect 8916 158 9100 222
rect 7822 156 9100 158
rect 9160 222 11650 224
rect 9160 158 9344 222
rect 9408 158 9424 222
rect 9488 158 9504 222
rect 9568 158 9584 222
rect 9648 158 9950 222
rect 10014 158 10030 222
rect 10094 158 10110 222
rect 10174 158 10190 222
rect 10254 158 10556 222
rect 10620 158 10636 222
rect 10700 158 10716 222
rect 10780 158 10796 222
rect 10860 158 11162 222
rect 11226 158 11242 222
rect 11306 158 11322 222
rect 11386 158 11402 222
rect 11466 158 11650 222
rect 9160 156 11650 158
rect 11710 222 12382 224
rect 11710 158 11894 222
rect 11958 158 11974 222
rect 12038 158 12054 222
rect 12118 158 12134 222
rect 12198 158 12382 222
rect 11710 156 12382 158
rect 12645 161 12676 225
rect 12740 161 12770 225
rect 5487 -936 5547 96
rect 5607 2 5673 92
rect 5607 -62 5608 2
rect 5672 -62 5673 2
rect 5607 -78 5673 -62
rect 5607 -142 5608 -78
rect 5672 -142 5673 -78
rect 5607 -158 5673 -142
rect 5607 -222 5608 -158
rect 5672 -222 5673 -158
rect 5607 -238 5673 -222
rect 5607 -302 5608 -238
rect 5672 -302 5673 -238
rect 5607 -318 5673 -302
rect 5607 -382 5608 -318
rect 5672 -382 5673 -318
rect 5607 -398 5673 -382
rect 5607 -462 5608 -398
rect 5672 -462 5673 -398
rect 5607 -478 5673 -462
rect 5607 -542 5608 -478
rect 5672 -542 5673 -478
rect 5607 -558 5673 -542
rect 5607 -622 5608 -558
rect 5672 -622 5673 -558
rect 5607 -638 5673 -622
rect 5607 -702 5608 -638
rect 5672 -702 5673 -638
rect 7088 2 7154 92
rect 7088 -62 7089 2
rect 7153 -62 7154 2
rect 7088 -78 7154 -62
rect 7088 -142 7089 -78
rect 7153 -142 7154 -78
rect 7088 -158 7154 -142
rect 7088 -222 7089 -158
rect 7153 -222 7154 -158
rect 7088 -238 7154 -222
rect 7088 -302 7089 -238
rect 7153 -302 7154 -238
rect 7088 -318 7154 -302
rect 7088 -382 7089 -318
rect 7153 -382 7154 -318
rect 7088 -398 7154 -382
rect 7088 -462 7089 -398
rect 7153 -462 7154 -398
rect 7088 -478 7154 -462
rect 7088 -542 7089 -478
rect 7153 -542 7154 -478
rect 7088 -558 7154 -542
rect 7088 -622 7089 -558
rect 7153 -622 7154 -558
rect 7088 -638 7154 -622
rect 5607 -718 5673 -702
rect 5607 -782 5608 -718
rect 5672 -782 5673 -718
rect 6902 -700 7027 -690
rect 6902 -764 6933 -700
rect 6997 -764 7027 -700
rect 6902 -774 7027 -764
rect 7088 -702 7089 -638
rect 7153 -702 7154 -638
rect 7088 -718 7154 -702
rect 5607 -936 5673 -782
rect 5001 -938 5673 -936
rect 5001 -1002 5105 -938
rect 5169 -961 5185 -938
rect 5175 -1002 5185 -961
rect 5249 -1002 5265 -938
rect 5329 -1002 5345 -938
rect 5409 -1002 5425 -938
rect 5489 -1002 5505 -938
rect 5569 -1002 5673 -938
rect 7088 -782 7089 -718
rect 7153 -782 7154 -718
rect 7088 -936 7154 -782
rect 7214 -936 7274 96
rect 7334 -874 7394 156
rect 7454 -936 7514 96
rect 7574 -874 7634 156
rect 7694 2 7760 92
rect 7694 -62 7695 2
rect 7759 -62 7760 2
rect 7694 -78 7760 -62
rect 7694 -142 7695 -78
rect 7759 -142 7760 -78
rect 7694 -158 7760 -142
rect 7694 -222 7695 -158
rect 7759 -222 7760 -158
rect 7694 -238 7760 -222
rect 7694 -302 7695 -238
rect 7759 -302 7760 -238
rect 7694 -318 7760 -302
rect 7694 -382 7695 -318
rect 7759 -382 7760 -318
rect 7694 -398 7760 -382
rect 7694 -462 7695 -398
rect 7759 -462 7760 -398
rect 7694 -478 7760 -462
rect 7694 -542 7695 -478
rect 7759 -542 7760 -478
rect 7694 -558 7760 -542
rect 7694 -622 7695 -558
rect 7759 -622 7760 -558
rect 7694 -638 7760 -622
rect 7694 -702 7695 -638
rect 7759 -702 7760 -638
rect 7694 -718 7760 -702
rect 7694 -782 7695 -718
rect 7759 -782 7760 -718
rect 7694 -936 7760 -782
rect 7088 -938 7760 -936
rect 6837 -952 6911 -951
rect 5001 -1004 5111 -1002
rect 4443 -1025 4452 -1004
rect 4370 -1031 4452 -1025
rect 5102 -1025 5111 -1004
rect 5175 -1004 5673 -1002
rect 6811 -962 6937 -952
rect 5175 -1025 5184 -1004
rect 5102 -1031 5184 -1025
rect 6811 -1026 6842 -962
rect 6906 -1026 6937 -962
rect 7088 -1002 7192 -938
rect 7256 -1002 7272 -938
rect 7336 -1002 7352 -938
rect 7416 -1002 7432 -938
rect 7496 -1002 7512 -938
rect 7576 -961 7592 -938
rect 7576 -1002 7586 -961
rect 7656 -1002 7760 -938
rect 7088 -1004 7586 -1002
rect 6811 -1036 6937 -1026
rect 7577 -1025 7586 -1004
rect 7650 -1004 7760 -1002
rect 7822 2 7888 92
rect 7822 -62 7823 2
rect 7887 -62 7888 2
rect 7822 -78 7888 -62
rect 7822 -142 7823 -78
rect 7887 -142 7888 -78
rect 7822 -158 7888 -142
rect 7822 -222 7823 -158
rect 7887 -222 7888 -158
rect 7822 -238 7888 -222
rect 7822 -302 7823 -238
rect 7887 -302 7888 -238
rect 7822 -318 7888 -302
rect 7822 -382 7823 -318
rect 7887 -382 7888 -318
rect 7822 -398 7888 -382
rect 7822 -462 7823 -398
rect 7887 -462 7888 -398
rect 7822 -478 7888 -462
rect 7822 -542 7823 -478
rect 7887 -542 7888 -478
rect 7822 -558 7888 -542
rect 7822 -622 7823 -558
rect 7887 -622 7888 -558
rect 7822 -638 7888 -622
rect 7822 -702 7823 -638
rect 7887 -702 7888 -638
rect 7822 -718 7888 -702
rect 7822 -782 7823 -718
rect 7887 -782 7888 -718
rect 7822 -936 7888 -782
rect 7948 -936 8008 96
rect 8068 -874 8128 156
rect 8188 -936 8248 96
rect 8308 -874 8368 156
rect 8428 2 8494 92
rect 8428 -62 8429 2
rect 8493 -62 8494 2
rect 8428 -78 8494 -62
rect 8428 -142 8429 -78
rect 8493 -142 8494 -78
rect 8428 -158 8494 -142
rect 8428 -222 8429 -158
rect 8493 -222 8494 -158
rect 8428 -238 8494 -222
rect 8428 -302 8429 -238
rect 8493 -302 8494 -238
rect 8428 -318 8494 -302
rect 8428 -382 8429 -318
rect 8493 -382 8494 -318
rect 8428 -398 8494 -382
rect 8428 -462 8429 -398
rect 8493 -462 8494 -398
rect 8428 -478 8494 -462
rect 8428 -542 8429 -478
rect 8493 -542 8494 -478
rect 8428 -558 8494 -542
rect 8428 -622 8429 -558
rect 8493 -622 8494 -558
rect 8428 -638 8494 -622
rect 8428 -702 8429 -638
rect 8493 -702 8494 -638
rect 8428 -718 8494 -702
rect 8428 -782 8429 -718
rect 8493 -782 8494 -718
rect 8428 -936 8494 -782
rect 8554 -874 8614 156
rect 8674 -936 8734 96
rect 8794 -874 8854 156
rect 8914 -936 8974 96
rect 9034 2 9100 92
rect 9034 -62 9035 2
rect 9099 -62 9100 2
rect 9034 -78 9100 -62
rect 9034 -142 9035 -78
rect 9099 -142 9100 -78
rect 9034 -158 9100 -142
rect 9034 -222 9035 -158
rect 9099 -222 9100 -158
rect 9034 -238 9100 -222
rect 9034 -302 9035 -238
rect 9099 -302 9100 -238
rect 9034 -318 9100 -302
rect 9034 -382 9035 -318
rect 9099 -382 9100 -318
rect 9034 -398 9100 -382
rect 9034 -462 9035 -398
rect 9099 -462 9100 -398
rect 9034 -478 9100 -462
rect 9034 -542 9035 -478
rect 9099 -542 9100 -478
rect 9034 -558 9100 -542
rect 9034 -622 9035 -558
rect 9099 -622 9100 -558
rect 9034 -638 9100 -622
rect 9034 -702 9035 -638
rect 9099 -702 9100 -638
rect 9034 -718 9100 -702
rect 9034 -782 9035 -718
rect 9099 -782 9100 -718
rect 9034 -936 9100 -782
rect 7822 -938 9100 -936
rect 7822 -1002 7926 -938
rect 7990 -1002 8006 -938
rect 8070 -1002 8086 -938
rect 8150 -1002 8166 -938
rect 8230 -1002 8246 -938
rect 8310 -961 8326 -938
rect 8310 -1002 8320 -961
rect 8390 -1002 8532 -938
rect 8596 -961 8612 -938
rect 8602 -1002 8612 -961
rect 8676 -1002 8692 -938
rect 8756 -1002 8772 -938
rect 8836 -1002 8852 -938
rect 8916 -1002 8932 -938
rect 8996 -1002 9100 -938
rect 7822 -1004 8320 -1002
rect 7650 -1025 7659 -1004
rect 7577 -1031 7659 -1025
rect 8311 -1025 8320 -1004
rect 8384 -1004 8538 -1002
rect 8384 -1025 8393 -1004
rect 8311 -1031 8393 -1025
rect 8529 -1025 8538 -1004
rect 8602 -1004 9100 -1002
rect 9160 2 9226 92
rect 9160 -62 9161 2
rect 9225 -62 9226 2
rect 9160 -78 9226 -62
rect 9160 -142 9161 -78
rect 9225 -142 9226 -78
rect 9160 -158 9226 -142
rect 9160 -222 9161 -158
rect 9225 -222 9226 -158
rect 9160 -238 9226 -222
rect 9160 -302 9161 -238
rect 9225 -302 9226 -238
rect 9160 -318 9226 -302
rect 9160 -382 9161 -318
rect 9225 -382 9226 -318
rect 9160 -398 9226 -382
rect 9160 -462 9161 -398
rect 9225 -462 9226 -398
rect 9160 -478 9226 -462
rect 9160 -542 9161 -478
rect 9225 -542 9226 -478
rect 9160 -558 9226 -542
rect 9160 -622 9161 -558
rect 9225 -622 9226 -558
rect 9160 -638 9226 -622
rect 9160 -702 9161 -638
rect 9225 -702 9226 -638
rect 9160 -718 9226 -702
rect 9160 -782 9161 -718
rect 9225 -782 9226 -718
rect 9160 -936 9226 -782
rect 9286 -936 9346 96
rect 9406 -874 9466 156
rect 9526 -936 9586 96
rect 9646 -874 9706 156
rect 9766 2 9832 92
rect 9766 -62 9767 2
rect 9831 -62 9832 2
rect 9766 -78 9832 -62
rect 9766 -142 9767 -78
rect 9831 -142 9832 -78
rect 9766 -158 9832 -142
rect 9766 -222 9767 -158
rect 9831 -222 9832 -158
rect 9766 -238 9832 -222
rect 9766 -302 9767 -238
rect 9831 -302 9832 -238
rect 9766 -318 9832 -302
rect 9766 -382 9767 -318
rect 9831 -382 9832 -318
rect 9766 -398 9832 -382
rect 9766 -462 9767 -398
rect 9831 -462 9832 -398
rect 9766 -478 9832 -462
rect 9766 -542 9767 -478
rect 9831 -542 9832 -478
rect 9766 -558 9832 -542
rect 9766 -622 9767 -558
rect 9831 -622 9832 -558
rect 9766 -638 9832 -622
rect 9766 -702 9767 -638
rect 9831 -702 9832 -638
rect 9766 -718 9832 -702
rect 9766 -782 9767 -718
rect 9831 -782 9832 -718
rect 9766 -936 9832 -782
rect 9892 -874 9952 156
rect 10012 -936 10072 96
rect 10132 -874 10192 156
rect 10252 -936 10312 96
rect 10372 2 10438 92
rect 10372 -62 10373 2
rect 10437 -62 10438 2
rect 10372 -78 10438 -62
rect 10372 -142 10373 -78
rect 10437 -142 10438 -78
rect 10372 -158 10438 -142
rect 10372 -222 10373 -158
rect 10437 -222 10438 -158
rect 10372 -238 10438 -222
rect 10372 -302 10373 -238
rect 10437 -302 10438 -238
rect 10372 -318 10438 -302
rect 10372 -382 10373 -318
rect 10437 -382 10438 -318
rect 10372 -398 10438 -382
rect 10372 -462 10373 -398
rect 10437 -462 10438 -398
rect 10372 -478 10438 -462
rect 10372 -542 10373 -478
rect 10437 -542 10438 -478
rect 10372 -558 10438 -542
rect 10372 -622 10373 -558
rect 10437 -622 10438 -558
rect 10372 -638 10438 -622
rect 10372 -702 10373 -638
rect 10437 -702 10438 -638
rect 10372 -718 10438 -702
rect 10372 -782 10373 -718
rect 10437 -782 10438 -718
rect 10372 -936 10438 -782
rect 10498 -936 10558 96
rect 10618 -874 10678 156
rect 10738 -936 10798 96
rect 10858 -874 10918 156
rect 10978 2 11044 92
rect 10978 -62 10979 2
rect 11043 -62 11044 2
rect 10978 -78 11044 -62
rect 10978 -142 10979 -78
rect 11043 -142 11044 -78
rect 10978 -158 11044 -142
rect 10978 -222 10979 -158
rect 11043 -222 11044 -158
rect 10978 -238 11044 -222
rect 10978 -302 10979 -238
rect 11043 -302 11044 -238
rect 10978 -318 11044 -302
rect 10978 -382 10979 -318
rect 11043 -382 11044 -318
rect 10978 -398 11044 -382
rect 10978 -462 10979 -398
rect 11043 -462 11044 -398
rect 10978 -478 11044 -462
rect 10978 -542 10979 -478
rect 11043 -542 11044 -478
rect 10978 -558 11044 -542
rect 10978 -622 10979 -558
rect 11043 -622 11044 -558
rect 10978 -638 11044 -622
rect 10978 -702 10979 -638
rect 11043 -702 11044 -638
rect 10978 -718 11044 -702
rect 10978 -782 10979 -718
rect 11043 -782 11044 -718
rect 10978 -936 11044 -782
rect 11104 -874 11164 156
rect 11224 -936 11284 96
rect 11344 -874 11404 156
rect 11464 -936 11524 96
rect 11584 2 11650 92
rect 11584 -62 11585 2
rect 11649 -62 11650 2
rect 11584 -78 11650 -62
rect 11584 -142 11585 -78
rect 11649 -142 11650 -78
rect 11584 -158 11650 -142
rect 11584 -222 11585 -158
rect 11649 -222 11650 -158
rect 11584 -238 11650 -222
rect 11584 -302 11585 -238
rect 11649 -302 11650 -238
rect 11584 -318 11650 -302
rect 11584 -382 11585 -318
rect 11649 -382 11650 -318
rect 11584 -398 11650 -382
rect 11584 -462 11585 -398
rect 11649 -462 11650 -398
rect 11584 -478 11650 -462
rect 11584 -542 11585 -478
rect 11649 -542 11650 -478
rect 11584 -558 11650 -542
rect 11584 -622 11585 -558
rect 11649 -622 11650 -558
rect 11584 -638 11650 -622
rect 11584 -702 11585 -638
rect 11649 -702 11650 -638
rect 11584 -718 11650 -702
rect 11584 -782 11585 -718
rect 11649 -782 11650 -718
rect 11584 -936 11650 -782
rect 9160 -938 11650 -936
rect 9160 -1002 9264 -938
rect 9328 -1002 9344 -938
rect 9408 -1002 9424 -938
rect 9488 -1002 9504 -938
rect 9568 -1002 9584 -938
rect 9648 -961 9664 -938
rect 9648 -1002 9658 -961
rect 9728 -1002 9870 -938
rect 9934 -961 9950 -938
rect 9940 -1002 9950 -961
rect 10014 -1002 10030 -938
rect 10094 -1002 10110 -938
rect 10174 -1002 10190 -938
rect 10254 -1002 10270 -938
rect 10334 -1002 10476 -938
rect 10540 -1002 10556 -938
rect 10620 -1002 10636 -938
rect 10700 -1002 10716 -938
rect 10780 -1002 10796 -938
rect 10860 -961 10876 -938
rect 10860 -1002 10870 -961
rect 10940 -1002 11082 -938
rect 11146 -961 11162 -938
rect 11152 -1002 11162 -961
rect 11226 -1002 11242 -938
rect 11306 -1002 11322 -938
rect 11386 -1002 11402 -938
rect 11466 -1002 11482 -938
rect 11546 -1002 11650 -938
rect 9160 -1004 9658 -1002
rect 8602 -1025 8611 -1004
rect 8529 -1031 8611 -1025
rect 9649 -1025 9658 -1004
rect 9722 -1004 9876 -1002
rect 9722 -1025 9731 -1004
rect 9649 -1031 9731 -1025
rect 9867 -1025 9876 -1004
rect 9940 -1004 10870 -1002
rect 9940 -1025 9949 -1004
rect 9867 -1031 9949 -1025
rect 10861 -1025 10870 -1004
rect 10934 -1004 11088 -1002
rect 10934 -1025 10943 -1004
rect 10861 -1031 10943 -1025
rect 11079 -1025 11088 -1004
rect 11152 -1004 11650 -1002
rect 11710 2 11776 92
rect 11710 -62 11711 2
rect 11775 -62 11776 2
rect 11710 -78 11776 -62
rect 11710 -142 11711 -78
rect 11775 -142 11776 -78
rect 11710 -158 11776 -142
rect 11710 -222 11711 -158
rect 11775 -222 11776 -158
rect 11710 -238 11776 -222
rect 11710 -302 11711 -238
rect 11775 -302 11776 -238
rect 11710 -318 11776 -302
rect 11710 -382 11711 -318
rect 11775 -382 11776 -318
rect 11710 -398 11776 -382
rect 11710 -462 11711 -398
rect 11775 -462 11776 -398
rect 11710 -478 11776 -462
rect 11710 -542 11711 -478
rect 11775 -542 11776 -478
rect 11710 -558 11776 -542
rect 11710 -622 11711 -558
rect 11775 -622 11776 -558
rect 11710 -638 11776 -622
rect 11710 -702 11711 -638
rect 11775 -702 11776 -638
rect 11710 -718 11776 -702
rect 11710 -782 11711 -718
rect 11775 -782 11776 -718
rect 11710 -936 11776 -782
rect 11836 -874 11896 156
rect 11956 -936 12016 96
rect 12076 -874 12136 156
rect 12645 151 12770 161
rect 12196 -936 12256 96
rect 12316 2 12382 92
rect 12316 -62 12317 2
rect 12381 -62 12382 2
rect 12316 -78 12382 -62
rect 12316 -142 12317 -78
rect 12381 -142 12382 -78
rect 12316 -158 12382 -142
rect 12316 -222 12317 -158
rect 12381 -222 12382 -158
rect 12316 -238 12382 -222
rect 12316 -302 12317 -238
rect 12381 -302 12382 -238
rect 12316 -318 12382 -302
rect 12316 -382 12317 -318
rect 12381 -382 12382 -318
rect 12316 -398 12382 -382
rect 12316 -462 12317 -398
rect 12381 -462 12382 -398
rect 12316 -478 12382 -462
rect 12316 -542 12317 -478
rect 12381 -542 12382 -478
rect 12316 -558 12382 -542
rect 12316 -622 12317 -558
rect 12381 -622 12382 -558
rect 12316 -638 12382 -622
rect 12316 -702 12317 -638
rect 12381 -702 12382 -638
rect 12316 -718 12382 -702
rect 12316 -782 12317 -718
rect 12381 -782 12382 -718
rect 12316 -936 12382 -782
rect 11710 -938 12382 -936
rect 11710 -1002 11814 -938
rect 11878 -961 11894 -938
rect 11884 -1002 11894 -961
rect 11958 -1002 11974 -938
rect 12038 -1002 12054 -938
rect 12118 -1002 12134 -938
rect 12198 -1002 12214 -938
rect 12278 -1002 12382 -938
rect 11710 -1004 11820 -1002
rect 11152 -1025 11161 -1004
rect 11079 -1031 11161 -1025
rect 11811 -1025 11820 -1004
rect 11884 -1004 12382 -1002
rect 11884 -1025 11893 -1004
rect 11811 -1031 11893 -1025
rect 102 -1165 228 -1155
rect 102 -1229 133 -1165
rect 197 -1229 228 -1165
rect 861 -1163 944 -1158
rect 861 -1184 871 -1163
rect 102 -1239 228 -1229
rect 378 -1186 871 -1184
rect 935 -1184 944 -1163
rect 1090 -1163 1173 -1158
rect 1090 -1184 1099 -1163
rect 935 -1186 1099 -1184
rect 1163 -1184 1173 -1163
rect 2073 -1163 2156 -1158
rect 2073 -1184 2083 -1163
rect 1163 -1186 2083 -1184
rect 2147 -1184 2156 -1163
rect 2302 -1163 2385 -1158
rect 2302 -1184 2311 -1163
rect 2147 -1186 2311 -1184
rect 2375 -1184 2385 -1163
rect 3285 -1163 3368 -1158
rect 3285 -1184 3295 -1163
rect 2375 -1186 3295 -1184
rect 3359 -1184 3368 -1163
rect 3514 -1163 3597 -1158
rect 3514 -1184 3523 -1163
rect 3359 -1186 3523 -1184
rect 3587 -1184 3597 -1163
rect 4497 -1163 4580 -1158
rect 4497 -1184 4507 -1163
rect 3587 -1186 4507 -1184
rect 4571 -1184 4580 -1163
rect 4726 -1163 4809 -1158
rect 4726 -1184 4735 -1163
rect 4571 -1186 4735 -1184
rect 4799 -1184 4809 -1163
rect 5458 -1160 5541 -1155
rect 5458 -1181 5467 -1160
rect 5352 -1183 5467 -1181
rect 5531 -1181 5541 -1160
rect 6811 -1165 6937 -1155
rect 5531 -1183 6024 -1181
rect 4799 -1186 5292 -1184
rect 378 -1250 482 -1186
rect 546 -1250 562 -1186
rect 626 -1250 642 -1186
rect 706 -1250 722 -1186
rect 786 -1250 802 -1186
rect 866 -1227 871 -1186
rect 866 -1250 882 -1227
rect 946 -1250 1088 -1186
rect 1163 -1227 1168 -1186
rect 1152 -1250 1168 -1227
rect 1232 -1250 1248 -1186
rect 1312 -1250 1328 -1186
rect 1392 -1250 1408 -1186
rect 1472 -1250 1488 -1186
rect 1552 -1250 1694 -1186
rect 1758 -1250 1774 -1186
rect 1838 -1250 1854 -1186
rect 1918 -1250 1934 -1186
rect 1998 -1250 2014 -1186
rect 2078 -1227 2083 -1186
rect 2078 -1250 2094 -1227
rect 2158 -1250 2300 -1186
rect 2375 -1227 2380 -1186
rect 2364 -1250 2380 -1227
rect 2444 -1250 2460 -1186
rect 2524 -1250 2540 -1186
rect 2604 -1250 2620 -1186
rect 2684 -1250 2700 -1186
rect 2764 -1250 2906 -1186
rect 2970 -1250 2986 -1186
rect 3050 -1250 3066 -1186
rect 3130 -1250 3146 -1186
rect 3210 -1250 3226 -1186
rect 3290 -1227 3295 -1186
rect 3290 -1250 3306 -1227
rect 3370 -1250 3512 -1186
rect 3587 -1227 3592 -1186
rect 3576 -1250 3592 -1227
rect 3656 -1250 3672 -1186
rect 3736 -1250 3752 -1186
rect 3816 -1250 3832 -1186
rect 3896 -1250 3912 -1186
rect 3976 -1250 4118 -1186
rect 4182 -1250 4198 -1186
rect 4262 -1250 4278 -1186
rect 4342 -1250 4358 -1186
rect 4422 -1250 4438 -1186
rect 4502 -1227 4507 -1186
rect 4502 -1250 4518 -1227
rect 4582 -1250 4724 -1186
rect 4799 -1227 4804 -1186
rect 4788 -1250 4804 -1227
rect 4868 -1250 4884 -1186
rect 4948 -1250 4964 -1186
rect 5028 -1250 5044 -1186
rect 5108 -1250 5124 -1186
rect 5188 -1250 5292 -1186
rect 378 -1252 5292 -1250
rect 378 -1406 444 -1252
rect 190 -1426 316 -1416
rect 190 -1490 221 -1426
rect 285 -1490 316 -1426
rect 190 -1500 316 -1490
rect 378 -1470 379 -1406
rect 443 -1470 444 -1406
rect 378 -1486 444 -1470
rect 378 -1550 379 -1486
rect 443 -1550 444 -1486
rect 378 -1566 444 -1550
rect 378 -1630 379 -1566
rect 443 -1630 444 -1566
rect 378 -1646 444 -1630
rect 108 -1668 234 -1658
rect 108 -1732 139 -1668
rect 203 -1732 234 -1668
rect 108 -1742 234 -1732
rect 378 -1710 379 -1646
rect 443 -1710 444 -1646
rect 378 -1726 444 -1710
rect 378 -1790 379 -1726
rect 443 -1790 444 -1726
rect 378 -1806 444 -1790
rect 107 -1825 233 -1815
rect 107 -1889 138 -1825
rect 202 -1889 233 -1825
rect 107 -1899 233 -1889
rect 378 -1870 379 -1806
rect 443 -1870 444 -1806
rect 378 -1886 444 -1870
rect 378 -1950 379 -1886
rect 443 -1950 444 -1886
rect 378 -1966 444 -1950
rect 107 -1995 233 -1985
rect 107 -2059 138 -1995
rect 202 -2059 233 -1995
rect 107 -2069 233 -2059
rect 378 -2030 379 -1966
rect 443 -2030 444 -1966
rect 378 -2046 444 -2030
rect 378 -2110 379 -2046
rect 443 -2110 444 -2046
rect 378 -2126 444 -2110
rect 108 -2147 234 -2137
rect 108 -2211 139 -2147
rect 203 -2211 234 -2147
rect 108 -2221 234 -2211
rect 378 -2190 379 -2126
rect 443 -2190 444 -2126
rect 378 -2280 444 -2190
rect 113 -2291 239 -2281
rect 504 -2284 564 -1252
rect 113 -2355 144 -2291
rect 208 -2355 239 -2291
rect 624 -2344 684 -1314
rect 744 -2284 804 -1252
rect 864 -2344 924 -1314
rect 984 -1406 1050 -1252
rect 984 -1470 985 -1406
rect 1049 -1470 1050 -1406
rect 984 -1486 1050 -1470
rect 984 -1550 985 -1486
rect 1049 -1550 1050 -1486
rect 984 -1566 1050 -1550
rect 984 -1630 985 -1566
rect 1049 -1630 1050 -1566
rect 984 -1646 1050 -1630
rect 984 -1710 985 -1646
rect 1049 -1710 1050 -1646
rect 984 -1726 1050 -1710
rect 984 -1790 985 -1726
rect 1049 -1790 1050 -1726
rect 984 -1806 1050 -1790
rect 984 -1870 985 -1806
rect 1049 -1870 1050 -1806
rect 984 -1886 1050 -1870
rect 984 -1950 985 -1886
rect 1049 -1950 1050 -1886
rect 984 -1966 1050 -1950
rect 984 -2030 985 -1966
rect 1049 -2030 1050 -1966
rect 984 -2046 1050 -2030
rect 984 -2110 985 -2046
rect 1049 -2110 1050 -2046
rect 984 -2126 1050 -2110
rect 984 -2190 985 -2126
rect 1049 -2190 1050 -2126
rect 984 -2280 1050 -2190
rect 1110 -2344 1170 -1314
rect 1230 -2284 1290 -1252
rect 1350 -2344 1410 -1314
rect 1470 -2284 1530 -1252
rect 1590 -1406 1656 -1252
rect 1590 -1470 1591 -1406
rect 1655 -1470 1656 -1406
rect 1590 -1486 1656 -1470
rect 1590 -1550 1591 -1486
rect 1655 -1550 1656 -1486
rect 1590 -1566 1656 -1550
rect 1590 -1630 1591 -1566
rect 1655 -1630 1656 -1566
rect 1590 -1646 1656 -1630
rect 1590 -1710 1591 -1646
rect 1655 -1710 1656 -1646
rect 1590 -1726 1656 -1710
rect 1590 -1790 1591 -1726
rect 1655 -1790 1656 -1726
rect 1590 -1806 1656 -1790
rect 1590 -1870 1591 -1806
rect 1655 -1870 1656 -1806
rect 1590 -1886 1656 -1870
rect 1590 -1950 1591 -1886
rect 1655 -1950 1656 -1886
rect 1590 -1966 1656 -1950
rect 1590 -2030 1591 -1966
rect 1655 -2030 1656 -1966
rect 1590 -2046 1656 -2030
rect 1590 -2110 1591 -2046
rect 1655 -2110 1656 -2046
rect 1590 -2126 1656 -2110
rect 1590 -2190 1591 -2126
rect 1655 -2190 1656 -2126
rect 1590 -2280 1656 -2190
rect 1716 -2284 1776 -1252
rect 1836 -2344 1896 -1314
rect 1956 -2284 2016 -1252
rect 2076 -2344 2136 -1314
rect 2196 -1406 2262 -1252
rect 2196 -1470 2197 -1406
rect 2261 -1470 2262 -1406
rect 2196 -1486 2262 -1470
rect 2196 -1550 2197 -1486
rect 2261 -1550 2262 -1486
rect 2196 -1566 2262 -1550
rect 2196 -1630 2197 -1566
rect 2261 -1630 2262 -1566
rect 2196 -1646 2262 -1630
rect 2196 -1710 2197 -1646
rect 2261 -1710 2262 -1646
rect 2196 -1726 2262 -1710
rect 2196 -1790 2197 -1726
rect 2261 -1790 2262 -1726
rect 2196 -1806 2262 -1790
rect 2196 -1870 2197 -1806
rect 2261 -1870 2262 -1806
rect 2196 -1886 2262 -1870
rect 2196 -1950 2197 -1886
rect 2261 -1950 2262 -1886
rect 2196 -1966 2262 -1950
rect 2196 -2030 2197 -1966
rect 2261 -2030 2262 -1966
rect 2196 -2046 2262 -2030
rect 2196 -2110 2197 -2046
rect 2261 -2110 2262 -2046
rect 2196 -2126 2262 -2110
rect 2196 -2190 2197 -2126
rect 2261 -2190 2262 -2126
rect 2196 -2280 2262 -2190
rect 2322 -2344 2382 -1314
rect 2442 -2284 2502 -1252
rect 2562 -2344 2622 -1314
rect 2682 -2284 2742 -1252
rect 2802 -1406 2868 -1252
rect 2802 -1470 2803 -1406
rect 2867 -1470 2868 -1406
rect 2802 -1486 2868 -1470
rect 2802 -1550 2803 -1486
rect 2867 -1550 2868 -1486
rect 2802 -1566 2868 -1550
rect 2802 -1630 2803 -1566
rect 2867 -1630 2868 -1566
rect 2802 -1646 2868 -1630
rect 2802 -1710 2803 -1646
rect 2867 -1710 2868 -1646
rect 2802 -1726 2868 -1710
rect 2802 -1790 2803 -1726
rect 2867 -1790 2868 -1726
rect 2802 -1806 2868 -1790
rect 2802 -1870 2803 -1806
rect 2867 -1870 2868 -1806
rect 2802 -1886 2868 -1870
rect 2802 -1950 2803 -1886
rect 2867 -1950 2868 -1886
rect 2802 -1966 2868 -1950
rect 2802 -2030 2803 -1966
rect 2867 -2030 2868 -1966
rect 2802 -2046 2868 -2030
rect 2802 -2110 2803 -2046
rect 2867 -2110 2868 -2046
rect 2802 -2126 2868 -2110
rect 2802 -2190 2803 -2126
rect 2867 -2190 2868 -2126
rect 2802 -2280 2868 -2190
rect 2928 -2284 2988 -1252
rect 3048 -2344 3108 -1314
rect 3168 -2284 3228 -1252
rect 3288 -2344 3348 -1314
rect 3408 -1406 3474 -1252
rect 3408 -1470 3409 -1406
rect 3473 -1470 3474 -1406
rect 3408 -1486 3474 -1470
rect 3408 -1550 3409 -1486
rect 3473 -1550 3474 -1486
rect 3408 -1566 3474 -1550
rect 3408 -1630 3409 -1566
rect 3473 -1630 3474 -1566
rect 3408 -1646 3474 -1630
rect 3408 -1710 3409 -1646
rect 3473 -1710 3474 -1646
rect 3408 -1726 3474 -1710
rect 3408 -1790 3409 -1726
rect 3473 -1790 3474 -1726
rect 3408 -1806 3474 -1790
rect 3408 -1870 3409 -1806
rect 3473 -1870 3474 -1806
rect 3408 -1886 3474 -1870
rect 3408 -1950 3409 -1886
rect 3473 -1950 3474 -1886
rect 3408 -1966 3474 -1950
rect 3408 -2030 3409 -1966
rect 3473 -2030 3474 -1966
rect 3408 -2046 3474 -2030
rect 3408 -2110 3409 -2046
rect 3473 -2110 3474 -2046
rect 3408 -2126 3474 -2110
rect 3408 -2190 3409 -2126
rect 3473 -2190 3474 -2126
rect 3408 -2280 3474 -2190
rect 3534 -2344 3594 -1314
rect 3654 -2284 3714 -1252
rect 3774 -2344 3834 -1314
rect 3894 -2284 3954 -1252
rect 4014 -1406 4080 -1252
rect 4014 -1470 4015 -1406
rect 4079 -1470 4080 -1406
rect 4014 -1486 4080 -1470
rect 4014 -1550 4015 -1486
rect 4079 -1550 4080 -1486
rect 4014 -1566 4080 -1550
rect 4014 -1630 4015 -1566
rect 4079 -1630 4080 -1566
rect 4014 -1646 4080 -1630
rect 4014 -1710 4015 -1646
rect 4079 -1710 4080 -1646
rect 4014 -1726 4080 -1710
rect 4014 -1790 4015 -1726
rect 4079 -1790 4080 -1726
rect 4014 -1806 4080 -1790
rect 4014 -1870 4015 -1806
rect 4079 -1870 4080 -1806
rect 4014 -1886 4080 -1870
rect 4014 -1950 4015 -1886
rect 4079 -1950 4080 -1886
rect 4014 -1966 4080 -1950
rect 4014 -2030 4015 -1966
rect 4079 -2030 4080 -1966
rect 4014 -2046 4080 -2030
rect 4014 -2110 4015 -2046
rect 4079 -2110 4080 -2046
rect 4014 -2126 4080 -2110
rect 4014 -2190 4015 -2126
rect 4079 -2190 4080 -2126
rect 4014 -2280 4080 -2190
rect 4140 -2284 4200 -1252
rect 4260 -2344 4320 -1314
rect 4380 -2284 4440 -1252
rect 4500 -2344 4560 -1314
rect 4620 -1406 4686 -1252
rect 4620 -1470 4621 -1406
rect 4685 -1470 4686 -1406
rect 4620 -1486 4686 -1470
rect 4620 -1550 4621 -1486
rect 4685 -1550 4686 -1486
rect 4620 -1566 4686 -1550
rect 4620 -1630 4621 -1566
rect 4685 -1630 4686 -1566
rect 4620 -1646 4686 -1630
rect 4620 -1710 4621 -1646
rect 4685 -1710 4686 -1646
rect 4620 -1726 4686 -1710
rect 4620 -1790 4621 -1726
rect 4685 -1790 4686 -1726
rect 4620 -1806 4686 -1790
rect 4620 -1870 4621 -1806
rect 4685 -1870 4686 -1806
rect 4620 -1886 4686 -1870
rect 4620 -1950 4621 -1886
rect 4685 -1950 4686 -1886
rect 4620 -1966 4686 -1950
rect 4620 -2030 4621 -1966
rect 4685 -2030 4686 -1966
rect 4620 -2046 4686 -2030
rect 4620 -2110 4621 -2046
rect 4685 -2110 4686 -2046
rect 4620 -2126 4686 -2110
rect 4620 -2190 4621 -2126
rect 4685 -2190 4686 -2126
rect 4620 -2280 4686 -2190
rect 4746 -2344 4806 -1314
rect 4866 -2284 4926 -1252
rect 4986 -2344 5046 -1314
rect 5106 -2284 5166 -1252
rect 5226 -1406 5292 -1252
rect 5226 -1470 5227 -1406
rect 5291 -1470 5292 -1406
rect 5226 -1486 5292 -1470
rect 5226 -1550 5227 -1486
rect 5291 -1550 5292 -1486
rect 5226 -1566 5292 -1550
rect 5226 -1630 5227 -1566
rect 5291 -1630 5292 -1566
rect 5226 -1646 5292 -1630
rect 5226 -1710 5227 -1646
rect 5291 -1710 5292 -1646
rect 5226 -1726 5292 -1710
rect 5226 -1790 5227 -1726
rect 5291 -1790 5292 -1726
rect 5226 -1806 5292 -1790
rect 5226 -1870 5227 -1806
rect 5291 -1870 5292 -1806
rect 5226 -1886 5292 -1870
rect 5226 -1950 5227 -1886
rect 5291 -1950 5292 -1886
rect 5226 -1966 5292 -1950
rect 5226 -2030 5227 -1966
rect 5291 -2030 5292 -1966
rect 5226 -2046 5292 -2030
rect 5226 -2110 5227 -2046
rect 5291 -2110 5292 -2046
rect 5226 -2126 5292 -2110
rect 5226 -2190 5227 -2126
rect 5291 -2190 5292 -2126
rect 5226 -2280 5292 -2190
rect 5352 -1247 5456 -1183
rect 5531 -1224 5536 -1183
rect 5520 -1247 5536 -1224
rect 5600 -1247 5616 -1183
rect 5680 -1247 5696 -1183
rect 5760 -1247 5776 -1183
rect 5840 -1247 5856 -1183
rect 5920 -1247 6024 -1183
rect 5352 -1249 6024 -1247
rect 5352 -1403 5418 -1249
rect 5352 -1467 5353 -1403
rect 5417 -1467 5418 -1403
rect 5352 -1483 5418 -1467
rect 5352 -1547 5353 -1483
rect 5417 -1547 5418 -1483
rect 5352 -1563 5418 -1547
rect 5352 -1627 5353 -1563
rect 5417 -1627 5418 -1563
rect 5352 -1643 5418 -1627
rect 5352 -1707 5353 -1643
rect 5417 -1707 5418 -1643
rect 5352 -1723 5418 -1707
rect 5352 -1787 5353 -1723
rect 5417 -1787 5418 -1723
rect 5352 -1803 5418 -1787
rect 5352 -1867 5353 -1803
rect 5417 -1867 5418 -1803
rect 5352 -1883 5418 -1867
rect 5352 -1947 5353 -1883
rect 5417 -1947 5418 -1883
rect 5352 -1963 5418 -1947
rect 5352 -2027 5353 -1963
rect 5417 -2027 5418 -1963
rect 5352 -2043 5418 -2027
rect 5352 -2107 5353 -2043
rect 5417 -2107 5418 -2043
rect 5352 -2123 5418 -2107
rect 5352 -2187 5353 -2123
rect 5417 -2187 5418 -2123
rect 5352 -2277 5418 -2187
rect 5478 -2341 5538 -1311
rect 5598 -2281 5658 -1249
rect 5718 -2341 5778 -1311
rect 5838 -2281 5898 -1249
rect 5958 -1403 6024 -1249
rect 6250 -1202 6623 -1185
rect 6250 -1266 6289 -1202
rect 6353 -1266 6432 -1202
rect 6496 -1266 6552 -1202
rect 6616 -1266 6623 -1202
rect 6811 -1229 6842 -1165
rect 6906 -1229 6937 -1165
rect 7570 -1163 7653 -1158
rect 7570 -1184 7580 -1163
rect 6811 -1239 6937 -1229
rect 7087 -1186 7580 -1184
rect 7644 -1184 7653 -1163
rect 7799 -1163 7882 -1158
rect 7799 -1184 7808 -1163
rect 7644 -1186 7808 -1184
rect 7872 -1184 7882 -1163
rect 8782 -1163 8865 -1158
rect 8782 -1184 8792 -1163
rect 7872 -1186 8792 -1184
rect 8856 -1184 8865 -1163
rect 9011 -1163 9094 -1158
rect 9011 -1184 9020 -1163
rect 8856 -1186 9020 -1184
rect 9084 -1184 9094 -1163
rect 9994 -1163 10077 -1158
rect 9994 -1184 10004 -1163
rect 9084 -1186 10004 -1184
rect 10068 -1184 10077 -1163
rect 10223 -1163 10306 -1158
rect 10223 -1184 10232 -1163
rect 10068 -1186 10232 -1184
rect 10296 -1184 10306 -1163
rect 11206 -1163 11289 -1158
rect 11206 -1184 11216 -1163
rect 10296 -1186 11216 -1184
rect 11280 -1184 11289 -1163
rect 11435 -1163 11518 -1158
rect 11435 -1184 11444 -1163
rect 11280 -1186 11444 -1184
rect 11508 -1184 11518 -1163
rect 12167 -1160 12250 -1155
rect 12167 -1181 12176 -1160
rect 12061 -1183 12176 -1181
rect 12240 -1181 12250 -1160
rect 12240 -1183 12733 -1181
rect 11508 -1186 12001 -1184
rect 6250 -1281 6623 -1266
rect 7087 -1250 7191 -1186
rect 7255 -1250 7271 -1186
rect 7335 -1250 7351 -1186
rect 7415 -1250 7431 -1186
rect 7495 -1250 7511 -1186
rect 7575 -1227 7580 -1186
rect 7575 -1250 7591 -1227
rect 7655 -1250 7797 -1186
rect 7872 -1227 7877 -1186
rect 7861 -1250 7877 -1227
rect 7941 -1250 7957 -1186
rect 8021 -1250 8037 -1186
rect 8101 -1250 8117 -1186
rect 8181 -1250 8197 -1186
rect 8261 -1250 8403 -1186
rect 8467 -1250 8483 -1186
rect 8547 -1250 8563 -1186
rect 8627 -1250 8643 -1186
rect 8707 -1250 8723 -1186
rect 8787 -1227 8792 -1186
rect 8787 -1250 8803 -1227
rect 8867 -1250 9009 -1186
rect 9084 -1227 9089 -1186
rect 9073 -1250 9089 -1227
rect 9153 -1250 9169 -1186
rect 9233 -1250 9249 -1186
rect 9313 -1250 9329 -1186
rect 9393 -1250 9409 -1186
rect 9473 -1250 9615 -1186
rect 9679 -1250 9695 -1186
rect 9759 -1250 9775 -1186
rect 9839 -1250 9855 -1186
rect 9919 -1250 9935 -1186
rect 9999 -1227 10004 -1186
rect 9999 -1250 10015 -1227
rect 10079 -1250 10221 -1186
rect 10296 -1227 10301 -1186
rect 10285 -1250 10301 -1227
rect 10365 -1250 10381 -1186
rect 10445 -1250 10461 -1186
rect 10525 -1250 10541 -1186
rect 10605 -1250 10621 -1186
rect 10685 -1250 10827 -1186
rect 10891 -1250 10907 -1186
rect 10971 -1250 10987 -1186
rect 11051 -1250 11067 -1186
rect 11131 -1250 11147 -1186
rect 11211 -1227 11216 -1186
rect 11211 -1250 11227 -1227
rect 11291 -1250 11433 -1186
rect 11508 -1227 11513 -1186
rect 11497 -1250 11513 -1227
rect 11577 -1250 11593 -1186
rect 11657 -1250 11673 -1186
rect 11737 -1250 11753 -1186
rect 11817 -1250 11833 -1186
rect 11897 -1250 12001 -1186
rect 7087 -1252 12001 -1250
rect 6417 -1282 6509 -1281
rect 5958 -1467 5959 -1403
rect 6023 -1467 6024 -1403
rect 7087 -1406 7153 -1252
rect 5958 -1483 6024 -1467
rect 5958 -1547 5959 -1483
rect 6023 -1547 6024 -1483
rect 6899 -1426 7025 -1416
rect 6899 -1490 6930 -1426
rect 6994 -1490 7025 -1426
rect 6899 -1500 7025 -1490
rect 7087 -1470 7088 -1406
rect 7152 -1470 7153 -1406
rect 7087 -1486 7153 -1470
rect 5958 -1563 6024 -1547
rect 5958 -1627 5959 -1563
rect 6023 -1627 6024 -1563
rect 5958 -1643 6024 -1627
rect 5958 -1707 5959 -1643
rect 6023 -1707 6024 -1643
rect 7087 -1550 7088 -1486
rect 7152 -1550 7153 -1486
rect 7087 -1566 7153 -1550
rect 7087 -1630 7088 -1566
rect 7152 -1630 7153 -1566
rect 7087 -1646 7153 -1630
rect 5958 -1723 6024 -1707
rect 5958 -1787 5959 -1723
rect 6023 -1787 6024 -1723
rect 6817 -1668 6943 -1658
rect 6400 -1731 6544 -1730
rect 5958 -1803 6024 -1787
rect 5958 -1867 5959 -1803
rect 6023 -1867 6024 -1803
rect 6256 -1747 6649 -1731
rect 6817 -1732 6848 -1668
rect 6912 -1732 6943 -1668
rect 6817 -1742 6943 -1732
rect 7087 -1710 7088 -1646
rect 7152 -1710 7153 -1646
rect 7087 -1726 7153 -1710
rect 6256 -1748 6439 -1747
rect 6256 -1812 6295 -1748
rect 6359 -1811 6439 -1748
rect 6503 -1748 6649 -1747
rect 6503 -1811 6570 -1748
rect 6359 -1812 6570 -1811
rect 6634 -1812 6649 -1748
rect 6256 -1826 6649 -1812
rect 7087 -1790 7088 -1726
rect 7152 -1790 7153 -1726
rect 7087 -1806 7153 -1790
rect 6256 -1827 6400 -1826
rect 6531 -1827 6649 -1826
rect 6816 -1825 6942 -1815
rect 5958 -1883 6024 -1867
rect 5958 -1947 5959 -1883
rect 6023 -1947 6024 -1883
rect 5958 -1963 6024 -1947
rect 5958 -2027 5959 -1963
rect 6023 -2027 6024 -1963
rect 6394 -1897 6520 -1887
rect 6394 -1961 6425 -1897
rect 6489 -1961 6520 -1897
rect 6816 -1889 6847 -1825
rect 6911 -1889 6942 -1825
rect 6816 -1899 6942 -1889
rect 7087 -1870 7088 -1806
rect 7152 -1870 7153 -1806
rect 7087 -1886 7153 -1870
rect 6394 -1971 6520 -1961
rect 7087 -1950 7088 -1886
rect 7152 -1950 7153 -1886
rect 7087 -1966 7153 -1950
rect 5958 -2043 6024 -2027
rect 5958 -2107 5959 -2043
rect 6023 -2107 6024 -2043
rect 6816 -1995 6942 -1985
rect 6816 -2059 6847 -1995
rect 6911 -2059 6942 -1995
rect 6816 -2069 6942 -2059
rect 7087 -2030 7088 -1966
rect 7152 -2030 7153 -1966
rect 7087 -2046 7153 -2030
rect 5958 -2123 6024 -2107
rect 5958 -2187 5959 -2123
rect 6023 -2187 6024 -2123
rect 6394 -2093 6520 -2083
rect 6394 -2157 6425 -2093
rect 6489 -2157 6520 -2093
rect 7087 -2110 7088 -2046
rect 7152 -2110 7153 -2046
rect 7087 -2126 7153 -2110
rect 6394 -2167 6520 -2157
rect 6817 -2147 6943 -2137
rect 5958 -2277 6024 -2187
rect 6817 -2211 6848 -2147
rect 6912 -2211 6943 -2147
rect 6817 -2221 6943 -2211
rect 7087 -2190 7088 -2126
rect 7152 -2190 7153 -2126
rect 6394 -2268 6520 -2258
rect 6394 -2332 6425 -2268
rect 6489 -2332 6520 -2268
rect 7087 -2280 7153 -2190
rect 5352 -2343 6024 -2341
rect 6394 -2342 6520 -2332
rect 6822 -2291 6948 -2281
rect 7213 -2284 7273 -1252
rect 113 -2365 239 -2355
rect 378 -2346 5292 -2344
rect 378 -2410 482 -2346
rect 546 -2410 562 -2346
rect 626 -2410 642 -2346
rect 706 -2410 722 -2346
rect 786 -2410 802 -2346
rect 866 -2410 882 -2346
rect 946 -2410 1088 -2346
rect 1152 -2410 1168 -2346
rect 1232 -2410 1248 -2346
rect 1312 -2410 1328 -2346
rect 1392 -2410 1408 -2346
rect 1472 -2410 1488 -2346
rect 1552 -2410 1694 -2346
rect 1758 -2410 1774 -2346
rect 1838 -2410 1854 -2346
rect 1918 -2410 1934 -2346
rect 1998 -2410 2014 -2346
rect 2078 -2410 2094 -2346
rect 2158 -2410 2300 -2346
rect 2364 -2410 2380 -2346
rect 2444 -2410 2460 -2346
rect 2524 -2410 2540 -2346
rect 2604 -2410 2620 -2346
rect 2684 -2410 2700 -2346
rect 2764 -2410 2906 -2346
rect 2970 -2410 2986 -2346
rect 3050 -2410 3066 -2346
rect 3130 -2410 3146 -2346
rect 3210 -2410 3226 -2346
rect 3290 -2410 3306 -2346
rect 3370 -2410 3512 -2346
rect 3576 -2410 3592 -2346
rect 3656 -2410 3672 -2346
rect 3736 -2410 3752 -2346
rect 3816 -2410 3832 -2346
rect 3896 -2410 3912 -2346
rect 3976 -2410 4118 -2346
rect 4182 -2410 4198 -2346
rect 4262 -2410 4278 -2346
rect 4342 -2410 4358 -2346
rect 4422 -2410 4438 -2346
rect 4502 -2410 4518 -2346
rect 4582 -2410 4724 -2346
rect 4788 -2410 4804 -2346
rect 4868 -2410 4884 -2346
rect 4948 -2410 4964 -2346
rect 5028 -2410 5044 -2346
rect 5108 -2410 5124 -2346
rect 5188 -2410 5292 -2346
rect 5352 -2407 5456 -2343
rect 5520 -2407 5536 -2343
rect 5600 -2407 5616 -2343
rect 5680 -2407 5696 -2343
rect 5760 -2407 5776 -2343
rect 5840 -2407 5856 -2343
rect 5920 -2344 6024 -2343
rect 5920 -2353 6048 -2344
rect 5920 -2407 5953 -2353
rect 5352 -2409 5953 -2407
rect 378 -2412 5292 -2410
rect 5922 -2417 5953 -2409
rect 6017 -2417 6048 -2353
rect 6822 -2355 6853 -2291
rect 6917 -2355 6948 -2291
rect 7333 -2344 7393 -1314
rect 7453 -2284 7513 -1252
rect 7573 -2344 7633 -1314
rect 7693 -1406 7759 -1252
rect 7693 -1470 7694 -1406
rect 7758 -1470 7759 -1406
rect 7693 -1486 7759 -1470
rect 7693 -1550 7694 -1486
rect 7758 -1550 7759 -1486
rect 7693 -1566 7759 -1550
rect 7693 -1630 7694 -1566
rect 7758 -1630 7759 -1566
rect 7693 -1646 7759 -1630
rect 7693 -1710 7694 -1646
rect 7758 -1710 7759 -1646
rect 7693 -1726 7759 -1710
rect 7693 -1790 7694 -1726
rect 7758 -1790 7759 -1726
rect 7693 -1806 7759 -1790
rect 7693 -1870 7694 -1806
rect 7758 -1870 7759 -1806
rect 7693 -1886 7759 -1870
rect 7693 -1950 7694 -1886
rect 7758 -1950 7759 -1886
rect 7693 -1966 7759 -1950
rect 7693 -2030 7694 -1966
rect 7758 -2030 7759 -1966
rect 7693 -2046 7759 -2030
rect 7693 -2110 7694 -2046
rect 7758 -2110 7759 -2046
rect 7693 -2126 7759 -2110
rect 7693 -2190 7694 -2126
rect 7758 -2190 7759 -2126
rect 7693 -2280 7759 -2190
rect 7819 -2344 7879 -1314
rect 7939 -2284 7999 -1252
rect 8059 -2344 8119 -1314
rect 8179 -2284 8239 -1252
rect 8299 -1406 8365 -1252
rect 8299 -1470 8300 -1406
rect 8364 -1470 8365 -1406
rect 8299 -1486 8365 -1470
rect 8299 -1550 8300 -1486
rect 8364 -1550 8365 -1486
rect 8299 -1566 8365 -1550
rect 8299 -1630 8300 -1566
rect 8364 -1630 8365 -1566
rect 8299 -1646 8365 -1630
rect 8299 -1710 8300 -1646
rect 8364 -1710 8365 -1646
rect 8299 -1726 8365 -1710
rect 8299 -1790 8300 -1726
rect 8364 -1790 8365 -1726
rect 8299 -1806 8365 -1790
rect 8299 -1870 8300 -1806
rect 8364 -1870 8365 -1806
rect 8299 -1886 8365 -1870
rect 8299 -1950 8300 -1886
rect 8364 -1950 8365 -1886
rect 8299 -1966 8365 -1950
rect 8299 -2030 8300 -1966
rect 8364 -2030 8365 -1966
rect 8299 -2046 8365 -2030
rect 8299 -2110 8300 -2046
rect 8364 -2110 8365 -2046
rect 8299 -2126 8365 -2110
rect 8299 -2190 8300 -2126
rect 8364 -2190 8365 -2126
rect 8299 -2280 8365 -2190
rect 8425 -2284 8485 -1252
rect 8545 -2344 8605 -1314
rect 8665 -2284 8725 -1252
rect 8785 -2344 8845 -1314
rect 8905 -1406 8971 -1252
rect 8905 -1470 8906 -1406
rect 8970 -1470 8971 -1406
rect 8905 -1486 8971 -1470
rect 8905 -1550 8906 -1486
rect 8970 -1550 8971 -1486
rect 8905 -1566 8971 -1550
rect 8905 -1630 8906 -1566
rect 8970 -1630 8971 -1566
rect 8905 -1646 8971 -1630
rect 8905 -1710 8906 -1646
rect 8970 -1710 8971 -1646
rect 8905 -1726 8971 -1710
rect 8905 -1790 8906 -1726
rect 8970 -1790 8971 -1726
rect 8905 -1806 8971 -1790
rect 8905 -1870 8906 -1806
rect 8970 -1870 8971 -1806
rect 8905 -1886 8971 -1870
rect 8905 -1950 8906 -1886
rect 8970 -1950 8971 -1886
rect 8905 -1966 8971 -1950
rect 8905 -2030 8906 -1966
rect 8970 -2030 8971 -1966
rect 8905 -2046 8971 -2030
rect 8905 -2110 8906 -2046
rect 8970 -2110 8971 -2046
rect 8905 -2126 8971 -2110
rect 8905 -2190 8906 -2126
rect 8970 -2190 8971 -2126
rect 8905 -2280 8971 -2190
rect 9031 -2344 9091 -1314
rect 9151 -2284 9211 -1252
rect 9271 -2344 9331 -1314
rect 9391 -2284 9451 -1252
rect 9511 -1406 9577 -1252
rect 9511 -1470 9512 -1406
rect 9576 -1470 9577 -1406
rect 9511 -1486 9577 -1470
rect 9511 -1550 9512 -1486
rect 9576 -1550 9577 -1486
rect 9511 -1566 9577 -1550
rect 9511 -1630 9512 -1566
rect 9576 -1630 9577 -1566
rect 9511 -1646 9577 -1630
rect 9511 -1710 9512 -1646
rect 9576 -1710 9577 -1646
rect 9511 -1726 9577 -1710
rect 9511 -1790 9512 -1726
rect 9576 -1790 9577 -1726
rect 9511 -1806 9577 -1790
rect 9511 -1870 9512 -1806
rect 9576 -1870 9577 -1806
rect 9511 -1886 9577 -1870
rect 9511 -1950 9512 -1886
rect 9576 -1950 9577 -1886
rect 9511 -1966 9577 -1950
rect 9511 -2030 9512 -1966
rect 9576 -2030 9577 -1966
rect 9511 -2046 9577 -2030
rect 9511 -2110 9512 -2046
rect 9576 -2110 9577 -2046
rect 9511 -2126 9577 -2110
rect 9511 -2190 9512 -2126
rect 9576 -2190 9577 -2126
rect 9511 -2280 9577 -2190
rect 9637 -2284 9697 -1252
rect 9757 -2344 9817 -1314
rect 9877 -2284 9937 -1252
rect 9997 -2344 10057 -1314
rect 10117 -1406 10183 -1252
rect 10117 -1470 10118 -1406
rect 10182 -1470 10183 -1406
rect 10117 -1486 10183 -1470
rect 10117 -1550 10118 -1486
rect 10182 -1550 10183 -1486
rect 10117 -1566 10183 -1550
rect 10117 -1630 10118 -1566
rect 10182 -1630 10183 -1566
rect 10117 -1646 10183 -1630
rect 10117 -1710 10118 -1646
rect 10182 -1710 10183 -1646
rect 10117 -1726 10183 -1710
rect 10117 -1790 10118 -1726
rect 10182 -1790 10183 -1726
rect 10117 -1806 10183 -1790
rect 10117 -1870 10118 -1806
rect 10182 -1870 10183 -1806
rect 10117 -1886 10183 -1870
rect 10117 -1950 10118 -1886
rect 10182 -1950 10183 -1886
rect 10117 -1966 10183 -1950
rect 10117 -2030 10118 -1966
rect 10182 -2030 10183 -1966
rect 10117 -2046 10183 -2030
rect 10117 -2110 10118 -2046
rect 10182 -2110 10183 -2046
rect 10117 -2126 10183 -2110
rect 10117 -2190 10118 -2126
rect 10182 -2190 10183 -2126
rect 10117 -2280 10183 -2190
rect 10243 -2344 10303 -1314
rect 10363 -2284 10423 -1252
rect 10483 -2344 10543 -1314
rect 10603 -2284 10663 -1252
rect 10723 -1406 10789 -1252
rect 10723 -1470 10724 -1406
rect 10788 -1470 10789 -1406
rect 10723 -1486 10789 -1470
rect 10723 -1550 10724 -1486
rect 10788 -1550 10789 -1486
rect 10723 -1566 10789 -1550
rect 10723 -1630 10724 -1566
rect 10788 -1630 10789 -1566
rect 10723 -1646 10789 -1630
rect 10723 -1710 10724 -1646
rect 10788 -1710 10789 -1646
rect 10723 -1726 10789 -1710
rect 10723 -1790 10724 -1726
rect 10788 -1790 10789 -1726
rect 10723 -1806 10789 -1790
rect 10723 -1870 10724 -1806
rect 10788 -1870 10789 -1806
rect 10723 -1886 10789 -1870
rect 10723 -1950 10724 -1886
rect 10788 -1950 10789 -1886
rect 10723 -1966 10789 -1950
rect 10723 -2030 10724 -1966
rect 10788 -2030 10789 -1966
rect 10723 -2046 10789 -2030
rect 10723 -2110 10724 -2046
rect 10788 -2110 10789 -2046
rect 10723 -2126 10789 -2110
rect 10723 -2190 10724 -2126
rect 10788 -2190 10789 -2126
rect 10723 -2280 10789 -2190
rect 10849 -2284 10909 -1252
rect 10969 -2344 11029 -1314
rect 11089 -2284 11149 -1252
rect 11209 -2344 11269 -1314
rect 11329 -1406 11395 -1252
rect 11329 -1470 11330 -1406
rect 11394 -1470 11395 -1406
rect 11329 -1486 11395 -1470
rect 11329 -1550 11330 -1486
rect 11394 -1550 11395 -1486
rect 11329 -1566 11395 -1550
rect 11329 -1630 11330 -1566
rect 11394 -1630 11395 -1566
rect 11329 -1646 11395 -1630
rect 11329 -1710 11330 -1646
rect 11394 -1710 11395 -1646
rect 11329 -1726 11395 -1710
rect 11329 -1790 11330 -1726
rect 11394 -1790 11395 -1726
rect 11329 -1806 11395 -1790
rect 11329 -1870 11330 -1806
rect 11394 -1870 11395 -1806
rect 11329 -1886 11395 -1870
rect 11329 -1950 11330 -1886
rect 11394 -1950 11395 -1886
rect 11329 -1966 11395 -1950
rect 11329 -2030 11330 -1966
rect 11394 -2030 11395 -1966
rect 11329 -2046 11395 -2030
rect 11329 -2110 11330 -2046
rect 11394 -2110 11395 -2046
rect 11329 -2126 11395 -2110
rect 11329 -2190 11330 -2126
rect 11394 -2190 11395 -2126
rect 11329 -2280 11395 -2190
rect 11455 -2344 11515 -1314
rect 11575 -2284 11635 -1252
rect 11695 -2344 11755 -1314
rect 11815 -2284 11875 -1252
rect 11935 -1406 12001 -1252
rect 11935 -1470 11936 -1406
rect 12000 -1470 12001 -1406
rect 11935 -1486 12001 -1470
rect 11935 -1550 11936 -1486
rect 12000 -1550 12001 -1486
rect 11935 -1566 12001 -1550
rect 11935 -1630 11936 -1566
rect 12000 -1630 12001 -1566
rect 11935 -1646 12001 -1630
rect 11935 -1710 11936 -1646
rect 12000 -1710 12001 -1646
rect 11935 -1726 12001 -1710
rect 11935 -1790 11936 -1726
rect 12000 -1790 12001 -1726
rect 11935 -1806 12001 -1790
rect 11935 -1870 11936 -1806
rect 12000 -1870 12001 -1806
rect 11935 -1886 12001 -1870
rect 11935 -1950 11936 -1886
rect 12000 -1950 12001 -1886
rect 11935 -1966 12001 -1950
rect 11935 -2030 11936 -1966
rect 12000 -2030 12001 -1966
rect 11935 -2046 12001 -2030
rect 11935 -2110 11936 -2046
rect 12000 -2110 12001 -2046
rect 11935 -2126 12001 -2110
rect 11935 -2190 11936 -2126
rect 12000 -2190 12001 -2126
rect 11935 -2280 12001 -2190
rect 12061 -1247 12165 -1183
rect 12240 -1224 12245 -1183
rect 12229 -1247 12245 -1224
rect 12309 -1247 12325 -1183
rect 12389 -1247 12405 -1183
rect 12469 -1247 12485 -1183
rect 12549 -1247 12565 -1183
rect 12629 -1247 12733 -1183
rect 12061 -1249 12733 -1247
rect 12061 -1403 12127 -1249
rect 12061 -1467 12062 -1403
rect 12126 -1467 12127 -1403
rect 12061 -1483 12127 -1467
rect 12061 -1547 12062 -1483
rect 12126 -1547 12127 -1483
rect 12061 -1563 12127 -1547
rect 12061 -1627 12062 -1563
rect 12126 -1627 12127 -1563
rect 12061 -1643 12127 -1627
rect 12061 -1707 12062 -1643
rect 12126 -1707 12127 -1643
rect 12061 -1723 12127 -1707
rect 12061 -1787 12062 -1723
rect 12126 -1787 12127 -1723
rect 12061 -1803 12127 -1787
rect 12061 -1867 12062 -1803
rect 12126 -1867 12127 -1803
rect 12061 -1883 12127 -1867
rect 12061 -1947 12062 -1883
rect 12126 -1947 12127 -1883
rect 12061 -1963 12127 -1947
rect 12061 -2027 12062 -1963
rect 12126 -2027 12127 -1963
rect 12061 -2043 12127 -2027
rect 12061 -2107 12062 -2043
rect 12126 -2107 12127 -2043
rect 12061 -2123 12127 -2107
rect 12061 -2187 12062 -2123
rect 12126 -2187 12127 -2123
rect 12061 -2277 12127 -2187
rect 12187 -2341 12247 -1311
rect 12307 -2281 12367 -1249
rect 12427 -2341 12487 -1311
rect 12547 -2281 12607 -1249
rect 12667 -1403 12733 -1249
rect 12959 -1202 13332 -1185
rect 12959 -1266 12998 -1202
rect 13062 -1266 13141 -1202
rect 13205 -1266 13261 -1202
rect 13325 -1266 13332 -1202
rect 12959 -1281 13332 -1266
rect 13126 -1282 13218 -1281
rect 12667 -1467 12668 -1403
rect 12732 -1467 12733 -1403
rect 12667 -1483 12733 -1467
rect 12667 -1547 12668 -1483
rect 12732 -1547 12733 -1483
rect 12667 -1563 12733 -1547
rect 12667 -1627 12668 -1563
rect 12732 -1627 12733 -1563
rect 12667 -1643 12733 -1627
rect 12667 -1707 12668 -1643
rect 12732 -1707 12733 -1643
rect 12667 -1723 12733 -1707
rect 12667 -1787 12668 -1723
rect 12732 -1787 12733 -1723
rect 13109 -1731 13253 -1730
rect 12667 -1803 12733 -1787
rect 12667 -1867 12668 -1803
rect 12732 -1867 12733 -1803
rect 12965 -1747 13358 -1731
rect 12965 -1748 13148 -1747
rect 12965 -1812 13004 -1748
rect 13068 -1811 13148 -1748
rect 13212 -1748 13358 -1747
rect 13212 -1811 13279 -1748
rect 13068 -1812 13279 -1811
rect 13343 -1812 13358 -1748
rect 12965 -1826 13358 -1812
rect 12965 -1827 13109 -1826
rect 13240 -1827 13358 -1826
rect 12667 -1883 12733 -1867
rect 12667 -1947 12668 -1883
rect 12732 -1947 12733 -1883
rect 12667 -1963 12733 -1947
rect 12667 -2027 12668 -1963
rect 12732 -2027 12733 -1963
rect 12667 -2043 12733 -2027
rect 12667 -2107 12668 -2043
rect 12732 -2107 12733 -2043
rect 12667 -2123 12733 -2107
rect 12667 -2187 12668 -2123
rect 12732 -2187 12733 -2123
rect 12667 -2277 12733 -2187
rect 12061 -2343 12733 -2341
rect 6822 -2365 6948 -2355
rect 7087 -2346 12001 -2344
rect 7087 -2410 7191 -2346
rect 7255 -2410 7271 -2346
rect 7335 -2410 7351 -2346
rect 7415 -2410 7431 -2346
rect 7495 -2410 7511 -2346
rect 7575 -2410 7591 -2346
rect 7655 -2410 7797 -2346
rect 7861 -2410 7877 -2346
rect 7941 -2410 7957 -2346
rect 8021 -2410 8037 -2346
rect 8101 -2410 8117 -2346
rect 8181 -2410 8197 -2346
rect 8261 -2410 8403 -2346
rect 8467 -2410 8483 -2346
rect 8547 -2410 8563 -2346
rect 8627 -2410 8643 -2346
rect 8707 -2410 8723 -2346
rect 8787 -2410 8803 -2346
rect 8867 -2410 9009 -2346
rect 9073 -2410 9089 -2346
rect 9153 -2410 9169 -2346
rect 9233 -2410 9249 -2346
rect 9313 -2410 9329 -2346
rect 9393 -2410 9409 -2346
rect 9473 -2410 9615 -2346
rect 9679 -2410 9695 -2346
rect 9759 -2410 9775 -2346
rect 9839 -2410 9855 -2346
rect 9919 -2410 9935 -2346
rect 9999 -2410 10015 -2346
rect 10079 -2410 10221 -2346
rect 10285 -2410 10301 -2346
rect 10365 -2410 10381 -2346
rect 10445 -2410 10461 -2346
rect 10525 -2410 10541 -2346
rect 10605 -2410 10621 -2346
rect 10685 -2410 10827 -2346
rect 10891 -2410 10907 -2346
rect 10971 -2410 10987 -2346
rect 11051 -2410 11067 -2346
rect 11131 -2410 11147 -2346
rect 11211 -2410 11227 -2346
rect 11291 -2410 11433 -2346
rect 11497 -2410 11513 -2346
rect 11577 -2410 11593 -2346
rect 11657 -2410 11673 -2346
rect 11737 -2410 11753 -2346
rect 11817 -2410 11833 -2346
rect 11897 -2410 12001 -2346
rect 12061 -2407 12165 -2343
rect 12229 -2407 12245 -2343
rect 12309 -2407 12325 -2343
rect 12389 -2407 12405 -2343
rect 12469 -2407 12485 -2343
rect 12549 -2407 12565 -2343
rect 12629 -2344 12733 -2343
rect 12629 -2353 12757 -2344
rect 12629 -2407 12662 -2353
rect 12061 -2409 12662 -2407
rect 7087 -2412 12001 -2410
rect 5922 -2427 6048 -2417
rect 12631 -2417 12662 -2409
rect 12726 -2417 12757 -2353
rect 12631 -2427 12757 -2417
<< via3 >>
rect 738 3734 802 3738
rect 738 3678 742 3734
rect 742 3678 798 3734
rect 798 3678 802 3734
rect 738 3674 802 3678
rect 835 3725 899 3728
rect 835 3669 838 3725
rect 838 3669 894 3725
rect 894 3669 899 3725
rect 835 3664 899 3669
rect 915 3725 979 3728
rect 915 3669 918 3725
rect 918 3669 974 3725
rect 974 3669 979 3725
rect 915 3664 979 3669
rect 995 3725 1059 3728
rect 995 3669 998 3725
rect 998 3669 1054 3725
rect 1054 3669 1059 3725
rect 995 3664 1059 3669
rect 1075 3725 1139 3728
rect 1075 3669 1078 3725
rect 1078 3669 1134 3725
rect 1134 3669 1139 3725
rect 1075 3664 1139 3669
rect 1155 3725 1219 3728
rect 1155 3669 1158 3725
rect 1158 3669 1214 3725
rect 1214 3669 1219 3725
rect 1155 3664 1219 3669
rect 1235 3725 1299 3728
rect 1235 3669 1238 3725
rect 1238 3669 1294 3725
rect 1294 3669 1299 3725
rect 1235 3664 1299 3669
rect 1567 3728 1631 3731
rect 1567 3672 1570 3728
rect 1570 3672 1626 3728
rect 1626 3672 1631 3728
rect 1567 3667 1631 3672
rect 1647 3728 1711 3731
rect 1647 3672 1650 3728
rect 1650 3672 1706 3728
rect 1706 3672 1711 3728
rect 1647 3667 1711 3672
rect 1727 3728 1791 3731
rect 1727 3672 1730 3728
rect 1730 3672 1786 3728
rect 1786 3672 1791 3728
rect 1727 3667 1791 3672
rect 1807 3728 1871 3731
rect 1807 3672 1810 3728
rect 1810 3672 1866 3728
rect 1866 3672 1871 3728
rect 1807 3667 1871 3672
rect 1887 3728 1951 3731
rect 1887 3672 1890 3728
rect 1890 3672 1946 3728
rect 1946 3672 1951 3728
rect 1887 3667 1951 3672
rect 1967 3728 2031 3731
rect 1967 3672 1970 3728
rect 1970 3672 2026 3728
rect 2026 3672 2031 3728
rect 1967 3667 2031 3672
rect 2173 3728 2237 3731
rect 2173 3672 2178 3728
rect 2178 3672 2234 3728
rect 2234 3672 2237 3728
rect 2173 3667 2237 3672
rect 2253 3728 2317 3731
rect 2253 3672 2258 3728
rect 2258 3672 2314 3728
rect 2314 3672 2317 3728
rect 2253 3667 2317 3672
rect 2333 3728 2397 3731
rect 2333 3672 2338 3728
rect 2338 3672 2394 3728
rect 2394 3672 2397 3728
rect 2333 3667 2397 3672
rect 2413 3728 2477 3731
rect 2413 3672 2418 3728
rect 2418 3672 2474 3728
rect 2474 3672 2477 3728
rect 2413 3667 2477 3672
rect 2493 3728 2557 3731
rect 2493 3672 2498 3728
rect 2498 3672 2554 3728
rect 2554 3672 2557 3728
rect 2493 3667 2557 3672
rect 2573 3728 2637 3731
rect 2573 3672 2578 3728
rect 2578 3672 2634 3728
rect 2634 3672 2637 3728
rect 2573 3667 2637 3672
rect 2779 3728 2843 3731
rect 2779 3672 2782 3728
rect 2782 3672 2838 3728
rect 2838 3672 2843 3728
rect 2779 3667 2843 3672
rect 2859 3728 2923 3731
rect 2859 3672 2862 3728
rect 2862 3672 2918 3728
rect 2918 3672 2923 3728
rect 2859 3667 2923 3672
rect 2939 3728 3003 3731
rect 2939 3672 2942 3728
rect 2942 3672 2998 3728
rect 2998 3672 3003 3728
rect 2939 3667 3003 3672
rect 3019 3728 3083 3731
rect 3019 3672 3022 3728
rect 3022 3672 3078 3728
rect 3078 3672 3083 3728
rect 3019 3667 3083 3672
rect 3099 3728 3163 3731
rect 3099 3672 3102 3728
rect 3102 3672 3158 3728
rect 3158 3672 3163 3728
rect 3099 3667 3163 3672
rect 3179 3728 3243 3731
rect 3179 3672 3182 3728
rect 3182 3672 3238 3728
rect 3238 3672 3243 3728
rect 3179 3667 3243 3672
rect 3385 3728 3449 3731
rect 3385 3672 3390 3728
rect 3390 3672 3446 3728
rect 3446 3672 3449 3728
rect 3385 3667 3449 3672
rect 3465 3728 3529 3731
rect 3465 3672 3470 3728
rect 3470 3672 3526 3728
rect 3526 3672 3529 3728
rect 3465 3667 3529 3672
rect 3545 3728 3609 3731
rect 3545 3672 3550 3728
rect 3550 3672 3606 3728
rect 3606 3672 3609 3728
rect 3545 3667 3609 3672
rect 3625 3728 3689 3731
rect 3625 3672 3630 3728
rect 3630 3672 3686 3728
rect 3686 3672 3689 3728
rect 3625 3667 3689 3672
rect 3705 3728 3769 3731
rect 3705 3672 3710 3728
rect 3710 3672 3766 3728
rect 3766 3672 3769 3728
rect 3705 3667 3769 3672
rect 3785 3728 3849 3731
rect 3785 3672 3790 3728
rect 3790 3672 3846 3728
rect 3846 3672 3849 3728
rect 3785 3667 3849 3672
rect 3991 3728 4055 3731
rect 3991 3672 3994 3728
rect 3994 3672 4050 3728
rect 4050 3672 4055 3728
rect 3991 3667 4055 3672
rect 4071 3728 4135 3731
rect 4071 3672 4074 3728
rect 4074 3672 4130 3728
rect 4130 3672 4135 3728
rect 4071 3667 4135 3672
rect 4151 3728 4215 3731
rect 4151 3672 4154 3728
rect 4154 3672 4210 3728
rect 4210 3672 4215 3728
rect 4151 3667 4215 3672
rect 4231 3728 4295 3731
rect 4231 3672 4234 3728
rect 4234 3672 4290 3728
rect 4290 3672 4295 3728
rect 4231 3667 4295 3672
rect 4311 3728 4375 3731
rect 4311 3672 4314 3728
rect 4314 3672 4370 3728
rect 4370 3672 4375 3728
rect 4311 3667 4375 3672
rect 4391 3728 4455 3731
rect 4391 3672 4394 3728
rect 4394 3672 4450 3728
rect 4450 3672 4455 3728
rect 4391 3667 4455 3672
rect 4597 3728 4661 3731
rect 4597 3672 4602 3728
rect 4602 3672 4658 3728
rect 4658 3672 4661 3728
rect 4597 3667 4661 3672
rect 4677 3728 4741 3731
rect 4677 3672 4682 3728
rect 4682 3672 4738 3728
rect 4738 3672 4741 3728
rect 4677 3667 4741 3672
rect 4757 3728 4821 3731
rect 4757 3672 4762 3728
rect 4762 3672 4818 3728
rect 4818 3672 4821 3728
rect 4757 3667 4821 3672
rect 4837 3728 4901 3731
rect 4837 3672 4842 3728
rect 4842 3672 4898 3728
rect 4898 3672 4901 3728
rect 4837 3667 4901 3672
rect 4917 3728 4981 3731
rect 4917 3672 4922 3728
rect 4922 3672 4978 3728
rect 4978 3672 4981 3728
rect 4917 3667 4981 3672
rect 4997 3728 5061 3731
rect 4997 3672 5002 3728
rect 5002 3672 5058 3728
rect 5058 3672 5061 3728
rect 4997 3667 5061 3672
rect 5203 3728 5267 3731
rect 5203 3672 5206 3728
rect 5206 3672 5262 3728
rect 5262 3672 5267 3728
rect 5203 3667 5267 3672
rect 5283 3728 5347 3731
rect 5283 3672 5286 3728
rect 5286 3672 5342 3728
rect 5342 3672 5347 3728
rect 5283 3667 5347 3672
rect 5363 3728 5427 3731
rect 5363 3672 5366 3728
rect 5366 3672 5422 3728
rect 5422 3672 5427 3728
rect 5363 3667 5427 3672
rect 5443 3728 5507 3731
rect 5443 3672 5446 3728
rect 5446 3672 5502 3728
rect 5502 3672 5507 3728
rect 5443 3667 5507 3672
rect 5523 3728 5587 3731
rect 5523 3672 5526 3728
rect 5526 3672 5582 3728
rect 5582 3672 5587 3728
rect 5523 3667 5587 3672
rect 5603 3728 5667 3731
rect 5603 3672 5606 3728
rect 5606 3672 5662 3728
rect 5662 3672 5667 3728
rect 5603 3667 5667 3672
rect 5809 3728 5873 3731
rect 5809 3672 5814 3728
rect 5814 3672 5870 3728
rect 5870 3672 5873 3728
rect 5809 3667 5873 3672
rect 5889 3728 5953 3731
rect 5889 3672 5894 3728
rect 5894 3672 5950 3728
rect 5950 3672 5953 3728
rect 5889 3667 5953 3672
rect 5969 3728 6033 3731
rect 5969 3672 5974 3728
rect 5974 3672 6030 3728
rect 6030 3672 6033 3728
rect 5969 3667 6033 3672
rect 6049 3728 6113 3731
rect 6049 3672 6054 3728
rect 6054 3672 6110 3728
rect 6110 3672 6113 3728
rect 6049 3667 6113 3672
rect 6129 3728 6193 3731
rect 6129 3672 6134 3728
rect 6134 3672 6190 3728
rect 6190 3672 6193 3728
rect 6129 3667 6193 3672
rect 6209 3728 6273 3731
rect 6209 3672 6214 3728
rect 6214 3672 6270 3728
rect 6270 3672 6273 3728
rect 6209 3667 6273 3672
rect 732 3444 796 3508
rect 732 3364 796 3428
rect 732 3284 796 3348
rect 732 3204 796 3268
rect 121 3129 185 3133
rect 121 3073 125 3129
rect 125 3073 181 3129
rect 181 3073 185 3129
rect 121 3069 185 3073
rect 252 3128 316 3132
rect 252 3072 256 3128
rect 256 3072 312 3128
rect 312 3072 316 3128
rect 252 3068 316 3072
rect 396 3129 460 3133
rect 396 3073 400 3129
rect 400 3073 456 3129
rect 456 3073 460 3129
rect 396 3069 460 3073
rect 732 3124 796 3188
rect 732 3044 796 3108
rect 732 2964 796 3028
rect 732 2884 796 2948
rect 732 2804 796 2868
rect 732 2724 796 2788
rect 139 2583 203 2587
rect 139 2527 143 2583
rect 143 2527 199 2583
rect 199 2527 203 2583
rect 139 2523 203 2527
rect 259 2583 323 2587
rect 259 2527 263 2583
rect 263 2527 319 2583
rect 319 2527 323 2583
rect 259 2523 323 2527
rect 402 2583 466 2587
rect 402 2527 406 2583
rect 406 2527 462 2583
rect 462 2527 466 2583
rect 402 2523 466 2527
rect 1338 3444 1402 3508
rect 1338 3364 1402 3428
rect 1338 3284 1402 3348
rect 1338 3204 1402 3268
rect 1338 3124 1402 3188
rect 1338 3044 1402 3108
rect 1338 2964 1402 3028
rect 1338 2884 1402 2948
rect 1338 2804 1402 2868
rect 1338 2724 1402 2788
rect 835 2504 899 2568
rect 915 2504 979 2568
rect 995 2504 1059 2568
rect 1075 2504 1139 2568
rect 1155 2504 1219 2568
rect 1235 2545 1299 2568
rect 1235 2504 1288 2545
rect 1288 2504 1299 2545
rect 1464 3447 1528 3511
rect 1464 3367 1528 3431
rect 1464 3287 1528 3351
rect 1464 3207 1528 3271
rect 1464 3127 1528 3191
rect 1464 3047 1528 3111
rect 1464 2967 1528 3031
rect 1464 2887 1528 2951
rect 1464 2807 1528 2871
rect 1464 2727 1528 2791
rect 2070 3447 2134 3511
rect 2070 3367 2134 3431
rect 2070 3287 2134 3351
rect 2070 3207 2134 3271
rect 2070 3127 2134 3191
rect 2070 3047 2134 3111
rect 2070 2967 2134 3031
rect 2070 2887 2134 2951
rect 2070 2807 2134 2871
rect 2070 2727 2134 2791
rect 2676 3447 2740 3511
rect 2676 3367 2740 3431
rect 2676 3287 2740 3351
rect 2676 3207 2740 3271
rect 2676 3127 2740 3191
rect 2676 3047 2740 3111
rect 2676 2967 2740 3031
rect 2676 2887 2740 2951
rect 2676 2807 2740 2871
rect 2676 2727 2740 2791
rect 3282 3447 3346 3511
rect 3282 3367 3346 3431
rect 3282 3287 3346 3351
rect 3282 3207 3346 3271
rect 3282 3127 3346 3191
rect 3282 3047 3346 3111
rect 3282 2967 3346 3031
rect 3282 2887 3346 2951
rect 3282 2807 3346 2871
rect 3282 2727 3346 2791
rect 3888 3447 3952 3511
rect 3888 3367 3952 3431
rect 3888 3287 3952 3351
rect 3888 3207 3952 3271
rect 3888 3127 3952 3191
rect 3888 3047 3952 3111
rect 3888 2967 3952 3031
rect 3888 2887 3952 2951
rect 3888 2807 3952 2871
rect 3888 2727 3952 2791
rect 4494 3447 4558 3511
rect 4494 3367 4558 3431
rect 4494 3287 4558 3351
rect 4494 3207 4558 3271
rect 4494 3127 4558 3191
rect 4494 3047 4558 3111
rect 4494 2967 4558 3031
rect 4494 2887 4558 2951
rect 4494 2807 4558 2871
rect 4494 2727 4558 2791
rect 5100 3447 5164 3511
rect 5100 3367 5164 3431
rect 5100 3287 5164 3351
rect 5100 3207 5164 3271
rect 5100 3127 5164 3191
rect 5100 3047 5164 3111
rect 5100 2967 5164 3031
rect 5100 2887 5164 2951
rect 5100 2807 5164 2871
rect 5100 2727 5164 2791
rect 5706 3447 5770 3511
rect 5706 3367 5770 3431
rect 5706 3287 5770 3351
rect 5706 3207 5770 3271
rect 5706 3127 5770 3191
rect 5706 3047 5770 3111
rect 5706 2967 5770 3031
rect 5706 2887 5770 2951
rect 5706 2807 5770 2871
rect 5706 2727 5770 2791
rect 6547 3672 6611 3676
rect 6547 3616 6551 3672
rect 6551 3616 6607 3672
rect 6607 3616 6611 3672
rect 6547 3612 6611 3616
rect 7024 3675 7088 3679
rect 7024 3619 7028 3675
rect 7028 3619 7084 3675
rect 7084 3619 7088 3675
rect 7024 3615 7088 3619
rect 7447 3734 7511 3738
rect 7447 3678 7451 3734
rect 7451 3678 7507 3734
rect 7507 3678 7511 3734
rect 7447 3674 7511 3678
rect 7544 3725 7608 3728
rect 7544 3669 7547 3725
rect 7547 3669 7603 3725
rect 7603 3669 7608 3725
rect 7544 3664 7608 3669
rect 7624 3725 7688 3728
rect 7624 3669 7627 3725
rect 7627 3669 7683 3725
rect 7683 3669 7688 3725
rect 7624 3664 7688 3669
rect 7704 3725 7768 3728
rect 7704 3669 7707 3725
rect 7707 3669 7763 3725
rect 7763 3669 7768 3725
rect 7704 3664 7768 3669
rect 7784 3725 7848 3728
rect 7784 3669 7787 3725
rect 7787 3669 7843 3725
rect 7843 3669 7848 3725
rect 7784 3664 7848 3669
rect 7864 3725 7928 3728
rect 7864 3669 7867 3725
rect 7867 3669 7923 3725
rect 7923 3669 7928 3725
rect 7864 3664 7928 3669
rect 7944 3725 8008 3728
rect 7944 3669 7947 3725
rect 7947 3669 8003 3725
rect 8003 3669 8008 3725
rect 7944 3664 8008 3669
rect 8276 3728 8340 3731
rect 8276 3672 8279 3728
rect 8279 3672 8335 3728
rect 8335 3672 8340 3728
rect 8276 3667 8340 3672
rect 8356 3728 8420 3731
rect 8356 3672 8359 3728
rect 8359 3672 8415 3728
rect 8415 3672 8420 3728
rect 8356 3667 8420 3672
rect 8436 3728 8500 3731
rect 8436 3672 8439 3728
rect 8439 3672 8495 3728
rect 8495 3672 8500 3728
rect 8436 3667 8500 3672
rect 8516 3728 8580 3731
rect 8516 3672 8519 3728
rect 8519 3672 8575 3728
rect 8575 3672 8580 3728
rect 8516 3667 8580 3672
rect 8596 3728 8660 3731
rect 8596 3672 8599 3728
rect 8599 3672 8655 3728
rect 8655 3672 8660 3728
rect 8596 3667 8660 3672
rect 8676 3728 8740 3731
rect 8676 3672 8679 3728
rect 8679 3672 8735 3728
rect 8735 3672 8740 3728
rect 8676 3667 8740 3672
rect 8882 3728 8946 3731
rect 8882 3672 8887 3728
rect 8887 3672 8943 3728
rect 8943 3672 8946 3728
rect 8882 3667 8946 3672
rect 8962 3728 9026 3731
rect 8962 3672 8967 3728
rect 8967 3672 9023 3728
rect 9023 3672 9026 3728
rect 8962 3667 9026 3672
rect 9042 3728 9106 3731
rect 9042 3672 9047 3728
rect 9047 3672 9103 3728
rect 9103 3672 9106 3728
rect 9042 3667 9106 3672
rect 9122 3728 9186 3731
rect 9122 3672 9127 3728
rect 9127 3672 9183 3728
rect 9183 3672 9186 3728
rect 9122 3667 9186 3672
rect 9202 3728 9266 3731
rect 9202 3672 9207 3728
rect 9207 3672 9263 3728
rect 9263 3672 9266 3728
rect 9202 3667 9266 3672
rect 9282 3728 9346 3731
rect 9282 3672 9287 3728
rect 9287 3672 9343 3728
rect 9343 3672 9346 3728
rect 9282 3667 9346 3672
rect 9488 3728 9552 3731
rect 9488 3672 9491 3728
rect 9491 3672 9547 3728
rect 9547 3672 9552 3728
rect 9488 3667 9552 3672
rect 9568 3728 9632 3731
rect 9568 3672 9571 3728
rect 9571 3672 9627 3728
rect 9627 3672 9632 3728
rect 9568 3667 9632 3672
rect 9648 3728 9712 3731
rect 9648 3672 9651 3728
rect 9651 3672 9707 3728
rect 9707 3672 9712 3728
rect 9648 3667 9712 3672
rect 9728 3728 9792 3731
rect 9728 3672 9731 3728
rect 9731 3672 9787 3728
rect 9787 3672 9792 3728
rect 9728 3667 9792 3672
rect 9808 3728 9872 3731
rect 9808 3672 9811 3728
rect 9811 3672 9867 3728
rect 9867 3672 9872 3728
rect 9808 3667 9872 3672
rect 9888 3728 9952 3731
rect 9888 3672 9891 3728
rect 9891 3672 9947 3728
rect 9947 3672 9952 3728
rect 9888 3667 9952 3672
rect 10094 3728 10158 3731
rect 10094 3672 10099 3728
rect 10099 3672 10155 3728
rect 10155 3672 10158 3728
rect 10094 3667 10158 3672
rect 10174 3728 10238 3731
rect 10174 3672 10179 3728
rect 10179 3672 10235 3728
rect 10235 3672 10238 3728
rect 10174 3667 10238 3672
rect 10254 3728 10318 3731
rect 10254 3672 10259 3728
rect 10259 3672 10315 3728
rect 10315 3672 10318 3728
rect 10254 3667 10318 3672
rect 10334 3728 10398 3731
rect 10334 3672 10339 3728
rect 10339 3672 10395 3728
rect 10395 3672 10398 3728
rect 10334 3667 10398 3672
rect 10414 3728 10478 3731
rect 10414 3672 10419 3728
rect 10419 3672 10475 3728
rect 10475 3672 10478 3728
rect 10414 3667 10478 3672
rect 10494 3728 10558 3731
rect 10494 3672 10499 3728
rect 10499 3672 10555 3728
rect 10555 3672 10558 3728
rect 10494 3667 10558 3672
rect 10700 3728 10764 3731
rect 10700 3672 10703 3728
rect 10703 3672 10759 3728
rect 10759 3672 10764 3728
rect 10700 3667 10764 3672
rect 10780 3728 10844 3731
rect 10780 3672 10783 3728
rect 10783 3672 10839 3728
rect 10839 3672 10844 3728
rect 10780 3667 10844 3672
rect 10860 3728 10924 3731
rect 10860 3672 10863 3728
rect 10863 3672 10919 3728
rect 10919 3672 10924 3728
rect 10860 3667 10924 3672
rect 10940 3728 11004 3731
rect 10940 3672 10943 3728
rect 10943 3672 10999 3728
rect 10999 3672 11004 3728
rect 10940 3667 11004 3672
rect 11020 3728 11084 3731
rect 11020 3672 11023 3728
rect 11023 3672 11079 3728
rect 11079 3672 11084 3728
rect 11020 3667 11084 3672
rect 11100 3728 11164 3731
rect 11100 3672 11103 3728
rect 11103 3672 11159 3728
rect 11159 3672 11164 3728
rect 11100 3667 11164 3672
rect 11306 3728 11370 3731
rect 11306 3672 11311 3728
rect 11311 3672 11367 3728
rect 11367 3672 11370 3728
rect 11306 3667 11370 3672
rect 11386 3728 11450 3731
rect 11386 3672 11391 3728
rect 11391 3672 11447 3728
rect 11447 3672 11450 3728
rect 11386 3667 11450 3672
rect 11466 3728 11530 3731
rect 11466 3672 11471 3728
rect 11471 3672 11527 3728
rect 11527 3672 11530 3728
rect 11466 3667 11530 3672
rect 11546 3728 11610 3731
rect 11546 3672 11551 3728
rect 11551 3672 11607 3728
rect 11607 3672 11610 3728
rect 11546 3667 11610 3672
rect 11626 3728 11690 3731
rect 11626 3672 11631 3728
rect 11631 3672 11687 3728
rect 11687 3672 11690 3728
rect 11626 3667 11690 3672
rect 11706 3728 11770 3731
rect 11706 3672 11711 3728
rect 11711 3672 11767 3728
rect 11767 3672 11770 3728
rect 11706 3667 11770 3672
rect 11912 3728 11976 3731
rect 11912 3672 11915 3728
rect 11915 3672 11971 3728
rect 11971 3672 11976 3728
rect 11912 3667 11976 3672
rect 11992 3728 12056 3731
rect 11992 3672 11995 3728
rect 11995 3672 12051 3728
rect 12051 3672 12056 3728
rect 11992 3667 12056 3672
rect 12072 3728 12136 3731
rect 12072 3672 12075 3728
rect 12075 3672 12131 3728
rect 12131 3672 12136 3728
rect 12072 3667 12136 3672
rect 12152 3728 12216 3731
rect 12152 3672 12155 3728
rect 12155 3672 12211 3728
rect 12211 3672 12216 3728
rect 12152 3667 12216 3672
rect 12232 3728 12296 3731
rect 12232 3672 12235 3728
rect 12235 3672 12291 3728
rect 12291 3672 12296 3728
rect 12232 3667 12296 3672
rect 12312 3728 12376 3731
rect 12312 3672 12315 3728
rect 12315 3672 12371 3728
rect 12371 3672 12376 3728
rect 12312 3667 12376 3672
rect 12518 3728 12582 3731
rect 12518 3672 12523 3728
rect 12523 3672 12579 3728
rect 12579 3672 12582 3728
rect 12518 3667 12582 3672
rect 12598 3728 12662 3731
rect 12598 3672 12603 3728
rect 12603 3672 12659 3728
rect 12659 3672 12662 3728
rect 12598 3667 12662 3672
rect 12678 3728 12742 3731
rect 12678 3672 12683 3728
rect 12683 3672 12739 3728
rect 12739 3672 12742 3728
rect 12678 3667 12742 3672
rect 12758 3728 12822 3731
rect 12758 3672 12763 3728
rect 12763 3672 12819 3728
rect 12819 3672 12822 3728
rect 12758 3667 12822 3672
rect 12838 3728 12902 3731
rect 12838 3672 12843 3728
rect 12843 3672 12899 3728
rect 12899 3672 12902 3728
rect 12838 3667 12902 3672
rect 12918 3728 12982 3731
rect 12918 3672 12923 3728
rect 12923 3672 12979 3728
rect 12979 3672 12982 3728
rect 12918 3667 12982 3672
rect 6312 3447 6376 3511
rect 6552 3528 6616 3532
rect 6552 3472 6556 3528
rect 6556 3472 6612 3528
rect 6612 3472 6616 3528
rect 6552 3468 6616 3472
rect 7013 3503 7077 3507
rect 7013 3447 7017 3503
rect 7017 3447 7073 3503
rect 7073 3447 7077 3503
rect 7013 3443 7077 3447
rect 7441 3444 7505 3508
rect 6312 3367 6376 3431
rect 6312 3287 6376 3351
rect 6553 3376 6617 3380
rect 6553 3320 6557 3376
rect 6557 3320 6613 3376
rect 6613 3320 6617 3376
rect 6553 3316 6617 3320
rect 7441 3364 7505 3428
rect 6312 3207 6376 3271
rect 7013 3311 7077 3315
rect 7013 3255 7017 3311
rect 7017 3255 7073 3311
rect 7073 3255 7077 3311
rect 7013 3251 7077 3255
rect 7441 3284 7505 3348
rect 6312 3127 6376 3191
rect 6553 3206 6617 3210
rect 6553 3150 6557 3206
rect 6557 3150 6613 3206
rect 6613 3150 6617 3206
rect 6553 3146 6617 3150
rect 7441 3204 7505 3268
rect 6312 3047 6376 3111
rect 6830 3129 6894 3133
rect 6830 3073 6834 3129
rect 6834 3073 6890 3129
rect 6890 3073 6894 3129
rect 6830 3069 6894 3073
rect 6961 3128 7025 3132
rect 6961 3072 6965 3128
rect 6965 3072 7021 3128
rect 7021 3072 7025 3128
rect 6961 3068 7025 3072
rect 7105 3129 7169 3133
rect 7105 3073 7109 3129
rect 7109 3073 7165 3129
rect 7165 3073 7169 3129
rect 7105 3069 7169 3073
rect 6312 2967 6376 3031
rect 6552 3049 6616 3053
rect 6552 2993 6556 3049
rect 6556 2993 6612 3049
rect 6612 2993 6616 3049
rect 6552 2989 6616 2993
rect 7441 3124 7505 3188
rect 7441 3044 7505 3108
rect 6312 2887 6376 2951
rect 6312 2807 6376 2871
rect 7441 2964 7505 3028
rect 7441 2884 7505 2948
rect 6312 2727 6376 2791
rect 6470 2807 6534 2811
rect 6470 2751 6474 2807
rect 6474 2751 6530 2807
rect 6530 2751 6534 2807
rect 6470 2747 6534 2751
rect 7441 2804 7505 2868
rect 7441 2724 7505 2788
rect 1567 2507 1631 2571
rect 1647 2507 1711 2571
rect 1727 2507 1791 2571
rect 1807 2507 1871 2571
rect 1887 2507 1951 2571
rect 1967 2548 2031 2571
rect 1967 2507 2020 2548
rect 2020 2507 2031 2548
rect 2173 2548 2237 2571
rect 2173 2507 2184 2548
rect 2184 2507 2237 2548
rect 2253 2507 2317 2571
rect 2333 2507 2397 2571
rect 2413 2507 2477 2571
rect 2493 2507 2557 2571
rect 2573 2507 2637 2571
rect 2779 2507 2843 2571
rect 2859 2507 2923 2571
rect 2939 2507 3003 2571
rect 3019 2507 3083 2571
rect 3099 2507 3163 2571
rect 3179 2548 3243 2571
rect 3179 2507 3232 2548
rect 3232 2507 3243 2548
rect 3385 2548 3449 2571
rect 3385 2507 3396 2548
rect 3396 2507 3449 2548
rect 3465 2507 3529 2571
rect 3545 2507 3609 2571
rect 3625 2507 3689 2571
rect 3705 2507 3769 2571
rect 3785 2507 3849 2571
rect 3991 2507 4055 2571
rect 4071 2507 4135 2571
rect 4151 2507 4215 2571
rect 4231 2507 4295 2571
rect 4311 2507 4375 2571
rect 4391 2548 4455 2571
rect 4391 2507 4444 2548
rect 4444 2507 4455 2548
rect 4597 2548 4661 2571
rect 4597 2507 4608 2548
rect 4608 2507 4661 2548
rect 4677 2507 4741 2571
rect 4757 2507 4821 2571
rect 4837 2507 4901 2571
rect 4917 2507 4981 2571
rect 4997 2507 5061 2571
rect 5203 2507 5267 2571
rect 5283 2507 5347 2571
rect 5363 2507 5427 2571
rect 5443 2507 5507 2571
rect 5523 2507 5587 2571
rect 5603 2548 5667 2571
rect 5603 2507 5656 2548
rect 5656 2507 5667 2548
rect 5809 2548 5873 2571
rect 5809 2507 5820 2548
rect 5820 2507 5873 2548
rect 5889 2507 5953 2571
rect 5969 2507 6033 2571
rect 6049 2507 6113 2571
rect 6129 2507 6193 2571
rect 6209 2507 6273 2571
rect 6558 2546 6622 2550
rect 6558 2490 6562 2546
rect 6562 2490 6618 2546
rect 6618 2490 6622 2546
rect 6558 2486 6622 2490
rect 6848 2583 6912 2587
rect 6848 2527 6852 2583
rect 6852 2527 6908 2583
rect 6908 2527 6912 2583
rect 6848 2523 6912 2527
rect 6968 2583 7032 2587
rect 6968 2527 6972 2583
rect 6972 2527 7028 2583
rect 7028 2527 7032 2583
rect 6968 2523 7032 2527
rect 7111 2583 7175 2587
rect 7111 2527 7115 2583
rect 7115 2527 7171 2583
rect 7171 2527 7175 2583
rect 7111 2523 7175 2527
rect 8047 3444 8111 3508
rect 8047 3364 8111 3428
rect 8047 3284 8111 3348
rect 8047 3204 8111 3268
rect 8047 3124 8111 3188
rect 8047 3044 8111 3108
rect 8047 2964 8111 3028
rect 8047 2884 8111 2948
rect 8047 2804 8111 2868
rect 8047 2724 8111 2788
rect 7544 2504 7608 2568
rect 7624 2504 7688 2568
rect 7704 2504 7768 2568
rect 7784 2504 7848 2568
rect 7864 2504 7928 2568
rect 7944 2545 8008 2568
rect 7944 2504 7997 2545
rect 7997 2504 8008 2545
rect 8173 3447 8237 3511
rect 8173 3367 8237 3431
rect 8173 3287 8237 3351
rect 8173 3207 8237 3271
rect 8173 3127 8237 3191
rect 8173 3047 8237 3111
rect 8173 2967 8237 3031
rect 8173 2887 8237 2951
rect 8173 2807 8237 2871
rect 8173 2727 8237 2791
rect 8779 3447 8843 3511
rect 8779 3367 8843 3431
rect 8779 3287 8843 3351
rect 8779 3207 8843 3271
rect 8779 3127 8843 3191
rect 8779 3047 8843 3111
rect 8779 2967 8843 3031
rect 8779 2887 8843 2951
rect 8779 2807 8843 2871
rect 8779 2727 8843 2791
rect 9385 3447 9449 3511
rect 9385 3367 9449 3431
rect 9385 3287 9449 3351
rect 9385 3207 9449 3271
rect 9385 3127 9449 3191
rect 9385 3047 9449 3111
rect 9385 2967 9449 3031
rect 9385 2887 9449 2951
rect 9385 2807 9449 2871
rect 9385 2727 9449 2791
rect 9991 3447 10055 3511
rect 9991 3367 10055 3431
rect 9991 3287 10055 3351
rect 9991 3207 10055 3271
rect 9991 3127 10055 3191
rect 9991 3047 10055 3111
rect 9991 2967 10055 3031
rect 9991 2887 10055 2951
rect 9991 2807 10055 2871
rect 9991 2727 10055 2791
rect 10597 3447 10661 3511
rect 10597 3367 10661 3431
rect 10597 3287 10661 3351
rect 10597 3207 10661 3271
rect 10597 3127 10661 3191
rect 10597 3047 10661 3111
rect 10597 2967 10661 3031
rect 10597 2887 10661 2951
rect 10597 2807 10661 2871
rect 10597 2727 10661 2791
rect 11203 3447 11267 3511
rect 11203 3367 11267 3431
rect 11203 3287 11267 3351
rect 11203 3207 11267 3271
rect 11203 3127 11267 3191
rect 11203 3047 11267 3111
rect 11203 2967 11267 3031
rect 11203 2887 11267 2951
rect 11203 2807 11267 2871
rect 11203 2727 11267 2791
rect 11809 3447 11873 3511
rect 11809 3367 11873 3431
rect 11809 3287 11873 3351
rect 11809 3207 11873 3271
rect 11809 3127 11873 3191
rect 11809 3047 11873 3111
rect 11809 2967 11873 3031
rect 11809 2887 11873 2951
rect 11809 2807 11873 2871
rect 11809 2727 11873 2791
rect 12415 3447 12479 3511
rect 12415 3367 12479 3431
rect 12415 3287 12479 3351
rect 12415 3207 12479 3271
rect 12415 3127 12479 3191
rect 12415 3047 12479 3111
rect 12415 2967 12479 3031
rect 12415 2887 12479 2951
rect 12415 2807 12479 2871
rect 12415 2727 12479 2791
rect 13256 3672 13320 3676
rect 13256 3616 13260 3672
rect 13260 3616 13316 3672
rect 13316 3616 13320 3672
rect 13256 3612 13320 3616
rect 13021 3447 13085 3511
rect 13261 3528 13325 3532
rect 13261 3472 13265 3528
rect 13265 3472 13321 3528
rect 13321 3472 13325 3528
rect 13261 3468 13325 3472
rect 13021 3367 13085 3431
rect 13021 3287 13085 3351
rect 13262 3376 13326 3380
rect 13262 3320 13266 3376
rect 13266 3320 13322 3376
rect 13322 3320 13326 3376
rect 13262 3316 13326 3320
rect 13021 3207 13085 3271
rect 13021 3127 13085 3191
rect 13262 3206 13326 3210
rect 13262 3150 13266 3206
rect 13266 3150 13322 3206
rect 13322 3150 13326 3206
rect 13262 3146 13326 3150
rect 13021 3047 13085 3111
rect 13021 2967 13085 3031
rect 13261 3049 13325 3053
rect 13261 2993 13265 3049
rect 13265 2993 13321 3049
rect 13321 2993 13325 3049
rect 13261 2989 13325 2993
rect 13021 2887 13085 2951
rect 13021 2807 13085 2871
rect 13021 2727 13085 2791
rect 13179 2807 13243 2811
rect 13179 2751 13183 2807
rect 13183 2751 13239 2807
rect 13239 2751 13243 2807
rect 13179 2747 13243 2751
rect 8276 2507 8340 2571
rect 8356 2507 8420 2571
rect 8436 2507 8500 2571
rect 8516 2507 8580 2571
rect 8596 2507 8660 2571
rect 8676 2548 8740 2571
rect 8676 2507 8729 2548
rect 8729 2507 8740 2548
rect 8882 2548 8946 2571
rect 8882 2507 8893 2548
rect 8893 2507 8946 2548
rect 8962 2507 9026 2571
rect 9042 2507 9106 2571
rect 9122 2507 9186 2571
rect 9202 2507 9266 2571
rect 9282 2507 9346 2571
rect 9488 2507 9552 2571
rect 9568 2507 9632 2571
rect 9648 2507 9712 2571
rect 9728 2507 9792 2571
rect 9808 2507 9872 2571
rect 9888 2548 9952 2571
rect 9888 2507 9941 2548
rect 9941 2507 9952 2548
rect 10094 2548 10158 2571
rect 10094 2507 10105 2548
rect 10105 2507 10158 2548
rect 10174 2507 10238 2571
rect 10254 2507 10318 2571
rect 10334 2507 10398 2571
rect 10414 2507 10478 2571
rect 10494 2507 10558 2571
rect 10700 2507 10764 2571
rect 10780 2507 10844 2571
rect 10860 2507 10924 2571
rect 10940 2507 11004 2571
rect 11020 2507 11084 2571
rect 11100 2548 11164 2571
rect 11100 2507 11153 2548
rect 11153 2507 11164 2548
rect 11306 2548 11370 2571
rect 11306 2507 11317 2548
rect 11317 2507 11370 2548
rect 11386 2507 11450 2571
rect 11466 2507 11530 2571
rect 11546 2507 11610 2571
rect 11626 2507 11690 2571
rect 11706 2507 11770 2571
rect 11912 2507 11976 2571
rect 11992 2507 12056 2571
rect 12072 2507 12136 2571
rect 12152 2507 12216 2571
rect 12232 2507 12296 2571
rect 12312 2548 12376 2571
rect 12312 2507 12365 2548
rect 12365 2507 12376 2548
rect 12518 2548 12582 2571
rect 12518 2507 12529 2548
rect 12529 2507 12582 2548
rect 12598 2507 12662 2571
rect 12678 2507 12742 2571
rect 12758 2507 12822 2571
rect 12838 2507 12902 2571
rect 12918 2507 12982 2571
rect 13267 2546 13331 2550
rect 13267 2490 13271 2546
rect 13271 2490 13327 2546
rect 13327 2490 13331 2546
rect 13267 2486 13331 2490
rect 1186 2259 1250 2323
rect 1266 2259 1330 2323
rect 1346 2259 1410 2323
rect 1426 2259 1490 2323
rect 1506 2259 1570 2323
rect 1586 2282 1644 2323
rect 1644 2282 1650 2323
rect 1586 2259 1650 2282
rect 1083 2039 1147 2103
rect 1083 1959 1147 2023
rect 1083 1879 1147 1943
rect 1083 1799 1147 1863
rect 106 1701 171 1707
rect 106 1643 169 1701
rect 169 1643 171 1701
rect 1083 1719 1147 1783
rect 1083 1639 1147 1703
rect 1083 1559 1147 1623
rect 1083 1479 1147 1543
rect 1083 1399 1147 1463
rect 1083 1319 1147 1383
rect 1689 2039 1753 2103
rect 1689 1959 1753 2023
rect 1689 1879 1753 1943
rect 1689 1799 1753 1863
rect 1689 1719 1753 1783
rect 1689 1639 1753 1703
rect 1689 1559 1753 1623
rect 1689 1479 1753 1543
rect 1689 1399 1753 1463
rect 1689 1319 1753 1383
rect 1918 2259 1982 2323
rect 1998 2259 2062 2323
rect 2078 2259 2142 2323
rect 2158 2259 2222 2323
rect 2238 2259 2302 2323
rect 2318 2282 2376 2323
rect 2376 2282 2382 2323
rect 2318 2259 2382 2282
rect 2524 2282 2530 2323
rect 2530 2282 2588 2323
rect 2524 2259 2588 2282
rect 2604 2259 2668 2323
rect 2684 2259 2748 2323
rect 2764 2259 2828 2323
rect 2844 2259 2908 2323
rect 2924 2259 2988 2323
rect 3130 2259 3194 2323
rect 3210 2259 3274 2323
rect 3290 2259 3354 2323
rect 3370 2259 3434 2323
rect 3450 2259 3514 2323
rect 3530 2282 3588 2323
rect 3588 2282 3594 2323
rect 3530 2259 3594 2282
rect 3736 2282 3742 2323
rect 3742 2282 3800 2323
rect 3736 2259 3800 2282
rect 3816 2259 3880 2323
rect 3896 2259 3960 2323
rect 3976 2259 4040 2323
rect 4056 2259 4120 2323
rect 4136 2259 4200 2323
rect 1815 2039 1879 2103
rect 1815 1959 1879 2023
rect 1815 1879 1879 1943
rect 1815 1799 1879 1863
rect 1815 1719 1879 1783
rect 1815 1639 1879 1703
rect 1815 1559 1879 1623
rect 1815 1479 1879 1543
rect 1815 1399 1879 1463
rect 1815 1319 1879 1383
rect 2421 2039 2485 2103
rect 2421 1959 2485 2023
rect 2421 1879 2485 1943
rect 2421 1799 2485 1863
rect 2421 1719 2485 1783
rect 2421 1639 2485 1703
rect 2421 1559 2485 1623
rect 2421 1479 2485 1543
rect 2421 1399 2485 1463
rect 2421 1319 2485 1383
rect 3027 2039 3091 2103
rect 3027 1959 3091 2023
rect 3027 1879 3091 1943
rect 3027 1799 3091 1863
rect 3027 1719 3091 1783
rect 3027 1639 3091 1703
rect 3027 1559 3091 1623
rect 3027 1479 3091 1543
rect 3027 1399 3091 1463
rect 3027 1319 3091 1383
rect 3633 2039 3697 2103
rect 3633 1959 3697 2023
rect 3633 1879 3697 1943
rect 3633 1799 3697 1863
rect 3633 1719 3697 1783
rect 3633 1639 3697 1703
rect 3633 1559 3697 1623
rect 3633 1479 3697 1543
rect 3633 1399 3697 1463
rect 3633 1319 3697 1383
rect 4239 2039 4303 2103
rect 4239 1959 4303 2023
rect 4239 1879 4303 1943
rect 4239 1799 4303 1863
rect 4239 1719 4303 1783
rect 4239 1639 4303 1703
rect 4239 1559 4303 1623
rect 4239 1479 4303 1543
rect 4239 1399 4303 1463
rect 4239 1319 4303 1383
rect 4468 2259 4532 2323
rect 4548 2259 4612 2323
rect 4628 2259 4692 2323
rect 4708 2259 4772 2323
rect 4788 2259 4852 2323
rect 4868 2282 4926 2323
rect 4926 2282 4932 2323
rect 4868 2259 4932 2282
rect 5074 2282 5080 2323
rect 5080 2282 5138 2323
rect 5074 2259 5138 2282
rect 5154 2259 5218 2323
rect 5234 2259 5298 2323
rect 5314 2259 5378 2323
rect 5394 2259 5458 2323
rect 5474 2259 5538 2323
rect 4365 2039 4429 2103
rect 4365 1959 4429 2023
rect 4365 1879 4429 1943
rect 4365 1799 4429 1863
rect 4365 1719 4429 1783
rect 4365 1639 4429 1703
rect 4365 1559 4429 1623
rect 4365 1479 4429 1543
rect 4365 1399 4429 1463
rect 4365 1319 4429 1383
rect 4971 2039 5035 2103
rect 4971 1959 5035 2023
rect 4971 1879 5035 1943
rect 4971 1799 5035 1863
rect 4971 1719 5035 1783
rect 4971 1639 5035 1703
rect 4971 1559 5035 1623
rect 4971 1479 5035 1543
rect 4971 1399 5035 1463
rect 4971 1319 5035 1383
rect 5577 2039 5641 2103
rect 5577 1959 5641 2023
rect 5577 1879 5641 1943
rect 5577 1799 5641 1863
rect 5577 1719 5641 1783
rect 5577 1639 5641 1703
rect 5577 1559 5641 1623
rect 5577 1479 5641 1543
rect 5577 1399 5641 1463
rect 5577 1319 5641 1383
rect 5808 2282 5814 2323
rect 5814 2282 5872 2323
rect 5808 2259 5872 2282
rect 5888 2259 5952 2323
rect 5968 2259 6032 2323
rect 6048 2259 6112 2323
rect 6128 2259 6192 2323
rect 6208 2259 6272 2323
rect 6558 2343 6622 2347
rect 6558 2287 6562 2343
rect 6562 2287 6618 2343
rect 6618 2287 6622 2343
rect 6558 2283 6622 2287
rect 5705 2039 5769 2103
rect 5705 1959 5769 2023
rect 5705 1879 5769 1943
rect 5705 1799 5769 1863
rect 5705 1719 5769 1783
rect 5705 1639 5769 1703
rect 5705 1559 5769 1623
rect 5705 1479 5769 1543
rect 5705 1399 5769 1463
rect 5705 1319 5769 1383
rect 6311 2039 6375 2103
rect 7895 2259 7959 2323
rect 7975 2259 8039 2323
rect 8055 2259 8119 2323
rect 8135 2259 8199 2323
rect 8215 2259 8279 2323
rect 8295 2282 8353 2323
rect 8353 2282 8359 2323
rect 8295 2259 8359 2282
rect 6311 1959 6375 2023
rect 6467 2081 6531 2085
rect 6467 2025 6471 2081
rect 6471 2025 6527 2081
rect 6527 2025 6531 2081
rect 6467 2021 6531 2025
rect 7792 2039 7856 2103
rect 6311 1879 6375 1943
rect 6311 1799 6375 1863
rect 6311 1719 6375 1783
rect 6311 1639 6375 1703
rect 6311 1559 6375 1623
rect 6311 1479 6375 1543
rect 6311 1399 6375 1463
rect 6311 1319 6375 1383
rect 7792 1959 7856 2023
rect 7792 1879 7856 1943
rect 7792 1799 7856 1863
rect 7792 1719 7856 1783
rect 7792 1639 7856 1703
rect 7792 1559 7856 1623
rect 7792 1479 7856 1543
rect 7792 1399 7856 1463
rect 7792 1319 7856 1383
rect 724 1156 788 1160
rect 724 1100 728 1156
rect 728 1100 784 1156
rect 784 1100 788 1156
rect 724 1096 788 1100
rect 1266 1159 1330 1163
rect 1266 1103 1270 1159
rect 1270 1103 1326 1159
rect 1326 1103 1330 1159
rect 1266 1099 1330 1103
rect 1346 1159 1410 1163
rect 1346 1103 1350 1159
rect 1350 1103 1406 1159
rect 1406 1103 1410 1159
rect 1346 1099 1410 1103
rect 1426 1159 1490 1163
rect 1426 1103 1430 1159
rect 1430 1103 1486 1159
rect 1486 1103 1490 1159
rect 1426 1099 1490 1103
rect 1506 1159 1570 1163
rect 1506 1103 1510 1159
rect 1510 1103 1566 1159
rect 1566 1103 1570 1159
rect 1506 1099 1570 1103
rect 1998 1159 2062 1163
rect 1998 1103 2002 1159
rect 2002 1103 2058 1159
rect 2058 1103 2062 1159
rect 1998 1099 2062 1103
rect 2078 1159 2142 1163
rect 2078 1103 2082 1159
rect 2082 1103 2138 1159
rect 2138 1103 2142 1159
rect 2078 1099 2142 1103
rect 2158 1159 2222 1163
rect 2158 1103 2162 1159
rect 2162 1103 2218 1159
rect 2218 1103 2222 1159
rect 2158 1099 2222 1103
rect 2238 1159 2302 1163
rect 2238 1103 2242 1159
rect 2242 1103 2298 1159
rect 2298 1103 2302 1159
rect 2238 1099 2302 1103
rect 2604 1159 2668 1163
rect 2604 1103 2608 1159
rect 2608 1103 2664 1159
rect 2664 1103 2668 1159
rect 2604 1099 2668 1103
rect 2684 1159 2748 1163
rect 2684 1103 2688 1159
rect 2688 1103 2744 1159
rect 2744 1103 2748 1159
rect 2684 1099 2748 1103
rect 2764 1159 2828 1163
rect 2764 1103 2768 1159
rect 2768 1103 2824 1159
rect 2824 1103 2828 1159
rect 2764 1099 2828 1103
rect 2844 1159 2908 1163
rect 2844 1103 2848 1159
rect 2848 1103 2904 1159
rect 2904 1103 2908 1159
rect 2844 1099 2908 1103
rect 3210 1159 3274 1163
rect 3210 1103 3214 1159
rect 3214 1103 3270 1159
rect 3270 1103 3274 1159
rect 3210 1099 3274 1103
rect 3290 1159 3354 1163
rect 3290 1103 3294 1159
rect 3294 1103 3350 1159
rect 3350 1103 3354 1159
rect 3290 1099 3354 1103
rect 3370 1159 3434 1163
rect 3370 1103 3374 1159
rect 3374 1103 3430 1159
rect 3430 1103 3434 1159
rect 3370 1099 3434 1103
rect 3450 1159 3514 1163
rect 3450 1103 3454 1159
rect 3454 1103 3510 1159
rect 3510 1103 3514 1159
rect 3450 1099 3514 1103
rect 3816 1159 3880 1163
rect 3816 1103 3820 1159
rect 3820 1103 3876 1159
rect 3876 1103 3880 1159
rect 3816 1099 3880 1103
rect 3896 1159 3960 1163
rect 3896 1103 3900 1159
rect 3900 1103 3956 1159
rect 3956 1103 3960 1159
rect 3896 1099 3960 1103
rect 3976 1159 4040 1163
rect 3976 1103 3980 1159
rect 3980 1103 4036 1159
rect 4036 1103 4040 1159
rect 3976 1099 4040 1103
rect 4056 1159 4120 1163
rect 4056 1103 4060 1159
rect 4060 1103 4116 1159
rect 4116 1103 4120 1159
rect 4056 1099 4120 1103
rect 4548 1159 4612 1163
rect 4548 1103 4552 1159
rect 4552 1103 4608 1159
rect 4608 1103 4612 1159
rect 4548 1099 4612 1103
rect 4628 1159 4692 1163
rect 4628 1103 4632 1159
rect 4632 1103 4688 1159
rect 4688 1103 4692 1159
rect 4628 1099 4692 1103
rect 4708 1159 4772 1163
rect 4708 1103 4712 1159
rect 4712 1103 4768 1159
rect 4768 1103 4772 1159
rect 4708 1099 4772 1103
rect 4788 1159 4852 1163
rect 4788 1103 4792 1159
rect 4792 1103 4848 1159
rect 4848 1103 4852 1159
rect 4788 1099 4852 1103
rect 5154 1159 5218 1163
rect 5154 1103 5158 1159
rect 5158 1103 5214 1159
rect 5214 1103 5218 1159
rect 5154 1099 5218 1103
rect 5234 1159 5298 1163
rect 5234 1103 5238 1159
rect 5238 1103 5294 1159
rect 5294 1103 5298 1159
rect 5234 1099 5298 1103
rect 5314 1159 5378 1163
rect 5314 1103 5318 1159
rect 5318 1103 5374 1159
rect 5374 1103 5378 1159
rect 5314 1099 5378 1103
rect 5394 1159 5458 1163
rect 5394 1103 5398 1159
rect 5398 1103 5454 1159
rect 5454 1103 5458 1159
rect 5394 1099 5458 1103
rect 5888 1159 5952 1163
rect 5888 1103 5892 1159
rect 5892 1103 5948 1159
rect 5948 1103 5952 1159
rect 5888 1099 5952 1103
rect 5968 1159 6032 1163
rect 5968 1103 5972 1159
rect 5972 1103 6028 1159
rect 6028 1103 6032 1159
rect 5968 1099 6032 1103
rect 6048 1159 6112 1163
rect 6048 1103 6052 1159
rect 6052 1103 6108 1159
rect 6108 1103 6112 1159
rect 6048 1099 6112 1103
rect 6128 1159 6192 1163
rect 6128 1103 6132 1159
rect 6132 1103 6188 1159
rect 6188 1103 6192 1159
rect 6128 1099 6192 1103
rect 8398 2039 8462 2103
rect 8398 1959 8462 2023
rect 8398 1879 8462 1943
rect 8398 1799 8462 1863
rect 8398 1719 8462 1783
rect 8398 1639 8462 1703
rect 8398 1559 8462 1623
rect 8398 1479 8462 1543
rect 8398 1399 8462 1463
rect 8398 1319 8462 1383
rect 8627 2259 8691 2323
rect 8707 2259 8771 2323
rect 8787 2259 8851 2323
rect 8867 2259 8931 2323
rect 8947 2259 9011 2323
rect 9027 2282 9085 2323
rect 9085 2282 9091 2323
rect 9027 2259 9091 2282
rect 9233 2282 9239 2323
rect 9239 2282 9297 2323
rect 9233 2259 9297 2282
rect 9313 2259 9377 2323
rect 9393 2259 9457 2323
rect 9473 2259 9537 2323
rect 9553 2259 9617 2323
rect 9633 2259 9697 2323
rect 9839 2259 9903 2323
rect 9919 2259 9983 2323
rect 9999 2259 10063 2323
rect 10079 2259 10143 2323
rect 10159 2259 10223 2323
rect 10239 2282 10297 2323
rect 10297 2282 10303 2323
rect 10239 2259 10303 2282
rect 10445 2282 10451 2323
rect 10451 2282 10509 2323
rect 10445 2259 10509 2282
rect 10525 2259 10589 2323
rect 10605 2259 10669 2323
rect 10685 2259 10749 2323
rect 10765 2259 10829 2323
rect 10845 2259 10909 2323
rect 8524 2039 8588 2103
rect 8524 1959 8588 2023
rect 8524 1879 8588 1943
rect 8524 1799 8588 1863
rect 8524 1719 8588 1783
rect 8524 1639 8588 1703
rect 8524 1559 8588 1623
rect 8524 1479 8588 1543
rect 8524 1399 8588 1463
rect 8524 1319 8588 1383
rect 9130 2039 9194 2103
rect 9130 1959 9194 2023
rect 9130 1879 9194 1943
rect 9130 1799 9194 1863
rect 9130 1719 9194 1783
rect 9130 1639 9194 1703
rect 9130 1559 9194 1623
rect 9130 1479 9194 1543
rect 9130 1399 9194 1463
rect 9130 1319 9194 1383
rect 9736 2039 9800 2103
rect 9736 1959 9800 2023
rect 9736 1879 9800 1943
rect 9736 1799 9800 1863
rect 9736 1719 9800 1783
rect 9736 1639 9800 1703
rect 9736 1559 9800 1623
rect 9736 1479 9800 1543
rect 9736 1399 9800 1463
rect 9736 1319 9800 1383
rect 10342 2039 10406 2103
rect 10342 1959 10406 2023
rect 10342 1879 10406 1943
rect 10342 1799 10406 1863
rect 10342 1719 10406 1783
rect 10342 1639 10406 1703
rect 10342 1559 10406 1623
rect 10342 1479 10406 1543
rect 10342 1399 10406 1463
rect 10342 1319 10406 1383
rect 10948 2039 11012 2103
rect 10948 1959 11012 2023
rect 10948 1879 11012 1943
rect 10948 1799 11012 1863
rect 10948 1719 11012 1783
rect 10948 1639 11012 1703
rect 10948 1559 11012 1623
rect 10948 1479 11012 1543
rect 10948 1399 11012 1463
rect 10948 1319 11012 1383
rect 11177 2259 11241 2323
rect 11257 2259 11321 2323
rect 11337 2259 11401 2323
rect 11417 2259 11481 2323
rect 11497 2259 11561 2323
rect 11577 2282 11635 2323
rect 11635 2282 11641 2323
rect 11577 2259 11641 2282
rect 11783 2282 11789 2323
rect 11789 2282 11847 2323
rect 11783 2259 11847 2282
rect 11863 2259 11927 2323
rect 11943 2259 12007 2323
rect 12023 2259 12087 2323
rect 12103 2259 12167 2323
rect 12183 2259 12247 2323
rect 11074 2039 11138 2103
rect 11074 1959 11138 2023
rect 11074 1879 11138 1943
rect 11074 1799 11138 1863
rect 11074 1719 11138 1783
rect 11074 1639 11138 1703
rect 11074 1559 11138 1623
rect 11074 1479 11138 1543
rect 11074 1399 11138 1463
rect 11074 1319 11138 1383
rect 11680 2039 11744 2103
rect 11680 1959 11744 2023
rect 11680 1879 11744 1943
rect 11680 1799 11744 1863
rect 11680 1719 11744 1783
rect 11680 1639 11744 1703
rect 11680 1559 11744 1623
rect 11680 1479 11744 1543
rect 11680 1399 11744 1463
rect 11680 1319 11744 1383
rect 12286 2039 12350 2103
rect 12286 1959 12350 2023
rect 12286 1879 12350 1943
rect 12286 1799 12350 1863
rect 12286 1719 12350 1783
rect 12286 1639 12350 1703
rect 12286 1559 12350 1623
rect 12286 1479 12350 1543
rect 12286 1399 12350 1463
rect 12286 1319 12350 1383
rect 12517 2282 12523 2323
rect 12523 2282 12581 2323
rect 12517 2259 12581 2282
rect 12597 2259 12661 2323
rect 12677 2259 12741 2323
rect 12757 2259 12821 2323
rect 12837 2259 12901 2323
rect 12917 2259 12981 2323
rect 13267 2343 13331 2347
rect 13267 2287 13271 2343
rect 13271 2287 13327 2343
rect 13327 2287 13331 2343
rect 13267 2283 13331 2287
rect 12414 2039 12478 2103
rect 12414 1959 12478 2023
rect 12414 1879 12478 1943
rect 12414 1799 12478 1863
rect 12414 1719 12478 1783
rect 12414 1639 12478 1703
rect 12414 1559 12478 1623
rect 12414 1479 12478 1543
rect 12414 1399 12478 1463
rect 12414 1319 12478 1383
rect 13020 2039 13084 2103
rect 13020 1959 13084 2023
rect 13176 2081 13240 2085
rect 13176 2025 13180 2081
rect 13180 2025 13236 2081
rect 13236 2025 13240 2081
rect 13176 2021 13240 2025
rect 13020 1879 13084 1943
rect 13020 1799 13084 1863
rect 13020 1719 13084 1783
rect 13020 1639 13084 1703
rect 13020 1559 13084 1623
rect 13020 1479 13084 1543
rect 13020 1399 13084 1463
rect 13020 1319 13084 1383
rect 7433 1156 7497 1160
rect 7433 1100 7437 1156
rect 7437 1100 7493 1156
rect 7493 1100 7497 1156
rect 7433 1096 7497 1100
rect 7975 1159 8039 1163
rect 7975 1103 7979 1159
rect 7979 1103 8035 1159
rect 8035 1103 8039 1159
rect 7975 1099 8039 1103
rect 8055 1159 8119 1163
rect 8055 1103 8059 1159
rect 8059 1103 8115 1159
rect 8115 1103 8119 1159
rect 8055 1099 8119 1103
rect 8135 1159 8199 1163
rect 8135 1103 8139 1159
rect 8139 1103 8195 1159
rect 8195 1103 8199 1159
rect 8135 1099 8199 1103
rect 8215 1159 8279 1163
rect 8215 1103 8219 1159
rect 8219 1103 8275 1159
rect 8275 1103 8279 1159
rect 8215 1099 8279 1103
rect 8707 1159 8771 1163
rect 8707 1103 8711 1159
rect 8711 1103 8767 1159
rect 8767 1103 8771 1159
rect 8707 1099 8771 1103
rect 8787 1159 8851 1163
rect 8787 1103 8791 1159
rect 8791 1103 8847 1159
rect 8847 1103 8851 1159
rect 8787 1099 8851 1103
rect 8867 1159 8931 1163
rect 8867 1103 8871 1159
rect 8871 1103 8927 1159
rect 8927 1103 8931 1159
rect 8867 1099 8931 1103
rect 8947 1159 9011 1163
rect 8947 1103 8951 1159
rect 8951 1103 9007 1159
rect 9007 1103 9011 1159
rect 8947 1099 9011 1103
rect 9313 1159 9377 1163
rect 9313 1103 9317 1159
rect 9317 1103 9373 1159
rect 9373 1103 9377 1159
rect 9313 1099 9377 1103
rect 9393 1159 9457 1163
rect 9393 1103 9397 1159
rect 9397 1103 9453 1159
rect 9453 1103 9457 1159
rect 9393 1099 9457 1103
rect 9473 1159 9537 1163
rect 9473 1103 9477 1159
rect 9477 1103 9533 1159
rect 9533 1103 9537 1159
rect 9473 1099 9537 1103
rect 9553 1159 9617 1163
rect 9553 1103 9557 1159
rect 9557 1103 9613 1159
rect 9613 1103 9617 1159
rect 9553 1099 9617 1103
rect 9919 1159 9983 1163
rect 9919 1103 9923 1159
rect 9923 1103 9979 1159
rect 9979 1103 9983 1159
rect 9919 1099 9983 1103
rect 9999 1159 10063 1163
rect 9999 1103 10003 1159
rect 10003 1103 10059 1159
rect 10059 1103 10063 1159
rect 9999 1099 10063 1103
rect 10079 1159 10143 1163
rect 10079 1103 10083 1159
rect 10083 1103 10139 1159
rect 10139 1103 10143 1159
rect 10079 1099 10143 1103
rect 10159 1159 10223 1163
rect 10159 1103 10163 1159
rect 10163 1103 10219 1159
rect 10219 1103 10223 1159
rect 10159 1099 10223 1103
rect 10525 1159 10589 1163
rect 10525 1103 10529 1159
rect 10529 1103 10585 1159
rect 10585 1103 10589 1159
rect 10525 1099 10589 1103
rect 10605 1159 10669 1163
rect 10605 1103 10609 1159
rect 10609 1103 10665 1159
rect 10665 1103 10669 1159
rect 10605 1099 10669 1103
rect 10685 1159 10749 1163
rect 10685 1103 10689 1159
rect 10689 1103 10745 1159
rect 10745 1103 10749 1159
rect 10685 1099 10749 1103
rect 10765 1159 10829 1163
rect 10765 1103 10769 1159
rect 10769 1103 10825 1159
rect 10825 1103 10829 1159
rect 10765 1099 10829 1103
rect 11257 1159 11321 1163
rect 11257 1103 11261 1159
rect 11261 1103 11317 1159
rect 11317 1103 11321 1159
rect 11257 1099 11321 1103
rect 11337 1159 11401 1163
rect 11337 1103 11341 1159
rect 11341 1103 11397 1159
rect 11397 1103 11401 1159
rect 11337 1099 11401 1103
rect 11417 1159 11481 1163
rect 11417 1103 11421 1159
rect 11421 1103 11477 1159
rect 11477 1103 11481 1159
rect 11417 1099 11481 1103
rect 11497 1159 11561 1163
rect 11497 1103 11501 1159
rect 11501 1103 11557 1159
rect 11557 1103 11561 1159
rect 11497 1099 11561 1103
rect 11863 1159 11927 1163
rect 11863 1103 11867 1159
rect 11867 1103 11923 1159
rect 11923 1103 11927 1159
rect 11863 1099 11927 1103
rect 11943 1159 12007 1163
rect 11943 1103 11947 1159
rect 11947 1103 12003 1159
rect 12003 1103 12007 1159
rect 11943 1099 12007 1103
rect 12023 1159 12087 1163
rect 12023 1103 12027 1159
rect 12027 1103 12083 1159
rect 12083 1103 12087 1159
rect 12023 1099 12087 1103
rect 12103 1159 12167 1163
rect 12103 1103 12107 1159
rect 12107 1103 12163 1159
rect 12163 1103 12167 1159
rect 12103 1099 12167 1103
rect 12597 1159 12661 1163
rect 12597 1103 12601 1159
rect 12601 1103 12657 1159
rect 12657 1103 12661 1159
rect 12597 1099 12661 1103
rect 12677 1159 12741 1163
rect 12677 1103 12681 1159
rect 12681 1103 12737 1159
rect 12737 1103 12741 1159
rect 12677 1099 12741 1103
rect 12757 1159 12821 1163
rect 12757 1103 12761 1159
rect 12761 1103 12817 1159
rect 12817 1103 12821 1159
rect 12757 1099 12821 1103
rect 12837 1159 12901 1163
rect 12837 1103 12841 1159
rect 12841 1103 12897 1159
rect 12897 1103 12901 1159
rect 12837 1099 12901 1103
rect 563 218 627 222
rect 563 162 567 218
rect 567 162 623 218
rect 623 162 627 218
rect 563 158 627 162
rect 643 218 707 222
rect 643 162 647 218
rect 647 162 703 218
rect 703 162 707 218
rect 643 158 707 162
rect 723 218 787 222
rect 723 162 727 218
rect 727 162 783 218
rect 783 162 787 218
rect 723 158 787 162
rect 803 218 867 222
rect 803 162 807 218
rect 807 162 863 218
rect 863 162 867 218
rect 803 158 867 162
rect 1297 218 1361 222
rect 1297 162 1301 218
rect 1301 162 1357 218
rect 1357 162 1361 218
rect 1297 158 1361 162
rect 1377 218 1441 222
rect 1377 162 1381 218
rect 1381 162 1437 218
rect 1437 162 1441 218
rect 1377 158 1441 162
rect 1457 218 1521 222
rect 1457 162 1461 218
rect 1461 162 1517 218
rect 1517 162 1521 218
rect 1457 158 1521 162
rect 1537 218 1601 222
rect 1537 162 1541 218
rect 1541 162 1597 218
rect 1597 162 1601 218
rect 1537 158 1601 162
rect 1903 218 1967 222
rect 1903 162 1907 218
rect 1907 162 1963 218
rect 1963 162 1967 218
rect 1903 158 1967 162
rect 1983 218 2047 222
rect 1983 162 1987 218
rect 1987 162 2043 218
rect 2043 162 2047 218
rect 1983 158 2047 162
rect 2063 218 2127 222
rect 2063 162 2067 218
rect 2067 162 2123 218
rect 2123 162 2127 218
rect 2063 158 2127 162
rect 2143 218 2207 222
rect 2143 162 2147 218
rect 2147 162 2203 218
rect 2203 162 2207 218
rect 2143 158 2207 162
rect 2635 218 2699 222
rect 2635 162 2639 218
rect 2639 162 2695 218
rect 2695 162 2699 218
rect 2635 158 2699 162
rect 2715 218 2779 222
rect 2715 162 2719 218
rect 2719 162 2775 218
rect 2775 162 2779 218
rect 2715 158 2779 162
rect 2795 218 2859 222
rect 2795 162 2799 218
rect 2799 162 2855 218
rect 2855 162 2859 218
rect 2795 158 2859 162
rect 2875 218 2939 222
rect 2875 162 2879 218
rect 2879 162 2935 218
rect 2935 162 2939 218
rect 2875 158 2939 162
rect 3241 218 3305 222
rect 3241 162 3245 218
rect 3245 162 3301 218
rect 3301 162 3305 218
rect 3241 158 3305 162
rect 3321 218 3385 222
rect 3321 162 3325 218
rect 3325 162 3381 218
rect 3381 162 3385 218
rect 3321 158 3385 162
rect 3401 218 3465 222
rect 3401 162 3405 218
rect 3405 162 3461 218
rect 3461 162 3465 218
rect 3401 158 3465 162
rect 3481 218 3545 222
rect 3481 162 3485 218
rect 3485 162 3541 218
rect 3541 162 3545 218
rect 3481 158 3545 162
rect 3847 218 3911 222
rect 3847 162 3851 218
rect 3851 162 3907 218
rect 3907 162 3911 218
rect 3847 158 3911 162
rect 3927 218 3991 222
rect 3927 162 3931 218
rect 3931 162 3987 218
rect 3987 162 3991 218
rect 3927 158 3991 162
rect 4007 218 4071 222
rect 4007 162 4011 218
rect 4011 162 4067 218
rect 4067 162 4071 218
rect 4007 158 4071 162
rect 4087 218 4151 222
rect 4087 162 4091 218
rect 4091 162 4147 218
rect 4147 162 4151 218
rect 4087 158 4151 162
rect 4453 218 4517 222
rect 4453 162 4457 218
rect 4457 162 4513 218
rect 4513 162 4517 218
rect 4453 158 4517 162
rect 4533 218 4597 222
rect 4533 162 4537 218
rect 4537 162 4593 218
rect 4593 162 4597 218
rect 4533 158 4597 162
rect 4613 218 4677 222
rect 4613 162 4617 218
rect 4617 162 4673 218
rect 4673 162 4677 218
rect 4613 158 4677 162
rect 4693 218 4757 222
rect 4693 162 4697 218
rect 4697 162 4753 218
rect 4753 162 4757 218
rect 4693 158 4757 162
rect 5185 218 5249 222
rect 5185 162 5189 218
rect 5189 162 5245 218
rect 5245 162 5249 218
rect 5185 158 5249 162
rect 5265 218 5329 222
rect 5265 162 5269 218
rect 5269 162 5325 218
rect 5325 162 5329 218
rect 5265 158 5329 162
rect 5345 218 5409 222
rect 5345 162 5349 218
rect 5349 162 5405 218
rect 5405 162 5409 218
rect 5345 158 5409 162
rect 5425 218 5489 222
rect 5425 162 5429 218
rect 5429 162 5485 218
rect 5485 162 5489 218
rect 5425 158 5489 162
rect 5967 221 6031 225
rect 5967 165 5971 221
rect 5971 165 6027 221
rect 6027 165 6031 221
rect 5967 161 6031 165
rect 380 -62 444 2
rect 380 -142 444 -78
rect 380 -222 444 -158
rect 380 -302 444 -238
rect 380 -382 444 -318
rect 380 -462 444 -398
rect 380 -542 444 -478
rect 380 -622 444 -558
rect 224 -704 288 -700
rect 224 -760 228 -704
rect 228 -760 284 -704
rect 284 -760 288 -704
rect 224 -764 288 -760
rect 380 -702 444 -638
rect 380 -782 444 -718
rect 986 -62 1050 2
rect 986 -142 1050 -78
rect 986 -222 1050 -158
rect 986 -302 1050 -238
rect 986 -382 1050 -318
rect 986 -462 1050 -398
rect 986 -542 1050 -478
rect 986 -622 1050 -558
rect 986 -702 1050 -638
rect 986 -782 1050 -718
rect 133 -966 197 -962
rect 133 -1022 137 -966
rect 137 -1022 193 -966
rect 193 -1022 197 -966
rect 133 -1026 197 -1022
rect 483 -1002 547 -938
rect 563 -1002 627 -938
rect 643 -1002 707 -938
rect 723 -1002 787 -938
rect 803 -1002 867 -938
rect 883 -961 947 -938
rect 883 -1002 941 -961
rect 941 -1002 947 -961
rect 1114 -62 1178 2
rect 1114 -142 1178 -78
rect 1114 -222 1178 -158
rect 1114 -302 1178 -238
rect 1114 -382 1178 -318
rect 1114 -462 1178 -398
rect 1114 -542 1178 -478
rect 1114 -622 1178 -558
rect 1114 -702 1178 -638
rect 1114 -782 1178 -718
rect 1720 -62 1784 2
rect 1720 -142 1784 -78
rect 1720 -222 1784 -158
rect 1720 -302 1784 -238
rect 1720 -382 1784 -318
rect 1720 -462 1784 -398
rect 1720 -542 1784 -478
rect 1720 -622 1784 -558
rect 1720 -702 1784 -638
rect 1720 -782 1784 -718
rect 2326 -62 2390 2
rect 2326 -142 2390 -78
rect 2326 -222 2390 -158
rect 2326 -302 2390 -238
rect 2326 -382 2390 -318
rect 2326 -462 2390 -398
rect 2326 -542 2390 -478
rect 2326 -622 2390 -558
rect 2326 -702 2390 -638
rect 2326 -782 2390 -718
rect 1217 -1002 1281 -938
rect 1297 -1002 1361 -938
rect 1377 -1002 1441 -938
rect 1457 -1002 1521 -938
rect 1537 -1002 1601 -938
rect 1617 -961 1681 -938
rect 1617 -1002 1675 -961
rect 1675 -1002 1681 -961
rect 1823 -961 1887 -938
rect 1823 -1002 1829 -961
rect 1829 -1002 1887 -961
rect 1903 -1002 1967 -938
rect 1983 -1002 2047 -938
rect 2063 -1002 2127 -938
rect 2143 -1002 2207 -938
rect 2223 -1002 2287 -938
rect 2452 -62 2516 2
rect 2452 -142 2516 -78
rect 2452 -222 2516 -158
rect 2452 -302 2516 -238
rect 2452 -382 2516 -318
rect 2452 -462 2516 -398
rect 2452 -542 2516 -478
rect 2452 -622 2516 -558
rect 2452 -702 2516 -638
rect 2452 -782 2516 -718
rect 3058 -62 3122 2
rect 3058 -142 3122 -78
rect 3058 -222 3122 -158
rect 3058 -302 3122 -238
rect 3058 -382 3122 -318
rect 3058 -462 3122 -398
rect 3058 -542 3122 -478
rect 3058 -622 3122 -558
rect 3058 -702 3122 -638
rect 3058 -782 3122 -718
rect 3664 -62 3728 2
rect 3664 -142 3728 -78
rect 3664 -222 3728 -158
rect 3664 -302 3728 -238
rect 3664 -382 3728 -318
rect 3664 -462 3728 -398
rect 3664 -542 3728 -478
rect 3664 -622 3728 -558
rect 3664 -702 3728 -638
rect 3664 -782 3728 -718
rect 4270 -62 4334 2
rect 4270 -142 4334 -78
rect 4270 -222 4334 -158
rect 4270 -302 4334 -238
rect 4270 -382 4334 -318
rect 4270 -462 4334 -398
rect 4270 -542 4334 -478
rect 4270 -622 4334 -558
rect 4270 -702 4334 -638
rect 4270 -782 4334 -718
rect 4876 -62 4940 2
rect 4876 -142 4940 -78
rect 4876 -222 4940 -158
rect 4876 -302 4940 -238
rect 4876 -382 4940 -318
rect 4876 -462 4940 -398
rect 4876 -542 4940 -478
rect 4876 -622 4940 -558
rect 4876 -702 4940 -638
rect 4876 -782 4940 -718
rect 2555 -1002 2619 -938
rect 2635 -1002 2699 -938
rect 2715 -1002 2779 -938
rect 2795 -1002 2859 -938
rect 2875 -1002 2939 -938
rect 2955 -961 3019 -938
rect 2955 -1002 3013 -961
rect 3013 -1002 3019 -961
rect 3161 -961 3225 -938
rect 3161 -1002 3167 -961
rect 3167 -1002 3225 -961
rect 3241 -1002 3305 -938
rect 3321 -1002 3385 -938
rect 3401 -1002 3465 -938
rect 3481 -1002 3545 -938
rect 3561 -1002 3625 -938
rect 3767 -1002 3831 -938
rect 3847 -1002 3911 -938
rect 3927 -1002 3991 -938
rect 4007 -1002 4071 -938
rect 4087 -1002 4151 -938
rect 4167 -961 4231 -938
rect 4167 -1002 4225 -961
rect 4225 -1002 4231 -961
rect 4373 -961 4437 -938
rect 4373 -1002 4379 -961
rect 4379 -1002 4437 -961
rect 4453 -1002 4517 -938
rect 4533 -1002 4597 -938
rect 4613 -1002 4677 -938
rect 4693 -1002 4757 -938
rect 4773 -1002 4837 -938
rect 5002 -62 5066 2
rect 5002 -142 5066 -78
rect 5002 -222 5066 -158
rect 5002 -302 5066 -238
rect 5002 -382 5066 -318
rect 5002 -462 5066 -398
rect 5002 -542 5066 -478
rect 5002 -622 5066 -558
rect 5002 -702 5066 -638
rect 5002 -782 5066 -718
rect 7272 218 7336 222
rect 7272 162 7276 218
rect 7276 162 7332 218
rect 7332 162 7336 218
rect 7272 158 7336 162
rect 7352 218 7416 222
rect 7352 162 7356 218
rect 7356 162 7412 218
rect 7412 162 7416 218
rect 7352 158 7416 162
rect 7432 218 7496 222
rect 7432 162 7436 218
rect 7436 162 7492 218
rect 7492 162 7496 218
rect 7432 158 7496 162
rect 7512 218 7576 222
rect 7512 162 7516 218
rect 7516 162 7572 218
rect 7572 162 7576 218
rect 7512 158 7576 162
rect 8006 218 8070 222
rect 8006 162 8010 218
rect 8010 162 8066 218
rect 8066 162 8070 218
rect 8006 158 8070 162
rect 8086 218 8150 222
rect 8086 162 8090 218
rect 8090 162 8146 218
rect 8146 162 8150 218
rect 8086 158 8150 162
rect 8166 218 8230 222
rect 8166 162 8170 218
rect 8170 162 8226 218
rect 8226 162 8230 218
rect 8166 158 8230 162
rect 8246 218 8310 222
rect 8246 162 8250 218
rect 8250 162 8306 218
rect 8306 162 8310 218
rect 8246 158 8310 162
rect 8612 218 8676 222
rect 8612 162 8616 218
rect 8616 162 8672 218
rect 8672 162 8676 218
rect 8612 158 8676 162
rect 8692 218 8756 222
rect 8692 162 8696 218
rect 8696 162 8752 218
rect 8752 162 8756 218
rect 8692 158 8756 162
rect 8772 218 8836 222
rect 8772 162 8776 218
rect 8776 162 8832 218
rect 8832 162 8836 218
rect 8772 158 8836 162
rect 8852 218 8916 222
rect 8852 162 8856 218
rect 8856 162 8912 218
rect 8912 162 8916 218
rect 8852 158 8916 162
rect 9344 218 9408 222
rect 9344 162 9348 218
rect 9348 162 9404 218
rect 9404 162 9408 218
rect 9344 158 9408 162
rect 9424 218 9488 222
rect 9424 162 9428 218
rect 9428 162 9484 218
rect 9484 162 9488 218
rect 9424 158 9488 162
rect 9504 218 9568 222
rect 9504 162 9508 218
rect 9508 162 9564 218
rect 9564 162 9568 218
rect 9504 158 9568 162
rect 9584 218 9648 222
rect 9584 162 9588 218
rect 9588 162 9644 218
rect 9644 162 9648 218
rect 9584 158 9648 162
rect 9950 218 10014 222
rect 9950 162 9954 218
rect 9954 162 10010 218
rect 10010 162 10014 218
rect 9950 158 10014 162
rect 10030 218 10094 222
rect 10030 162 10034 218
rect 10034 162 10090 218
rect 10090 162 10094 218
rect 10030 158 10094 162
rect 10110 218 10174 222
rect 10110 162 10114 218
rect 10114 162 10170 218
rect 10170 162 10174 218
rect 10110 158 10174 162
rect 10190 218 10254 222
rect 10190 162 10194 218
rect 10194 162 10250 218
rect 10250 162 10254 218
rect 10190 158 10254 162
rect 10556 218 10620 222
rect 10556 162 10560 218
rect 10560 162 10616 218
rect 10616 162 10620 218
rect 10556 158 10620 162
rect 10636 218 10700 222
rect 10636 162 10640 218
rect 10640 162 10696 218
rect 10696 162 10700 218
rect 10636 158 10700 162
rect 10716 218 10780 222
rect 10716 162 10720 218
rect 10720 162 10776 218
rect 10776 162 10780 218
rect 10716 158 10780 162
rect 10796 218 10860 222
rect 10796 162 10800 218
rect 10800 162 10856 218
rect 10856 162 10860 218
rect 10796 158 10860 162
rect 11162 218 11226 222
rect 11162 162 11166 218
rect 11166 162 11222 218
rect 11222 162 11226 218
rect 11162 158 11226 162
rect 11242 218 11306 222
rect 11242 162 11246 218
rect 11246 162 11302 218
rect 11302 162 11306 218
rect 11242 158 11306 162
rect 11322 218 11386 222
rect 11322 162 11326 218
rect 11326 162 11382 218
rect 11382 162 11386 218
rect 11322 158 11386 162
rect 11402 218 11466 222
rect 11402 162 11406 218
rect 11406 162 11462 218
rect 11462 162 11466 218
rect 11402 158 11466 162
rect 11894 218 11958 222
rect 11894 162 11898 218
rect 11898 162 11954 218
rect 11954 162 11958 218
rect 11894 158 11958 162
rect 11974 218 12038 222
rect 11974 162 11978 218
rect 11978 162 12034 218
rect 12034 162 12038 218
rect 11974 158 12038 162
rect 12054 218 12118 222
rect 12054 162 12058 218
rect 12058 162 12114 218
rect 12114 162 12118 218
rect 12054 158 12118 162
rect 12134 218 12198 222
rect 12134 162 12138 218
rect 12138 162 12194 218
rect 12194 162 12198 218
rect 12134 158 12198 162
rect 12676 221 12740 225
rect 12676 165 12680 221
rect 12680 165 12736 221
rect 12736 165 12740 221
rect 12676 161 12740 165
rect 5608 -62 5672 2
rect 5608 -142 5672 -78
rect 5608 -222 5672 -158
rect 5608 -302 5672 -238
rect 5608 -382 5672 -318
rect 5608 -462 5672 -398
rect 5608 -542 5672 -478
rect 5608 -622 5672 -558
rect 5608 -702 5672 -638
rect 7089 -62 7153 2
rect 7089 -142 7153 -78
rect 7089 -222 7153 -158
rect 7089 -302 7153 -238
rect 7089 -382 7153 -318
rect 7089 -462 7153 -398
rect 7089 -542 7153 -478
rect 7089 -622 7153 -558
rect 5608 -782 5672 -718
rect 6933 -704 6997 -700
rect 6933 -760 6937 -704
rect 6937 -760 6993 -704
rect 6993 -760 6997 -704
rect 6933 -764 6997 -760
rect 7089 -702 7153 -638
rect 5105 -961 5169 -938
rect 5105 -1002 5111 -961
rect 5111 -1002 5169 -961
rect 5185 -1002 5249 -938
rect 5265 -1002 5329 -938
rect 5345 -1002 5409 -938
rect 5425 -1002 5489 -938
rect 5505 -1002 5569 -938
rect 7089 -782 7153 -718
rect 7695 -62 7759 2
rect 7695 -142 7759 -78
rect 7695 -222 7759 -158
rect 7695 -302 7759 -238
rect 7695 -382 7759 -318
rect 7695 -462 7759 -398
rect 7695 -542 7759 -478
rect 7695 -622 7759 -558
rect 7695 -702 7759 -638
rect 7695 -782 7759 -718
rect 6842 -966 6906 -962
rect 6842 -1022 6846 -966
rect 6846 -1022 6902 -966
rect 6902 -1022 6906 -966
rect 6842 -1026 6906 -1022
rect 7192 -1002 7256 -938
rect 7272 -1002 7336 -938
rect 7352 -1002 7416 -938
rect 7432 -1002 7496 -938
rect 7512 -1002 7576 -938
rect 7592 -961 7656 -938
rect 7592 -1002 7650 -961
rect 7650 -1002 7656 -961
rect 7823 -62 7887 2
rect 7823 -142 7887 -78
rect 7823 -222 7887 -158
rect 7823 -302 7887 -238
rect 7823 -382 7887 -318
rect 7823 -462 7887 -398
rect 7823 -542 7887 -478
rect 7823 -622 7887 -558
rect 7823 -702 7887 -638
rect 7823 -782 7887 -718
rect 8429 -62 8493 2
rect 8429 -142 8493 -78
rect 8429 -222 8493 -158
rect 8429 -302 8493 -238
rect 8429 -382 8493 -318
rect 8429 -462 8493 -398
rect 8429 -542 8493 -478
rect 8429 -622 8493 -558
rect 8429 -702 8493 -638
rect 8429 -782 8493 -718
rect 9035 -62 9099 2
rect 9035 -142 9099 -78
rect 9035 -222 9099 -158
rect 9035 -302 9099 -238
rect 9035 -382 9099 -318
rect 9035 -462 9099 -398
rect 9035 -542 9099 -478
rect 9035 -622 9099 -558
rect 9035 -702 9099 -638
rect 9035 -782 9099 -718
rect 7926 -1002 7990 -938
rect 8006 -1002 8070 -938
rect 8086 -1002 8150 -938
rect 8166 -1002 8230 -938
rect 8246 -1002 8310 -938
rect 8326 -961 8390 -938
rect 8326 -1002 8384 -961
rect 8384 -1002 8390 -961
rect 8532 -961 8596 -938
rect 8532 -1002 8538 -961
rect 8538 -1002 8596 -961
rect 8612 -1002 8676 -938
rect 8692 -1002 8756 -938
rect 8772 -1002 8836 -938
rect 8852 -1002 8916 -938
rect 8932 -1002 8996 -938
rect 9161 -62 9225 2
rect 9161 -142 9225 -78
rect 9161 -222 9225 -158
rect 9161 -302 9225 -238
rect 9161 -382 9225 -318
rect 9161 -462 9225 -398
rect 9161 -542 9225 -478
rect 9161 -622 9225 -558
rect 9161 -702 9225 -638
rect 9161 -782 9225 -718
rect 9767 -62 9831 2
rect 9767 -142 9831 -78
rect 9767 -222 9831 -158
rect 9767 -302 9831 -238
rect 9767 -382 9831 -318
rect 9767 -462 9831 -398
rect 9767 -542 9831 -478
rect 9767 -622 9831 -558
rect 9767 -702 9831 -638
rect 9767 -782 9831 -718
rect 10373 -62 10437 2
rect 10373 -142 10437 -78
rect 10373 -222 10437 -158
rect 10373 -302 10437 -238
rect 10373 -382 10437 -318
rect 10373 -462 10437 -398
rect 10373 -542 10437 -478
rect 10373 -622 10437 -558
rect 10373 -702 10437 -638
rect 10373 -782 10437 -718
rect 10979 -62 11043 2
rect 10979 -142 11043 -78
rect 10979 -222 11043 -158
rect 10979 -302 11043 -238
rect 10979 -382 11043 -318
rect 10979 -462 11043 -398
rect 10979 -542 11043 -478
rect 10979 -622 11043 -558
rect 10979 -702 11043 -638
rect 10979 -782 11043 -718
rect 11585 -62 11649 2
rect 11585 -142 11649 -78
rect 11585 -222 11649 -158
rect 11585 -302 11649 -238
rect 11585 -382 11649 -318
rect 11585 -462 11649 -398
rect 11585 -542 11649 -478
rect 11585 -622 11649 -558
rect 11585 -702 11649 -638
rect 11585 -782 11649 -718
rect 9264 -1002 9328 -938
rect 9344 -1002 9408 -938
rect 9424 -1002 9488 -938
rect 9504 -1002 9568 -938
rect 9584 -1002 9648 -938
rect 9664 -961 9728 -938
rect 9664 -1002 9722 -961
rect 9722 -1002 9728 -961
rect 9870 -961 9934 -938
rect 9870 -1002 9876 -961
rect 9876 -1002 9934 -961
rect 9950 -1002 10014 -938
rect 10030 -1002 10094 -938
rect 10110 -1002 10174 -938
rect 10190 -1002 10254 -938
rect 10270 -1002 10334 -938
rect 10476 -1002 10540 -938
rect 10556 -1002 10620 -938
rect 10636 -1002 10700 -938
rect 10716 -1002 10780 -938
rect 10796 -1002 10860 -938
rect 10876 -961 10940 -938
rect 10876 -1002 10934 -961
rect 10934 -1002 10940 -961
rect 11082 -961 11146 -938
rect 11082 -1002 11088 -961
rect 11088 -1002 11146 -961
rect 11162 -1002 11226 -938
rect 11242 -1002 11306 -938
rect 11322 -1002 11386 -938
rect 11402 -1002 11466 -938
rect 11482 -1002 11546 -938
rect 11711 -62 11775 2
rect 11711 -142 11775 -78
rect 11711 -222 11775 -158
rect 11711 -302 11775 -238
rect 11711 -382 11775 -318
rect 11711 -462 11775 -398
rect 11711 -542 11775 -478
rect 11711 -622 11775 -558
rect 11711 -702 11775 -638
rect 11711 -782 11775 -718
rect 12317 -62 12381 2
rect 12317 -142 12381 -78
rect 12317 -222 12381 -158
rect 12317 -302 12381 -238
rect 12317 -382 12381 -318
rect 12317 -462 12381 -398
rect 12317 -542 12381 -478
rect 12317 -622 12381 -558
rect 12317 -702 12381 -638
rect 12317 -782 12381 -718
rect 11814 -961 11878 -938
rect 11814 -1002 11820 -961
rect 11820 -1002 11878 -961
rect 11894 -1002 11958 -938
rect 11974 -1002 12038 -938
rect 12054 -1002 12118 -938
rect 12134 -1002 12198 -938
rect 12214 -1002 12278 -938
rect 133 -1169 197 -1165
rect 133 -1225 137 -1169
rect 137 -1225 193 -1169
rect 193 -1225 197 -1169
rect 133 -1229 197 -1225
rect 482 -1250 546 -1186
rect 562 -1250 626 -1186
rect 642 -1250 706 -1186
rect 722 -1250 786 -1186
rect 802 -1250 866 -1186
rect 882 -1227 935 -1186
rect 935 -1227 946 -1186
rect 882 -1250 946 -1227
rect 1088 -1227 1099 -1186
rect 1099 -1227 1152 -1186
rect 1088 -1250 1152 -1227
rect 1168 -1250 1232 -1186
rect 1248 -1250 1312 -1186
rect 1328 -1250 1392 -1186
rect 1408 -1250 1472 -1186
rect 1488 -1250 1552 -1186
rect 1694 -1250 1758 -1186
rect 1774 -1250 1838 -1186
rect 1854 -1250 1918 -1186
rect 1934 -1250 1998 -1186
rect 2014 -1250 2078 -1186
rect 2094 -1227 2147 -1186
rect 2147 -1227 2158 -1186
rect 2094 -1250 2158 -1227
rect 2300 -1227 2311 -1186
rect 2311 -1227 2364 -1186
rect 2300 -1250 2364 -1227
rect 2380 -1250 2444 -1186
rect 2460 -1250 2524 -1186
rect 2540 -1250 2604 -1186
rect 2620 -1250 2684 -1186
rect 2700 -1250 2764 -1186
rect 2906 -1250 2970 -1186
rect 2986 -1250 3050 -1186
rect 3066 -1250 3130 -1186
rect 3146 -1250 3210 -1186
rect 3226 -1250 3290 -1186
rect 3306 -1227 3359 -1186
rect 3359 -1227 3370 -1186
rect 3306 -1250 3370 -1227
rect 3512 -1227 3523 -1186
rect 3523 -1227 3576 -1186
rect 3512 -1250 3576 -1227
rect 3592 -1250 3656 -1186
rect 3672 -1250 3736 -1186
rect 3752 -1250 3816 -1186
rect 3832 -1250 3896 -1186
rect 3912 -1250 3976 -1186
rect 4118 -1250 4182 -1186
rect 4198 -1250 4262 -1186
rect 4278 -1250 4342 -1186
rect 4358 -1250 4422 -1186
rect 4438 -1250 4502 -1186
rect 4518 -1227 4571 -1186
rect 4571 -1227 4582 -1186
rect 4518 -1250 4582 -1227
rect 4724 -1227 4735 -1186
rect 4735 -1227 4788 -1186
rect 4724 -1250 4788 -1227
rect 4804 -1250 4868 -1186
rect 4884 -1250 4948 -1186
rect 4964 -1250 5028 -1186
rect 5044 -1250 5108 -1186
rect 5124 -1250 5188 -1186
rect 221 -1430 285 -1426
rect 221 -1486 225 -1430
rect 225 -1486 281 -1430
rect 281 -1486 285 -1430
rect 221 -1490 285 -1486
rect 379 -1470 443 -1406
rect 379 -1550 443 -1486
rect 379 -1630 443 -1566
rect 139 -1672 203 -1668
rect 139 -1728 143 -1672
rect 143 -1728 199 -1672
rect 199 -1728 203 -1672
rect 139 -1732 203 -1728
rect 379 -1710 443 -1646
rect 379 -1790 443 -1726
rect 138 -1829 202 -1825
rect 138 -1885 142 -1829
rect 142 -1885 198 -1829
rect 198 -1885 202 -1829
rect 138 -1889 202 -1885
rect 379 -1870 443 -1806
rect 379 -1950 443 -1886
rect 138 -1999 202 -1995
rect 138 -2055 142 -1999
rect 142 -2055 198 -1999
rect 198 -2055 202 -1999
rect 138 -2059 202 -2055
rect 379 -2030 443 -1966
rect 379 -2110 443 -2046
rect 139 -2151 203 -2147
rect 139 -2207 143 -2151
rect 143 -2207 199 -2151
rect 199 -2207 203 -2151
rect 139 -2211 203 -2207
rect 379 -2190 443 -2126
rect 144 -2295 208 -2291
rect 144 -2351 148 -2295
rect 148 -2351 204 -2295
rect 204 -2351 208 -2295
rect 144 -2355 208 -2351
rect 985 -1470 1049 -1406
rect 985 -1550 1049 -1486
rect 985 -1630 1049 -1566
rect 985 -1710 1049 -1646
rect 985 -1790 1049 -1726
rect 985 -1870 1049 -1806
rect 985 -1950 1049 -1886
rect 985 -2030 1049 -1966
rect 985 -2110 1049 -2046
rect 985 -2190 1049 -2126
rect 1591 -1470 1655 -1406
rect 1591 -1550 1655 -1486
rect 1591 -1630 1655 -1566
rect 1591 -1710 1655 -1646
rect 1591 -1790 1655 -1726
rect 1591 -1870 1655 -1806
rect 1591 -1950 1655 -1886
rect 1591 -2030 1655 -1966
rect 1591 -2110 1655 -2046
rect 1591 -2190 1655 -2126
rect 2197 -1470 2261 -1406
rect 2197 -1550 2261 -1486
rect 2197 -1630 2261 -1566
rect 2197 -1710 2261 -1646
rect 2197 -1790 2261 -1726
rect 2197 -1870 2261 -1806
rect 2197 -1950 2261 -1886
rect 2197 -2030 2261 -1966
rect 2197 -2110 2261 -2046
rect 2197 -2190 2261 -2126
rect 2803 -1470 2867 -1406
rect 2803 -1550 2867 -1486
rect 2803 -1630 2867 -1566
rect 2803 -1710 2867 -1646
rect 2803 -1790 2867 -1726
rect 2803 -1870 2867 -1806
rect 2803 -1950 2867 -1886
rect 2803 -2030 2867 -1966
rect 2803 -2110 2867 -2046
rect 2803 -2190 2867 -2126
rect 3409 -1470 3473 -1406
rect 3409 -1550 3473 -1486
rect 3409 -1630 3473 -1566
rect 3409 -1710 3473 -1646
rect 3409 -1790 3473 -1726
rect 3409 -1870 3473 -1806
rect 3409 -1950 3473 -1886
rect 3409 -2030 3473 -1966
rect 3409 -2110 3473 -2046
rect 3409 -2190 3473 -2126
rect 4015 -1470 4079 -1406
rect 4015 -1550 4079 -1486
rect 4015 -1630 4079 -1566
rect 4015 -1710 4079 -1646
rect 4015 -1790 4079 -1726
rect 4015 -1870 4079 -1806
rect 4015 -1950 4079 -1886
rect 4015 -2030 4079 -1966
rect 4015 -2110 4079 -2046
rect 4015 -2190 4079 -2126
rect 4621 -1470 4685 -1406
rect 4621 -1550 4685 -1486
rect 4621 -1630 4685 -1566
rect 4621 -1710 4685 -1646
rect 4621 -1790 4685 -1726
rect 4621 -1870 4685 -1806
rect 4621 -1950 4685 -1886
rect 4621 -2030 4685 -1966
rect 4621 -2110 4685 -2046
rect 4621 -2190 4685 -2126
rect 5227 -1470 5291 -1406
rect 5227 -1550 5291 -1486
rect 5227 -1630 5291 -1566
rect 5227 -1710 5291 -1646
rect 5227 -1790 5291 -1726
rect 5227 -1870 5291 -1806
rect 5227 -1950 5291 -1886
rect 5227 -2030 5291 -1966
rect 5227 -2110 5291 -2046
rect 5227 -2190 5291 -2126
rect 5456 -1224 5467 -1183
rect 5467 -1224 5520 -1183
rect 5456 -1247 5520 -1224
rect 5536 -1247 5600 -1183
rect 5616 -1247 5680 -1183
rect 5696 -1247 5760 -1183
rect 5776 -1247 5840 -1183
rect 5856 -1247 5920 -1183
rect 5353 -1467 5417 -1403
rect 5353 -1547 5417 -1483
rect 5353 -1627 5417 -1563
rect 5353 -1707 5417 -1643
rect 5353 -1787 5417 -1723
rect 5353 -1867 5417 -1803
rect 5353 -1947 5417 -1883
rect 5353 -2027 5417 -1963
rect 5353 -2107 5417 -2043
rect 5353 -2187 5417 -2123
rect 6289 -1206 6353 -1202
rect 6289 -1262 6293 -1206
rect 6293 -1262 6349 -1206
rect 6349 -1262 6353 -1206
rect 6289 -1266 6353 -1262
rect 6432 -1206 6496 -1202
rect 6432 -1262 6436 -1206
rect 6436 -1262 6492 -1206
rect 6492 -1262 6496 -1206
rect 6432 -1266 6496 -1262
rect 6552 -1206 6616 -1202
rect 6552 -1262 6556 -1206
rect 6556 -1262 6612 -1206
rect 6612 -1262 6616 -1206
rect 6552 -1266 6616 -1262
rect 6842 -1169 6906 -1165
rect 6842 -1225 6846 -1169
rect 6846 -1225 6902 -1169
rect 6902 -1225 6906 -1169
rect 6842 -1229 6906 -1225
rect 7191 -1250 7255 -1186
rect 7271 -1250 7335 -1186
rect 7351 -1250 7415 -1186
rect 7431 -1250 7495 -1186
rect 7511 -1250 7575 -1186
rect 7591 -1227 7644 -1186
rect 7644 -1227 7655 -1186
rect 7591 -1250 7655 -1227
rect 7797 -1227 7808 -1186
rect 7808 -1227 7861 -1186
rect 7797 -1250 7861 -1227
rect 7877 -1250 7941 -1186
rect 7957 -1250 8021 -1186
rect 8037 -1250 8101 -1186
rect 8117 -1250 8181 -1186
rect 8197 -1250 8261 -1186
rect 8403 -1250 8467 -1186
rect 8483 -1250 8547 -1186
rect 8563 -1250 8627 -1186
rect 8643 -1250 8707 -1186
rect 8723 -1250 8787 -1186
rect 8803 -1227 8856 -1186
rect 8856 -1227 8867 -1186
rect 8803 -1250 8867 -1227
rect 9009 -1227 9020 -1186
rect 9020 -1227 9073 -1186
rect 9009 -1250 9073 -1227
rect 9089 -1250 9153 -1186
rect 9169 -1250 9233 -1186
rect 9249 -1250 9313 -1186
rect 9329 -1250 9393 -1186
rect 9409 -1250 9473 -1186
rect 9615 -1250 9679 -1186
rect 9695 -1250 9759 -1186
rect 9775 -1250 9839 -1186
rect 9855 -1250 9919 -1186
rect 9935 -1250 9999 -1186
rect 10015 -1227 10068 -1186
rect 10068 -1227 10079 -1186
rect 10015 -1250 10079 -1227
rect 10221 -1227 10232 -1186
rect 10232 -1227 10285 -1186
rect 10221 -1250 10285 -1227
rect 10301 -1250 10365 -1186
rect 10381 -1250 10445 -1186
rect 10461 -1250 10525 -1186
rect 10541 -1250 10605 -1186
rect 10621 -1250 10685 -1186
rect 10827 -1250 10891 -1186
rect 10907 -1250 10971 -1186
rect 10987 -1250 11051 -1186
rect 11067 -1250 11131 -1186
rect 11147 -1250 11211 -1186
rect 11227 -1227 11280 -1186
rect 11280 -1227 11291 -1186
rect 11227 -1250 11291 -1227
rect 11433 -1227 11444 -1186
rect 11444 -1227 11497 -1186
rect 11433 -1250 11497 -1227
rect 11513 -1250 11577 -1186
rect 11593 -1250 11657 -1186
rect 11673 -1250 11737 -1186
rect 11753 -1250 11817 -1186
rect 11833 -1250 11897 -1186
rect 5959 -1467 6023 -1403
rect 5959 -1547 6023 -1483
rect 6930 -1430 6994 -1426
rect 6930 -1486 6934 -1430
rect 6934 -1486 6990 -1430
rect 6990 -1486 6994 -1430
rect 6930 -1490 6994 -1486
rect 7088 -1470 7152 -1406
rect 5959 -1627 6023 -1563
rect 5959 -1707 6023 -1643
rect 7088 -1550 7152 -1486
rect 7088 -1630 7152 -1566
rect 5959 -1787 6023 -1723
rect 5959 -1867 6023 -1803
rect 6848 -1672 6912 -1668
rect 6848 -1728 6852 -1672
rect 6852 -1728 6908 -1672
rect 6908 -1728 6912 -1672
rect 6848 -1732 6912 -1728
rect 7088 -1710 7152 -1646
rect 6295 -1752 6359 -1748
rect 6295 -1808 6299 -1752
rect 6299 -1808 6355 -1752
rect 6355 -1808 6359 -1752
rect 6295 -1812 6359 -1808
rect 6439 -1751 6503 -1747
rect 6439 -1807 6443 -1751
rect 6443 -1807 6499 -1751
rect 6499 -1807 6503 -1751
rect 6439 -1811 6503 -1807
rect 6570 -1752 6634 -1748
rect 6570 -1808 6574 -1752
rect 6574 -1808 6630 -1752
rect 6630 -1808 6634 -1752
rect 6570 -1812 6634 -1808
rect 7088 -1790 7152 -1726
rect 5959 -1947 6023 -1883
rect 5959 -2027 6023 -1963
rect 6425 -1901 6489 -1897
rect 6425 -1957 6429 -1901
rect 6429 -1957 6485 -1901
rect 6485 -1957 6489 -1901
rect 6425 -1961 6489 -1957
rect 6847 -1829 6911 -1825
rect 6847 -1885 6851 -1829
rect 6851 -1885 6907 -1829
rect 6907 -1885 6911 -1829
rect 6847 -1889 6911 -1885
rect 7088 -1870 7152 -1806
rect 7088 -1950 7152 -1886
rect 5959 -2107 6023 -2043
rect 6847 -1999 6911 -1995
rect 6847 -2055 6851 -1999
rect 6851 -2055 6907 -1999
rect 6907 -2055 6911 -1999
rect 6847 -2059 6911 -2055
rect 7088 -2030 7152 -1966
rect 5959 -2187 6023 -2123
rect 6425 -2097 6489 -2093
rect 6425 -2153 6429 -2097
rect 6429 -2153 6485 -2097
rect 6485 -2153 6489 -2097
rect 6425 -2157 6489 -2153
rect 7088 -2110 7152 -2046
rect 6848 -2151 6912 -2147
rect 6848 -2207 6852 -2151
rect 6852 -2207 6908 -2151
rect 6908 -2207 6912 -2151
rect 6848 -2211 6912 -2207
rect 7088 -2190 7152 -2126
rect 6425 -2272 6489 -2268
rect 6425 -2328 6429 -2272
rect 6429 -2328 6485 -2272
rect 6485 -2328 6489 -2272
rect 6425 -2332 6489 -2328
rect 482 -2351 546 -2346
rect 482 -2407 485 -2351
rect 485 -2407 541 -2351
rect 541 -2407 546 -2351
rect 482 -2410 546 -2407
rect 562 -2351 626 -2346
rect 562 -2407 565 -2351
rect 565 -2407 621 -2351
rect 621 -2407 626 -2351
rect 562 -2410 626 -2407
rect 642 -2351 706 -2346
rect 642 -2407 645 -2351
rect 645 -2407 701 -2351
rect 701 -2407 706 -2351
rect 642 -2410 706 -2407
rect 722 -2351 786 -2346
rect 722 -2407 725 -2351
rect 725 -2407 781 -2351
rect 781 -2407 786 -2351
rect 722 -2410 786 -2407
rect 802 -2351 866 -2346
rect 802 -2407 805 -2351
rect 805 -2407 861 -2351
rect 861 -2407 866 -2351
rect 802 -2410 866 -2407
rect 882 -2351 946 -2346
rect 882 -2407 885 -2351
rect 885 -2407 941 -2351
rect 941 -2407 946 -2351
rect 882 -2410 946 -2407
rect 1088 -2351 1152 -2346
rect 1088 -2407 1093 -2351
rect 1093 -2407 1149 -2351
rect 1149 -2407 1152 -2351
rect 1088 -2410 1152 -2407
rect 1168 -2351 1232 -2346
rect 1168 -2407 1173 -2351
rect 1173 -2407 1229 -2351
rect 1229 -2407 1232 -2351
rect 1168 -2410 1232 -2407
rect 1248 -2351 1312 -2346
rect 1248 -2407 1253 -2351
rect 1253 -2407 1309 -2351
rect 1309 -2407 1312 -2351
rect 1248 -2410 1312 -2407
rect 1328 -2351 1392 -2346
rect 1328 -2407 1333 -2351
rect 1333 -2407 1389 -2351
rect 1389 -2407 1392 -2351
rect 1328 -2410 1392 -2407
rect 1408 -2351 1472 -2346
rect 1408 -2407 1413 -2351
rect 1413 -2407 1469 -2351
rect 1469 -2407 1472 -2351
rect 1408 -2410 1472 -2407
rect 1488 -2351 1552 -2346
rect 1488 -2407 1493 -2351
rect 1493 -2407 1549 -2351
rect 1549 -2407 1552 -2351
rect 1488 -2410 1552 -2407
rect 1694 -2351 1758 -2346
rect 1694 -2407 1697 -2351
rect 1697 -2407 1753 -2351
rect 1753 -2407 1758 -2351
rect 1694 -2410 1758 -2407
rect 1774 -2351 1838 -2346
rect 1774 -2407 1777 -2351
rect 1777 -2407 1833 -2351
rect 1833 -2407 1838 -2351
rect 1774 -2410 1838 -2407
rect 1854 -2351 1918 -2346
rect 1854 -2407 1857 -2351
rect 1857 -2407 1913 -2351
rect 1913 -2407 1918 -2351
rect 1854 -2410 1918 -2407
rect 1934 -2351 1998 -2346
rect 1934 -2407 1937 -2351
rect 1937 -2407 1993 -2351
rect 1993 -2407 1998 -2351
rect 1934 -2410 1998 -2407
rect 2014 -2351 2078 -2346
rect 2014 -2407 2017 -2351
rect 2017 -2407 2073 -2351
rect 2073 -2407 2078 -2351
rect 2014 -2410 2078 -2407
rect 2094 -2351 2158 -2346
rect 2094 -2407 2097 -2351
rect 2097 -2407 2153 -2351
rect 2153 -2407 2158 -2351
rect 2094 -2410 2158 -2407
rect 2300 -2351 2364 -2346
rect 2300 -2407 2305 -2351
rect 2305 -2407 2361 -2351
rect 2361 -2407 2364 -2351
rect 2300 -2410 2364 -2407
rect 2380 -2351 2444 -2346
rect 2380 -2407 2385 -2351
rect 2385 -2407 2441 -2351
rect 2441 -2407 2444 -2351
rect 2380 -2410 2444 -2407
rect 2460 -2351 2524 -2346
rect 2460 -2407 2465 -2351
rect 2465 -2407 2521 -2351
rect 2521 -2407 2524 -2351
rect 2460 -2410 2524 -2407
rect 2540 -2351 2604 -2346
rect 2540 -2407 2545 -2351
rect 2545 -2407 2601 -2351
rect 2601 -2407 2604 -2351
rect 2540 -2410 2604 -2407
rect 2620 -2351 2684 -2346
rect 2620 -2407 2625 -2351
rect 2625 -2407 2681 -2351
rect 2681 -2407 2684 -2351
rect 2620 -2410 2684 -2407
rect 2700 -2351 2764 -2346
rect 2700 -2407 2705 -2351
rect 2705 -2407 2761 -2351
rect 2761 -2407 2764 -2351
rect 2700 -2410 2764 -2407
rect 2906 -2351 2970 -2346
rect 2906 -2407 2909 -2351
rect 2909 -2407 2965 -2351
rect 2965 -2407 2970 -2351
rect 2906 -2410 2970 -2407
rect 2986 -2351 3050 -2346
rect 2986 -2407 2989 -2351
rect 2989 -2407 3045 -2351
rect 3045 -2407 3050 -2351
rect 2986 -2410 3050 -2407
rect 3066 -2351 3130 -2346
rect 3066 -2407 3069 -2351
rect 3069 -2407 3125 -2351
rect 3125 -2407 3130 -2351
rect 3066 -2410 3130 -2407
rect 3146 -2351 3210 -2346
rect 3146 -2407 3149 -2351
rect 3149 -2407 3205 -2351
rect 3205 -2407 3210 -2351
rect 3146 -2410 3210 -2407
rect 3226 -2351 3290 -2346
rect 3226 -2407 3229 -2351
rect 3229 -2407 3285 -2351
rect 3285 -2407 3290 -2351
rect 3226 -2410 3290 -2407
rect 3306 -2351 3370 -2346
rect 3306 -2407 3309 -2351
rect 3309 -2407 3365 -2351
rect 3365 -2407 3370 -2351
rect 3306 -2410 3370 -2407
rect 3512 -2351 3576 -2346
rect 3512 -2407 3517 -2351
rect 3517 -2407 3573 -2351
rect 3573 -2407 3576 -2351
rect 3512 -2410 3576 -2407
rect 3592 -2351 3656 -2346
rect 3592 -2407 3597 -2351
rect 3597 -2407 3653 -2351
rect 3653 -2407 3656 -2351
rect 3592 -2410 3656 -2407
rect 3672 -2351 3736 -2346
rect 3672 -2407 3677 -2351
rect 3677 -2407 3733 -2351
rect 3733 -2407 3736 -2351
rect 3672 -2410 3736 -2407
rect 3752 -2351 3816 -2346
rect 3752 -2407 3757 -2351
rect 3757 -2407 3813 -2351
rect 3813 -2407 3816 -2351
rect 3752 -2410 3816 -2407
rect 3832 -2351 3896 -2346
rect 3832 -2407 3837 -2351
rect 3837 -2407 3893 -2351
rect 3893 -2407 3896 -2351
rect 3832 -2410 3896 -2407
rect 3912 -2351 3976 -2346
rect 3912 -2407 3917 -2351
rect 3917 -2407 3973 -2351
rect 3973 -2407 3976 -2351
rect 3912 -2410 3976 -2407
rect 4118 -2351 4182 -2346
rect 4118 -2407 4121 -2351
rect 4121 -2407 4177 -2351
rect 4177 -2407 4182 -2351
rect 4118 -2410 4182 -2407
rect 4198 -2351 4262 -2346
rect 4198 -2407 4201 -2351
rect 4201 -2407 4257 -2351
rect 4257 -2407 4262 -2351
rect 4198 -2410 4262 -2407
rect 4278 -2351 4342 -2346
rect 4278 -2407 4281 -2351
rect 4281 -2407 4337 -2351
rect 4337 -2407 4342 -2351
rect 4278 -2410 4342 -2407
rect 4358 -2351 4422 -2346
rect 4358 -2407 4361 -2351
rect 4361 -2407 4417 -2351
rect 4417 -2407 4422 -2351
rect 4358 -2410 4422 -2407
rect 4438 -2351 4502 -2346
rect 4438 -2407 4441 -2351
rect 4441 -2407 4497 -2351
rect 4497 -2407 4502 -2351
rect 4438 -2410 4502 -2407
rect 4518 -2351 4582 -2346
rect 4518 -2407 4521 -2351
rect 4521 -2407 4577 -2351
rect 4577 -2407 4582 -2351
rect 4518 -2410 4582 -2407
rect 4724 -2351 4788 -2346
rect 4724 -2407 4729 -2351
rect 4729 -2407 4785 -2351
rect 4785 -2407 4788 -2351
rect 4724 -2410 4788 -2407
rect 4804 -2351 4868 -2346
rect 4804 -2407 4809 -2351
rect 4809 -2407 4865 -2351
rect 4865 -2407 4868 -2351
rect 4804 -2410 4868 -2407
rect 4884 -2351 4948 -2346
rect 4884 -2407 4889 -2351
rect 4889 -2407 4945 -2351
rect 4945 -2407 4948 -2351
rect 4884 -2410 4948 -2407
rect 4964 -2351 5028 -2346
rect 4964 -2407 4969 -2351
rect 4969 -2407 5025 -2351
rect 5025 -2407 5028 -2351
rect 4964 -2410 5028 -2407
rect 5044 -2351 5108 -2346
rect 5044 -2407 5049 -2351
rect 5049 -2407 5105 -2351
rect 5105 -2407 5108 -2351
rect 5044 -2410 5108 -2407
rect 5124 -2351 5188 -2346
rect 5124 -2407 5129 -2351
rect 5129 -2407 5185 -2351
rect 5185 -2407 5188 -2351
rect 5124 -2410 5188 -2407
rect 5456 -2348 5520 -2343
rect 5456 -2404 5461 -2348
rect 5461 -2404 5517 -2348
rect 5517 -2404 5520 -2348
rect 5456 -2407 5520 -2404
rect 5536 -2348 5600 -2343
rect 5536 -2404 5541 -2348
rect 5541 -2404 5597 -2348
rect 5597 -2404 5600 -2348
rect 5536 -2407 5600 -2404
rect 5616 -2348 5680 -2343
rect 5616 -2404 5621 -2348
rect 5621 -2404 5677 -2348
rect 5677 -2404 5680 -2348
rect 5616 -2407 5680 -2404
rect 5696 -2348 5760 -2343
rect 5696 -2404 5701 -2348
rect 5701 -2404 5757 -2348
rect 5757 -2404 5760 -2348
rect 5696 -2407 5760 -2404
rect 5776 -2348 5840 -2343
rect 5776 -2404 5781 -2348
rect 5781 -2404 5837 -2348
rect 5837 -2404 5840 -2348
rect 5776 -2407 5840 -2404
rect 5856 -2348 5920 -2343
rect 5856 -2404 5861 -2348
rect 5861 -2404 5917 -2348
rect 5917 -2404 5920 -2348
rect 5856 -2407 5920 -2404
rect 5953 -2357 6017 -2353
rect 5953 -2413 5957 -2357
rect 5957 -2413 6013 -2357
rect 6013 -2413 6017 -2357
rect 5953 -2417 6017 -2413
rect 6853 -2295 6917 -2291
rect 6853 -2351 6857 -2295
rect 6857 -2351 6913 -2295
rect 6913 -2351 6917 -2295
rect 6853 -2355 6917 -2351
rect 7694 -1470 7758 -1406
rect 7694 -1550 7758 -1486
rect 7694 -1630 7758 -1566
rect 7694 -1710 7758 -1646
rect 7694 -1790 7758 -1726
rect 7694 -1870 7758 -1806
rect 7694 -1950 7758 -1886
rect 7694 -2030 7758 -1966
rect 7694 -2110 7758 -2046
rect 7694 -2190 7758 -2126
rect 8300 -1470 8364 -1406
rect 8300 -1550 8364 -1486
rect 8300 -1630 8364 -1566
rect 8300 -1710 8364 -1646
rect 8300 -1790 8364 -1726
rect 8300 -1870 8364 -1806
rect 8300 -1950 8364 -1886
rect 8300 -2030 8364 -1966
rect 8300 -2110 8364 -2046
rect 8300 -2190 8364 -2126
rect 8906 -1470 8970 -1406
rect 8906 -1550 8970 -1486
rect 8906 -1630 8970 -1566
rect 8906 -1710 8970 -1646
rect 8906 -1790 8970 -1726
rect 8906 -1870 8970 -1806
rect 8906 -1950 8970 -1886
rect 8906 -2030 8970 -1966
rect 8906 -2110 8970 -2046
rect 8906 -2190 8970 -2126
rect 9512 -1470 9576 -1406
rect 9512 -1550 9576 -1486
rect 9512 -1630 9576 -1566
rect 9512 -1710 9576 -1646
rect 9512 -1790 9576 -1726
rect 9512 -1870 9576 -1806
rect 9512 -1950 9576 -1886
rect 9512 -2030 9576 -1966
rect 9512 -2110 9576 -2046
rect 9512 -2190 9576 -2126
rect 10118 -1470 10182 -1406
rect 10118 -1550 10182 -1486
rect 10118 -1630 10182 -1566
rect 10118 -1710 10182 -1646
rect 10118 -1790 10182 -1726
rect 10118 -1870 10182 -1806
rect 10118 -1950 10182 -1886
rect 10118 -2030 10182 -1966
rect 10118 -2110 10182 -2046
rect 10118 -2190 10182 -2126
rect 10724 -1470 10788 -1406
rect 10724 -1550 10788 -1486
rect 10724 -1630 10788 -1566
rect 10724 -1710 10788 -1646
rect 10724 -1790 10788 -1726
rect 10724 -1870 10788 -1806
rect 10724 -1950 10788 -1886
rect 10724 -2030 10788 -1966
rect 10724 -2110 10788 -2046
rect 10724 -2190 10788 -2126
rect 11330 -1470 11394 -1406
rect 11330 -1550 11394 -1486
rect 11330 -1630 11394 -1566
rect 11330 -1710 11394 -1646
rect 11330 -1790 11394 -1726
rect 11330 -1870 11394 -1806
rect 11330 -1950 11394 -1886
rect 11330 -2030 11394 -1966
rect 11330 -2110 11394 -2046
rect 11330 -2190 11394 -2126
rect 11936 -1470 12000 -1406
rect 11936 -1550 12000 -1486
rect 11936 -1630 12000 -1566
rect 11936 -1710 12000 -1646
rect 11936 -1790 12000 -1726
rect 11936 -1870 12000 -1806
rect 11936 -1950 12000 -1886
rect 11936 -2030 12000 -1966
rect 11936 -2110 12000 -2046
rect 11936 -2190 12000 -2126
rect 12165 -1224 12176 -1183
rect 12176 -1224 12229 -1183
rect 12165 -1247 12229 -1224
rect 12245 -1247 12309 -1183
rect 12325 -1247 12389 -1183
rect 12405 -1247 12469 -1183
rect 12485 -1247 12549 -1183
rect 12565 -1247 12629 -1183
rect 12062 -1467 12126 -1403
rect 12062 -1547 12126 -1483
rect 12062 -1627 12126 -1563
rect 12062 -1707 12126 -1643
rect 12062 -1787 12126 -1723
rect 12062 -1867 12126 -1803
rect 12062 -1947 12126 -1883
rect 12062 -2027 12126 -1963
rect 12062 -2107 12126 -2043
rect 12062 -2187 12126 -2123
rect 12998 -1206 13062 -1202
rect 12998 -1262 13002 -1206
rect 13002 -1262 13058 -1206
rect 13058 -1262 13062 -1206
rect 12998 -1266 13062 -1262
rect 13141 -1206 13205 -1202
rect 13141 -1262 13145 -1206
rect 13145 -1262 13201 -1206
rect 13201 -1262 13205 -1206
rect 13141 -1266 13205 -1262
rect 13261 -1206 13325 -1202
rect 13261 -1262 13265 -1206
rect 13265 -1262 13321 -1206
rect 13321 -1262 13325 -1206
rect 13261 -1266 13325 -1262
rect 12668 -1467 12732 -1403
rect 12668 -1547 12732 -1483
rect 12668 -1627 12732 -1563
rect 12668 -1707 12732 -1643
rect 12668 -1787 12732 -1723
rect 12668 -1867 12732 -1803
rect 13004 -1752 13068 -1748
rect 13004 -1808 13008 -1752
rect 13008 -1808 13064 -1752
rect 13064 -1808 13068 -1752
rect 13004 -1812 13068 -1808
rect 13148 -1751 13212 -1747
rect 13148 -1807 13152 -1751
rect 13152 -1807 13208 -1751
rect 13208 -1807 13212 -1751
rect 13148 -1811 13212 -1807
rect 13279 -1752 13343 -1748
rect 13279 -1808 13283 -1752
rect 13283 -1808 13339 -1752
rect 13339 -1808 13343 -1752
rect 13279 -1812 13343 -1808
rect 12668 -1947 12732 -1883
rect 12668 -2027 12732 -1963
rect 12668 -2107 12732 -2043
rect 12668 -2187 12732 -2123
rect 7191 -2351 7255 -2346
rect 7191 -2407 7194 -2351
rect 7194 -2407 7250 -2351
rect 7250 -2407 7255 -2351
rect 7191 -2410 7255 -2407
rect 7271 -2351 7335 -2346
rect 7271 -2407 7274 -2351
rect 7274 -2407 7330 -2351
rect 7330 -2407 7335 -2351
rect 7271 -2410 7335 -2407
rect 7351 -2351 7415 -2346
rect 7351 -2407 7354 -2351
rect 7354 -2407 7410 -2351
rect 7410 -2407 7415 -2351
rect 7351 -2410 7415 -2407
rect 7431 -2351 7495 -2346
rect 7431 -2407 7434 -2351
rect 7434 -2407 7490 -2351
rect 7490 -2407 7495 -2351
rect 7431 -2410 7495 -2407
rect 7511 -2351 7575 -2346
rect 7511 -2407 7514 -2351
rect 7514 -2407 7570 -2351
rect 7570 -2407 7575 -2351
rect 7511 -2410 7575 -2407
rect 7591 -2351 7655 -2346
rect 7591 -2407 7594 -2351
rect 7594 -2407 7650 -2351
rect 7650 -2407 7655 -2351
rect 7591 -2410 7655 -2407
rect 7797 -2351 7861 -2346
rect 7797 -2407 7802 -2351
rect 7802 -2407 7858 -2351
rect 7858 -2407 7861 -2351
rect 7797 -2410 7861 -2407
rect 7877 -2351 7941 -2346
rect 7877 -2407 7882 -2351
rect 7882 -2407 7938 -2351
rect 7938 -2407 7941 -2351
rect 7877 -2410 7941 -2407
rect 7957 -2351 8021 -2346
rect 7957 -2407 7962 -2351
rect 7962 -2407 8018 -2351
rect 8018 -2407 8021 -2351
rect 7957 -2410 8021 -2407
rect 8037 -2351 8101 -2346
rect 8037 -2407 8042 -2351
rect 8042 -2407 8098 -2351
rect 8098 -2407 8101 -2351
rect 8037 -2410 8101 -2407
rect 8117 -2351 8181 -2346
rect 8117 -2407 8122 -2351
rect 8122 -2407 8178 -2351
rect 8178 -2407 8181 -2351
rect 8117 -2410 8181 -2407
rect 8197 -2351 8261 -2346
rect 8197 -2407 8202 -2351
rect 8202 -2407 8258 -2351
rect 8258 -2407 8261 -2351
rect 8197 -2410 8261 -2407
rect 8403 -2351 8467 -2346
rect 8403 -2407 8406 -2351
rect 8406 -2407 8462 -2351
rect 8462 -2407 8467 -2351
rect 8403 -2410 8467 -2407
rect 8483 -2351 8547 -2346
rect 8483 -2407 8486 -2351
rect 8486 -2407 8542 -2351
rect 8542 -2407 8547 -2351
rect 8483 -2410 8547 -2407
rect 8563 -2351 8627 -2346
rect 8563 -2407 8566 -2351
rect 8566 -2407 8622 -2351
rect 8622 -2407 8627 -2351
rect 8563 -2410 8627 -2407
rect 8643 -2351 8707 -2346
rect 8643 -2407 8646 -2351
rect 8646 -2407 8702 -2351
rect 8702 -2407 8707 -2351
rect 8643 -2410 8707 -2407
rect 8723 -2351 8787 -2346
rect 8723 -2407 8726 -2351
rect 8726 -2407 8782 -2351
rect 8782 -2407 8787 -2351
rect 8723 -2410 8787 -2407
rect 8803 -2351 8867 -2346
rect 8803 -2407 8806 -2351
rect 8806 -2407 8862 -2351
rect 8862 -2407 8867 -2351
rect 8803 -2410 8867 -2407
rect 9009 -2351 9073 -2346
rect 9009 -2407 9014 -2351
rect 9014 -2407 9070 -2351
rect 9070 -2407 9073 -2351
rect 9009 -2410 9073 -2407
rect 9089 -2351 9153 -2346
rect 9089 -2407 9094 -2351
rect 9094 -2407 9150 -2351
rect 9150 -2407 9153 -2351
rect 9089 -2410 9153 -2407
rect 9169 -2351 9233 -2346
rect 9169 -2407 9174 -2351
rect 9174 -2407 9230 -2351
rect 9230 -2407 9233 -2351
rect 9169 -2410 9233 -2407
rect 9249 -2351 9313 -2346
rect 9249 -2407 9254 -2351
rect 9254 -2407 9310 -2351
rect 9310 -2407 9313 -2351
rect 9249 -2410 9313 -2407
rect 9329 -2351 9393 -2346
rect 9329 -2407 9334 -2351
rect 9334 -2407 9390 -2351
rect 9390 -2407 9393 -2351
rect 9329 -2410 9393 -2407
rect 9409 -2351 9473 -2346
rect 9409 -2407 9414 -2351
rect 9414 -2407 9470 -2351
rect 9470 -2407 9473 -2351
rect 9409 -2410 9473 -2407
rect 9615 -2351 9679 -2346
rect 9615 -2407 9618 -2351
rect 9618 -2407 9674 -2351
rect 9674 -2407 9679 -2351
rect 9615 -2410 9679 -2407
rect 9695 -2351 9759 -2346
rect 9695 -2407 9698 -2351
rect 9698 -2407 9754 -2351
rect 9754 -2407 9759 -2351
rect 9695 -2410 9759 -2407
rect 9775 -2351 9839 -2346
rect 9775 -2407 9778 -2351
rect 9778 -2407 9834 -2351
rect 9834 -2407 9839 -2351
rect 9775 -2410 9839 -2407
rect 9855 -2351 9919 -2346
rect 9855 -2407 9858 -2351
rect 9858 -2407 9914 -2351
rect 9914 -2407 9919 -2351
rect 9855 -2410 9919 -2407
rect 9935 -2351 9999 -2346
rect 9935 -2407 9938 -2351
rect 9938 -2407 9994 -2351
rect 9994 -2407 9999 -2351
rect 9935 -2410 9999 -2407
rect 10015 -2351 10079 -2346
rect 10015 -2407 10018 -2351
rect 10018 -2407 10074 -2351
rect 10074 -2407 10079 -2351
rect 10015 -2410 10079 -2407
rect 10221 -2351 10285 -2346
rect 10221 -2407 10226 -2351
rect 10226 -2407 10282 -2351
rect 10282 -2407 10285 -2351
rect 10221 -2410 10285 -2407
rect 10301 -2351 10365 -2346
rect 10301 -2407 10306 -2351
rect 10306 -2407 10362 -2351
rect 10362 -2407 10365 -2351
rect 10301 -2410 10365 -2407
rect 10381 -2351 10445 -2346
rect 10381 -2407 10386 -2351
rect 10386 -2407 10442 -2351
rect 10442 -2407 10445 -2351
rect 10381 -2410 10445 -2407
rect 10461 -2351 10525 -2346
rect 10461 -2407 10466 -2351
rect 10466 -2407 10522 -2351
rect 10522 -2407 10525 -2351
rect 10461 -2410 10525 -2407
rect 10541 -2351 10605 -2346
rect 10541 -2407 10546 -2351
rect 10546 -2407 10602 -2351
rect 10602 -2407 10605 -2351
rect 10541 -2410 10605 -2407
rect 10621 -2351 10685 -2346
rect 10621 -2407 10626 -2351
rect 10626 -2407 10682 -2351
rect 10682 -2407 10685 -2351
rect 10621 -2410 10685 -2407
rect 10827 -2351 10891 -2346
rect 10827 -2407 10830 -2351
rect 10830 -2407 10886 -2351
rect 10886 -2407 10891 -2351
rect 10827 -2410 10891 -2407
rect 10907 -2351 10971 -2346
rect 10907 -2407 10910 -2351
rect 10910 -2407 10966 -2351
rect 10966 -2407 10971 -2351
rect 10907 -2410 10971 -2407
rect 10987 -2351 11051 -2346
rect 10987 -2407 10990 -2351
rect 10990 -2407 11046 -2351
rect 11046 -2407 11051 -2351
rect 10987 -2410 11051 -2407
rect 11067 -2351 11131 -2346
rect 11067 -2407 11070 -2351
rect 11070 -2407 11126 -2351
rect 11126 -2407 11131 -2351
rect 11067 -2410 11131 -2407
rect 11147 -2351 11211 -2346
rect 11147 -2407 11150 -2351
rect 11150 -2407 11206 -2351
rect 11206 -2407 11211 -2351
rect 11147 -2410 11211 -2407
rect 11227 -2351 11291 -2346
rect 11227 -2407 11230 -2351
rect 11230 -2407 11286 -2351
rect 11286 -2407 11291 -2351
rect 11227 -2410 11291 -2407
rect 11433 -2351 11497 -2346
rect 11433 -2407 11438 -2351
rect 11438 -2407 11494 -2351
rect 11494 -2407 11497 -2351
rect 11433 -2410 11497 -2407
rect 11513 -2351 11577 -2346
rect 11513 -2407 11518 -2351
rect 11518 -2407 11574 -2351
rect 11574 -2407 11577 -2351
rect 11513 -2410 11577 -2407
rect 11593 -2351 11657 -2346
rect 11593 -2407 11598 -2351
rect 11598 -2407 11654 -2351
rect 11654 -2407 11657 -2351
rect 11593 -2410 11657 -2407
rect 11673 -2351 11737 -2346
rect 11673 -2407 11678 -2351
rect 11678 -2407 11734 -2351
rect 11734 -2407 11737 -2351
rect 11673 -2410 11737 -2407
rect 11753 -2351 11817 -2346
rect 11753 -2407 11758 -2351
rect 11758 -2407 11814 -2351
rect 11814 -2407 11817 -2351
rect 11753 -2410 11817 -2407
rect 11833 -2351 11897 -2346
rect 11833 -2407 11838 -2351
rect 11838 -2407 11894 -2351
rect 11894 -2407 11897 -2351
rect 11833 -2410 11897 -2407
rect 12165 -2348 12229 -2343
rect 12165 -2404 12170 -2348
rect 12170 -2404 12226 -2348
rect 12226 -2404 12229 -2348
rect 12165 -2407 12229 -2404
rect 12245 -2348 12309 -2343
rect 12245 -2404 12250 -2348
rect 12250 -2404 12306 -2348
rect 12306 -2404 12309 -2348
rect 12245 -2407 12309 -2404
rect 12325 -2348 12389 -2343
rect 12325 -2404 12330 -2348
rect 12330 -2404 12386 -2348
rect 12386 -2404 12389 -2348
rect 12325 -2407 12389 -2404
rect 12405 -2348 12469 -2343
rect 12405 -2404 12410 -2348
rect 12410 -2404 12466 -2348
rect 12466 -2404 12469 -2348
rect 12405 -2407 12469 -2404
rect 12485 -2348 12549 -2343
rect 12485 -2404 12490 -2348
rect 12490 -2404 12546 -2348
rect 12546 -2404 12549 -2348
rect 12485 -2407 12549 -2404
rect 12565 -2348 12629 -2343
rect 12565 -2404 12570 -2348
rect 12570 -2404 12626 -2348
rect 12626 -2404 12629 -2348
rect 12565 -2407 12629 -2404
rect 12662 -2357 12726 -2353
rect 12662 -2413 12666 -2357
rect 12666 -2413 12722 -2357
rect 12722 -2413 12726 -2357
rect 12662 -2417 12726 -2413
<< metal4 >>
rect 106 3854 13893 3855
rect 106 3738 13943 3854
rect 106 3674 738 3738
rect 802 3732 7447 3738
rect 802 3731 6755 3732
rect 802 3728 1567 3731
rect 802 3674 835 3728
rect 106 3665 835 3674
rect 106 3133 524 3665
rect 731 3664 835 3665
rect 899 3664 915 3728
rect 979 3664 995 3728
rect 1059 3664 1075 3728
rect 1139 3664 1155 3728
rect 1219 3664 1235 3728
rect 1299 3667 1567 3728
rect 1631 3667 1647 3731
rect 1711 3667 1727 3731
rect 1791 3667 1807 3731
rect 1871 3667 1887 3731
rect 1951 3667 1967 3731
rect 2031 3667 2173 3731
rect 2237 3667 2253 3731
rect 2317 3667 2333 3731
rect 2397 3667 2413 3731
rect 2477 3667 2493 3731
rect 2557 3667 2573 3731
rect 2637 3667 2779 3731
rect 2843 3667 2859 3731
rect 2923 3667 2939 3731
rect 3003 3667 3019 3731
rect 3083 3667 3099 3731
rect 3163 3667 3179 3731
rect 3243 3667 3385 3731
rect 3449 3667 3465 3731
rect 3529 3667 3545 3731
rect 3609 3667 3625 3731
rect 3689 3667 3705 3731
rect 3769 3667 3785 3731
rect 3849 3667 3991 3731
rect 4055 3667 4071 3731
rect 4135 3667 4151 3731
rect 4215 3667 4231 3731
rect 4295 3667 4311 3731
rect 4375 3667 4391 3731
rect 4455 3667 4597 3731
rect 4661 3667 4677 3731
rect 4741 3667 4757 3731
rect 4821 3667 4837 3731
rect 4901 3667 4917 3731
rect 4981 3667 4997 3731
rect 5061 3667 5203 3731
rect 5267 3667 5283 3731
rect 5347 3667 5363 3731
rect 5427 3667 5443 3731
rect 5507 3667 5523 3731
rect 5587 3667 5603 3731
rect 5667 3667 5809 3731
rect 5873 3667 5889 3731
rect 5953 3667 5969 3731
rect 6033 3667 6049 3731
rect 6113 3667 6129 3731
rect 6193 3667 6209 3731
rect 6273 3676 6755 3731
rect 6273 3667 6547 3676
rect 1299 3665 6547 3667
rect 1299 3664 1404 3665
rect 731 3663 1404 3664
rect 731 3662 1403 3663
rect 106 3069 121 3133
rect 185 3132 396 3133
rect 185 3069 252 3132
rect 106 3068 252 3069
rect 316 3069 396 3132
rect 460 3127 524 3133
rect 731 3508 797 3598
rect 731 3444 732 3508
rect 796 3444 797 3508
rect 731 3428 797 3444
rect 731 3364 732 3428
rect 796 3364 797 3428
rect 731 3348 797 3364
rect 731 3284 732 3348
rect 796 3284 797 3348
rect 731 3268 797 3284
rect 731 3204 732 3268
rect 796 3204 797 3268
rect 731 3188 797 3204
rect 460 3069 523 3127
rect 316 3068 523 3069
rect 106 3050 523 3068
rect 731 3124 732 3188
rect 796 3124 797 3188
rect 731 3108 797 3124
rect 731 3044 732 3108
rect 796 3044 797 3108
rect 731 3028 797 3044
rect 731 2964 732 3028
rect 796 2964 797 3028
rect 731 2948 797 2964
rect 731 2884 732 2948
rect 796 2884 797 2948
rect 731 2868 797 2884
rect 731 2804 732 2868
rect 796 2804 797 2868
rect 731 2788 797 2804
rect 731 2724 732 2788
rect 796 2724 797 2788
rect 132 2587 509 2602
rect 132 2547 139 2587
rect 3 2523 139 2547
rect 203 2523 259 2587
rect 323 2523 402 2587
rect 466 2523 509 2587
rect 731 2570 797 2724
rect 857 3197 917 3662
rect 977 3197 1037 3602
rect 857 3137 1037 3197
rect 857 2632 917 3137
rect 977 2570 1037 3137
rect 1097 2632 1157 3662
rect 1217 2570 1277 3602
rect 1337 3508 1403 3598
rect 1337 3444 1338 3508
rect 1402 3444 1403 3508
rect 1337 3428 1403 3444
rect 1337 3364 1338 3428
rect 1402 3364 1403 3428
rect 1337 3348 1403 3364
rect 1337 3284 1338 3348
rect 1402 3284 1403 3348
rect 1337 3268 1403 3284
rect 1337 3204 1338 3268
rect 1402 3204 1403 3268
rect 1337 3188 1403 3204
rect 1337 3124 1338 3188
rect 1402 3124 1403 3188
rect 1337 3108 1403 3124
rect 1337 3044 1338 3108
rect 1402 3044 1403 3108
rect 1337 3028 1403 3044
rect 1337 2964 1338 3028
rect 1402 2964 1403 3028
rect 1337 2948 1403 2964
rect 1337 2884 1338 2948
rect 1402 2884 1403 2948
rect 1337 2868 1403 2884
rect 1337 2804 1338 2868
rect 1402 2804 1403 2868
rect 1337 2788 1403 2804
rect 1337 2724 1338 2788
rect 1402 2724 1403 2788
rect 1337 2570 1403 2724
rect 731 2568 1403 2570
rect 3 1707 510 2523
rect 731 2504 835 2568
rect 899 2504 915 2568
rect 979 2504 995 2568
rect 1059 2504 1075 2568
rect 1139 2504 1155 2568
rect 1219 2504 1235 2568
rect 1299 2504 1403 2568
rect 1463 3511 1529 3601
rect 1463 3447 1464 3511
rect 1528 3447 1529 3511
rect 1463 3431 1529 3447
rect 1463 3367 1464 3431
rect 1528 3367 1529 3431
rect 1463 3351 1529 3367
rect 1463 3287 1464 3351
rect 1528 3287 1529 3351
rect 1463 3271 1529 3287
rect 1463 3207 1464 3271
rect 1528 3207 1529 3271
rect 1463 3191 1529 3207
rect 1463 3127 1464 3191
rect 1528 3127 1529 3191
rect 1463 3111 1529 3127
rect 1463 3047 1464 3111
rect 1528 3047 1529 3111
rect 1463 3031 1529 3047
rect 1463 2967 1464 3031
rect 1528 2967 1529 3031
rect 1463 2951 1529 2967
rect 1463 2887 1464 2951
rect 1528 2887 1529 2951
rect 1463 2871 1529 2887
rect 1463 2807 1464 2871
rect 1528 2807 1529 2871
rect 1463 2791 1529 2807
rect 1463 2727 1464 2791
rect 1528 2727 1529 2791
rect 1463 2573 1529 2727
rect 1589 3200 1649 3665
rect 1709 3200 1769 3605
rect 1589 3140 1769 3200
rect 1589 2635 1649 3140
rect 1709 2573 1769 3140
rect 1829 2635 1889 3665
rect 1949 2573 2009 3605
rect 2069 3511 2135 3601
rect 2069 3447 2070 3511
rect 2134 3447 2135 3511
rect 2069 3431 2135 3447
rect 2069 3367 2070 3431
rect 2134 3367 2135 3431
rect 2069 3351 2135 3367
rect 2069 3287 2070 3351
rect 2134 3287 2135 3351
rect 2069 3271 2135 3287
rect 2069 3207 2070 3271
rect 2134 3207 2135 3271
rect 2069 3191 2135 3207
rect 2069 3127 2070 3191
rect 2134 3127 2135 3191
rect 2069 3111 2135 3127
rect 2069 3047 2070 3111
rect 2134 3047 2135 3111
rect 2069 3031 2135 3047
rect 2069 2967 2070 3031
rect 2134 2967 2135 3031
rect 2069 2951 2135 2967
rect 2069 2887 2070 2951
rect 2134 2887 2135 2951
rect 2069 2871 2135 2887
rect 2069 2807 2070 2871
rect 2134 2807 2135 2871
rect 2069 2791 2135 2807
rect 2069 2727 2070 2791
rect 2134 2727 2135 2791
rect 2069 2573 2135 2727
rect 2195 2573 2255 3605
rect 2315 2635 2375 3665
rect 2435 3200 2495 3605
rect 2555 3200 2615 3665
rect 2435 3140 2615 3200
rect 2435 2573 2495 3140
rect 2555 2635 2615 3140
rect 2675 3511 2741 3601
rect 2675 3447 2676 3511
rect 2740 3447 2741 3511
rect 2675 3431 2741 3447
rect 2675 3367 2676 3431
rect 2740 3367 2741 3431
rect 2675 3351 2741 3367
rect 2675 3287 2676 3351
rect 2740 3287 2741 3351
rect 2675 3271 2741 3287
rect 2675 3207 2676 3271
rect 2740 3207 2741 3271
rect 2675 3191 2741 3207
rect 2675 3127 2676 3191
rect 2740 3127 2741 3191
rect 2675 3111 2741 3127
rect 2675 3047 2676 3111
rect 2740 3047 2741 3111
rect 2675 3031 2741 3047
rect 2675 2967 2676 3031
rect 2740 2967 2741 3031
rect 2675 2951 2741 2967
rect 2675 2887 2676 2951
rect 2740 2887 2741 2951
rect 2675 2871 2741 2887
rect 2675 2807 2676 2871
rect 2740 2807 2741 2871
rect 2675 2791 2741 2807
rect 2675 2727 2676 2791
rect 2740 2727 2741 2791
rect 2675 2573 2741 2727
rect 2801 3200 2861 3665
rect 2921 3200 2981 3605
rect 2801 3140 2981 3200
rect 2801 2635 2861 3140
rect 2921 2573 2981 3140
rect 3041 2635 3101 3665
rect 3161 2573 3221 3605
rect 3281 3511 3347 3601
rect 3281 3447 3282 3511
rect 3346 3447 3347 3511
rect 3281 3431 3347 3447
rect 3281 3367 3282 3431
rect 3346 3367 3347 3431
rect 3281 3351 3347 3367
rect 3281 3287 3282 3351
rect 3346 3287 3347 3351
rect 3281 3271 3347 3287
rect 3281 3207 3282 3271
rect 3346 3207 3347 3271
rect 3281 3191 3347 3207
rect 3281 3127 3282 3191
rect 3346 3127 3347 3191
rect 3281 3111 3347 3127
rect 3281 3047 3282 3111
rect 3346 3047 3347 3111
rect 3281 3031 3347 3047
rect 3281 2967 3282 3031
rect 3346 2967 3347 3031
rect 3281 2951 3347 2967
rect 3281 2887 3282 2951
rect 3346 2887 3347 2951
rect 3281 2871 3347 2887
rect 3281 2807 3282 2871
rect 3346 2807 3347 2871
rect 3281 2791 3347 2807
rect 3281 2727 3282 2791
rect 3346 2727 3347 2791
rect 3281 2573 3347 2727
rect 3407 2573 3467 3605
rect 3527 2635 3587 3665
rect 3647 3200 3707 3605
rect 3767 3200 3827 3665
rect 3647 3140 3827 3200
rect 3647 2573 3707 3140
rect 3767 2635 3827 3140
rect 3887 3511 3953 3601
rect 3887 3447 3888 3511
rect 3952 3447 3953 3511
rect 3887 3431 3953 3447
rect 3887 3367 3888 3431
rect 3952 3367 3953 3431
rect 3887 3351 3953 3367
rect 3887 3287 3888 3351
rect 3952 3287 3953 3351
rect 3887 3271 3953 3287
rect 3887 3207 3888 3271
rect 3952 3207 3953 3271
rect 3887 3191 3953 3207
rect 3887 3127 3888 3191
rect 3952 3127 3953 3191
rect 3887 3111 3953 3127
rect 3887 3047 3888 3111
rect 3952 3047 3953 3111
rect 3887 3031 3953 3047
rect 3887 2967 3888 3031
rect 3952 2967 3953 3031
rect 3887 2951 3953 2967
rect 3887 2887 3888 2951
rect 3952 2887 3953 2951
rect 3887 2871 3953 2887
rect 3887 2807 3888 2871
rect 3952 2807 3953 2871
rect 3887 2791 3953 2807
rect 3887 2727 3888 2791
rect 3952 2727 3953 2791
rect 3887 2573 3953 2727
rect 4013 3200 4073 3665
rect 4133 3200 4193 3605
rect 4013 3140 4193 3200
rect 4013 2635 4073 3140
rect 4133 2573 4193 3140
rect 4253 2635 4313 3665
rect 4373 2573 4433 3605
rect 4493 3511 4559 3601
rect 4493 3447 4494 3511
rect 4558 3447 4559 3511
rect 4493 3431 4559 3447
rect 4493 3367 4494 3431
rect 4558 3367 4559 3431
rect 4493 3351 4559 3367
rect 4493 3287 4494 3351
rect 4558 3287 4559 3351
rect 4493 3271 4559 3287
rect 4493 3207 4494 3271
rect 4558 3207 4559 3271
rect 4493 3191 4559 3207
rect 4493 3127 4494 3191
rect 4558 3127 4559 3191
rect 4493 3111 4559 3127
rect 4493 3047 4494 3111
rect 4558 3047 4559 3111
rect 4493 3031 4559 3047
rect 4493 2967 4494 3031
rect 4558 2967 4559 3031
rect 4493 2951 4559 2967
rect 4493 2887 4494 2951
rect 4558 2887 4559 2951
rect 4493 2871 4559 2887
rect 4493 2807 4494 2871
rect 4558 2807 4559 2871
rect 4493 2791 4559 2807
rect 4493 2727 4494 2791
rect 4558 2727 4559 2791
rect 4493 2573 4559 2727
rect 4619 2573 4679 3605
rect 4739 2635 4799 3665
rect 4859 3200 4919 3605
rect 4979 3200 5039 3665
rect 4859 3140 5039 3200
rect 4859 2573 4919 3140
rect 4979 2635 5039 3140
rect 5099 3511 5165 3601
rect 5099 3447 5100 3511
rect 5164 3447 5165 3511
rect 5099 3431 5165 3447
rect 5099 3367 5100 3431
rect 5164 3367 5165 3431
rect 5099 3351 5165 3367
rect 5099 3287 5100 3351
rect 5164 3287 5165 3351
rect 5099 3271 5165 3287
rect 5099 3207 5100 3271
rect 5164 3207 5165 3271
rect 5099 3191 5165 3207
rect 5099 3127 5100 3191
rect 5164 3127 5165 3191
rect 5099 3111 5165 3127
rect 5099 3047 5100 3111
rect 5164 3047 5165 3111
rect 5099 3031 5165 3047
rect 5099 2967 5100 3031
rect 5164 2967 5165 3031
rect 5099 2951 5165 2967
rect 5099 2887 5100 2951
rect 5164 2887 5165 2951
rect 5099 2871 5165 2887
rect 5099 2807 5100 2871
rect 5164 2807 5165 2871
rect 5099 2791 5165 2807
rect 5099 2727 5100 2791
rect 5164 2727 5165 2791
rect 5099 2573 5165 2727
rect 5225 3200 5285 3665
rect 5345 3200 5405 3605
rect 5225 3140 5405 3200
rect 5225 2635 5285 3140
rect 5345 2573 5405 3140
rect 5465 2635 5525 3665
rect 5585 2573 5645 3605
rect 5705 3511 5771 3601
rect 5705 3447 5706 3511
rect 5770 3447 5771 3511
rect 5705 3431 5771 3447
rect 5705 3367 5706 3431
rect 5770 3367 5771 3431
rect 5705 3351 5771 3367
rect 5705 3287 5706 3351
rect 5770 3287 5771 3351
rect 5705 3271 5771 3287
rect 5705 3207 5706 3271
rect 5770 3207 5771 3271
rect 5705 3191 5771 3207
rect 5705 3127 5706 3191
rect 5770 3127 5771 3191
rect 5705 3111 5771 3127
rect 5705 3047 5706 3111
rect 5770 3047 5771 3111
rect 5705 3031 5771 3047
rect 5705 2967 5706 3031
rect 5770 2967 5771 3031
rect 5705 2951 5771 2967
rect 5705 2887 5706 2951
rect 5770 2887 5771 2951
rect 5705 2871 5771 2887
rect 5705 2807 5706 2871
rect 5770 2807 5771 2871
rect 5705 2791 5771 2807
rect 5705 2727 5706 2791
rect 5770 2727 5771 2791
rect 5705 2573 5771 2727
rect 5831 2573 5891 3605
rect 5951 2635 6011 3665
rect 6071 3200 6131 3605
rect 6191 3200 6251 3665
rect 6437 3612 6547 3665
rect 6611 3612 6755 3676
rect 6071 3140 6251 3200
rect 6071 2573 6131 3140
rect 6191 2635 6251 3140
rect 6311 3511 6377 3601
rect 6311 3447 6312 3511
rect 6376 3447 6377 3511
rect 6311 3431 6377 3447
rect 6311 3367 6312 3431
rect 6376 3367 6377 3431
rect 6311 3351 6377 3367
rect 6311 3287 6312 3351
rect 6376 3287 6377 3351
rect 6311 3271 6377 3287
rect 6311 3207 6312 3271
rect 6376 3207 6377 3271
rect 6311 3191 6377 3207
rect 6311 3127 6312 3191
rect 6376 3127 6377 3191
rect 6311 3111 6377 3127
rect 6311 3047 6312 3111
rect 6376 3047 6377 3111
rect 6311 3031 6377 3047
rect 6311 2967 6312 3031
rect 6376 2967 6377 3031
rect 6311 2951 6377 2967
rect 6311 2887 6312 2951
rect 6376 2887 6377 2951
rect 6311 2871 6377 2887
rect 6311 2807 6312 2871
rect 6376 2807 6377 2871
rect 6311 2791 6377 2807
rect 6311 2727 6312 2791
rect 6376 2727 6377 2791
rect 6437 3532 6755 3612
rect 6437 3468 6552 3532
rect 6616 3468 6755 3532
rect 6437 3380 6755 3468
rect 6437 3316 6553 3380
rect 6617 3316 6755 3380
rect 6437 3210 6755 3316
rect 6437 3146 6553 3210
rect 6617 3146 6755 3210
rect 6437 3053 6755 3146
rect 6437 2989 6552 3053
rect 6616 2989 6755 3053
rect 6815 3679 7447 3732
rect 6815 3615 7024 3679
rect 7088 3674 7447 3679
rect 7511 3731 13943 3738
rect 7511 3728 8276 3731
rect 7511 3674 7544 3728
rect 7088 3665 7544 3674
rect 7088 3615 7233 3665
rect 7440 3664 7544 3665
rect 7608 3664 7624 3728
rect 7688 3664 7704 3728
rect 7768 3664 7784 3728
rect 7848 3664 7864 3728
rect 7928 3664 7944 3728
rect 8008 3667 8276 3728
rect 8340 3667 8356 3731
rect 8420 3667 8436 3731
rect 8500 3667 8516 3731
rect 8580 3667 8596 3731
rect 8660 3667 8676 3731
rect 8740 3667 8882 3731
rect 8946 3667 8962 3731
rect 9026 3667 9042 3731
rect 9106 3667 9122 3731
rect 9186 3667 9202 3731
rect 9266 3667 9282 3731
rect 9346 3667 9488 3731
rect 9552 3667 9568 3731
rect 9632 3667 9648 3731
rect 9712 3667 9728 3731
rect 9792 3667 9808 3731
rect 9872 3667 9888 3731
rect 9952 3667 10094 3731
rect 10158 3667 10174 3731
rect 10238 3667 10254 3731
rect 10318 3667 10334 3731
rect 10398 3667 10414 3731
rect 10478 3667 10494 3731
rect 10558 3667 10700 3731
rect 10764 3667 10780 3731
rect 10844 3667 10860 3731
rect 10924 3667 10940 3731
rect 11004 3667 11020 3731
rect 11084 3667 11100 3731
rect 11164 3667 11306 3731
rect 11370 3667 11386 3731
rect 11450 3667 11466 3731
rect 11530 3667 11546 3731
rect 11610 3667 11626 3731
rect 11690 3667 11706 3731
rect 11770 3667 11912 3731
rect 11976 3667 11992 3731
rect 12056 3667 12072 3731
rect 12136 3667 12152 3731
rect 12216 3667 12232 3731
rect 12296 3667 12312 3731
rect 12376 3667 12518 3731
rect 12582 3667 12598 3731
rect 12662 3667 12678 3731
rect 12742 3667 12758 3731
rect 12822 3667 12838 3731
rect 12902 3667 12918 3731
rect 12982 3676 13464 3731
rect 12982 3667 13256 3676
rect 8008 3665 13256 3667
rect 8008 3664 8113 3665
rect 7440 3663 8113 3664
rect 7440 3662 8112 3663
rect 6815 3507 7233 3615
rect 6815 3443 7013 3507
rect 7077 3443 7233 3507
rect 6815 3315 7233 3443
rect 6815 3251 7013 3315
rect 7077 3251 7233 3315
rect 6815 3133 7233 3251
rect 6815 3069 6830 3133
rect 6894 3132 7105 3133
rect 6894 3069 6961 3132
rect 6815 3068 6961 3069
rect 7025 3069 7105 3132
rect 7169 3127 7233 3133
rect 7440 3508 7506 3598
rect 7440 3444 7441 3508
rect 7505 3444 7506 3508
rect 7440 3428 7506 3444
rect 7440 3364 7441 3428
rect 7505 3364 7506 3428
rect 7440 3348 7506 3364
rect 7440 3284 7441 3348
rect 7505 3284 7506 3348
rect 7440 3268 7506 3284
rect 7440 3204 7441 3268
rect 7505 3204 7506 3268
rect 7440 3188 7506 3204
rect 7169 3069 7232 3127
rect 7025 3068 7232 3069
rect 6815 3050 7232 3068
rect 7440 3124 7441 3188
rect 7505 3124 7506 3188
rect 7440 3108 7506 3124
rect 6437 2811 6755 2989
rect 6437 2747 6470 2811
rect 6534 2747 6755 2811
rect 6437 2735 6755 2747
rect 6311 2573 6377 2727
rect 1463 2571 6377 2573
rect 1463 2507 1567 2571
rect 1631 2507 1647 2571
rect 1711 2507 1727 2571
rect 1791 2507 1807 2571
rect 1871 2507 1887 2571
rect 1951 2507 1967 2571
rect 2031 2507 2173 2571
rect 2237 2507 2253 2571
rect 2317 2507 2333 2571
rect 2397 2507 2413 2571
rect 2477 2507 2493 2571
rect 2557 2507 2573 2571
rect 2637 2507 2779 2571
rect 2843 2507 2859 2571
rect 2923 2507 2939 2571
rect 3003 2507 3019 2571
rect 3083 2507 3099 2571
rect 3163 2507 3179 2571
rect 3243 2507 3385 2571
rect 3449 2507 3465 2571
rect 3529 2507 3545 2571
rect 3609 2507 3625 2571
rect 3689 2507 3705 2571
rect 3769 2507 3785 2571
rect 3849 2507 3991 2571
rect 4055 2507 4071 2571
rect 4135 2507 4151 2571
rect 4215 2507 4231 2571
rect 4295 2507 4311 2571
rect 4375 2507 4391 2571
rect 4455 2507 4597 2571
rect 4661 2507 4677 2571
rect 4741 2507 4757 2571
rect 4821 2507 4837 2571
rect 4901 2507 4917 2571
rect 4981 2507 4997 2571
rect 5061 2507 5203 2571
rect 5267 2507 5283 2571
rect 5347 2507 5363 2571
rect 5427 2507 5443 2571
rect 5507 2507 5523 2571
rect 5587 2507 5603 2571
rect 5667 2507 5809 2571
rect 5873 2507 5889 2571
rect 5953 2507 5969 2571
rect 6033 2507 6049 2571
rect 6113 2507 6129 2571
rect 6193 2507 6209 2571
rect 6273 2507 6377 2571
rect 1463 2505 6377 2507
rect 6437 2550 6635 2560
rect 731 2502 1403 2504
rect 6437 2486 6558 2550
rect 6622 2486 6635 2550
rect 6437 2476 6635 2486
rect 3 1643 106 1707
rect 171 1643 510 1707
rect 3 1164 510 1643
rect 1082 2323 1754 2325
rect 1082 2259 1186 2323
rect 1250 2259 1266 2323
rect 1330 2259 1346 2323
rect 1410 2259 1426 2323
rect 1490 2259 1506 2323
rect 1570 2259 1586 2323
rect 1650 2259 1754 2323
rect 1082 2257 1754 2259
rect 1082 2103 1148 2257
rect 1082 2039 1083 2103
rect 1147 2039 1148 2103
rect 1082 2023 1148 2039
rect 1082 1959 1083 2023
rect 1147 1959 1148 2023
rect 1082 1943 1148 1959
rect 1082 1879 1083 1943
rect 1147 1879 1148 1943
rect 1082 1863 1148 1879
rect 1082 1799 1083 1863
rect 1147 1799 1148 1863
rect 1082 1783 1148 1799
rect 1082 1719 1083 1783
rect 1147 1719 1148 1783
rect 1082 1703 1148 1719
rect 1082 1639 1083 1703
rect 1147 1639 1148 1703
rect 1082 1623 1148 1639
rect 1082 1559 1083 1623
rect 1147 1559 1148 1623
rect 1082 1543 1148 1559
rect 1082 1479 1083 1543
rect 1147 1479 1148 1543
rect 1082 1463 1148 1479
rect 1082 1399 1083 1463
rect 1147 1399 1148 1463
rect 1082 1383 1148 1399
rect 1082 1319 1083 1383
rect 1147 1319 1148 1383
rect 1082 1229 1148 1319
rect 1208 1563 1268 2195
rect 1328 1563 1388 2257
rect 1208 1487 1388 1563
rect 694 1164 819 1170
rect 1208 1165 1268 1487
rect 1328 1225 1388 1487
rect 1448 1165 1508 2195
rect 1568 1225 1628 2257
rect 1688 2103 1754 2257
rect 1688 2039 1689 2103
rect 1753 2039 1754 2103
rect 1688 2023 1754 2039
rect 1688 1959 1689 2023
rect 1753 1959 1754 2023
rect 1688 1943 1754 1959
rect 1688 1879 1689 1943
rect 1753 1879 1754 1943
rect 1688 1863 1754 1879
rect 1688 1799 1689 1863
rect 1753 1799 1754 1863
rect 1688 1783 1754 1799
rect 1688 1719 1689 1783
rect 1753 1719 1754 1783
rect 1688 1703 1754 1719
rect 1688 1639 1689 1703
rect 1753 1639 1754 1703
rect 1688 1623 1754 1639
rect 1688 1559 1689 1623
rect 1753 1559 1754 1623
rect 1688 1543 1754 1559
rect 1688 1479 1689 1543
rect 1753 1479 1754 1543
rect 1688 1463 1754 1479
rect 1688 1399 1689 1463
rect 1753 1399 1754 1463
rect 1688 1383 1754 1399
rect 1688 1319 1689 1383
rect 1753 1319 1754 1383
rect 1688 1229 1754 1319
rect 1814 2323 4304 2325
rect 1814 2259 1918 2323
rect 1982 2259 1998 2323
rect 2062 2259 2078 2323
rect 2142 2259 2158 2323
rect 2222 2259 2238 2323
rect 2302 2259 2318 2323
rect 2382 2259 2524 2323
rect 2588 2259 2604 2323
rect 2668 2259 2684 2323
rect 2748 2259 2764 2323
rect 2828 2259 2844 2323
rect 2908 2259 2924 2323
rect 2988 2259 3130 2323
rect 3194 2259 3210 2323
rect 3274 2259 3290 2323
rect 3354 2259 3370 2323
rect 3434 2259 3450 2323
rect 3514 2259 3530 2323
rect 3594 2259 3736 2323
rect 3800 2259 3816 2323
rect 3880 2259 3896 2323
rect 3960 2259 3976 2323
rect 4040 2259 4056 2323
rect 4120 2259 4136 2323
rect 4200 2259 4304 2323
rect 1814 2257 4304 2259
rect 1814 2103 1880 2257
rect 1814 2039 1815 2103
rect 1879 2039 1880 2103
rect 1814 2023 1880 2039
rect 1814 1959 1815 2023
rect 1879 1959 1880 2023
rect 1814 1943 1880 1959
rect 1814 1879 1815 1943
rect 1879 1879 1880 1943
rect 1814 1863 1880 1879
rect 1814 1799 1815 1863
rect 1879 1799 1880 1863
rect 1814 1783 1880 1799
rect 1814 1719 1815 1783
rect 1879 1719 1880 1783
rect 1814 1703 1880 1719
rect 1814 1639 1815 1703
rect 1879 1639 1880 1703
rect 1814 1623 1880 1639
rect 1814 1559 1815 1623
rect 1879 1559 1880 1623
rect 1814 1543 1880 1559
rect 1814 1479 1815 1543
rect 1879 1479 1880 1543
rect 1814 1463 1880 1479
rect 1814 1399 1815 1463
rect 1879 1399 1880 1463
rect 1814 1383 1880 1399
rect 1814 1319 1815 1383
rect 1879 1319 1880 1383
rect 1814 1229 1880 1319
rect 1940 1563 2000 2195
rect 2060 1563 2120 2257
rect 1940 1487 2120 1563
rect 1940 1165 2000 1487
rect 2060 1225 2120 1487
rect 2180 1165 2240 2195
rect 2300 1225 2360 2257
rect 2420 2103 2486 2257
rect 2420 2039 2421 2103
rect 2485 2039 2486 2103
rect 2420 2023 2486 2039
rect 2420 1959 2421 2023
rect 2485 1959 2486 2023
rect 2420 1943 2486 1959
rect 2420 1879 2421 1943
rect 2485 1879 2486 1943
rect 2420 1863 2486 1879
rect 2420 1799 2421 1863
rect 2485 1799 2486 1863
rect 2420 1783 2486 1799
rect 2420 1719 2421 1783
rect 2485 1719 2486 1783
rect 2420 1703 2486 1719
rect 2420 1639 2421 1703
rect 2485 1639 2486 1703
rect 2420 1623 2486 1639
rect 2420 1559 2421 1623
rect 2485 1559 2486 1623
rect 2420 1543 2486 1559
rect 2420 1479 2421 1543
rect 2485 1479 2486 1543
rect 2420 1463 2486 1479
rect 2420 1399 2421 1463
rect 2485 1399 2486 1463
rect 2420 1383 2486 1399
rect 2420 1319 2421 1383
rect 2485 1319 2486 1383
rect 2420 1229 2486 1319
rect 2546 1225 2606 2257
rect 2666 1165 2726 2195
rect 2786 1563 2846 2257
rect 2906 1563 2966 2195
rect 2786 1487 2966 1563
rect 2786 1225 2846 1487
rect 2906 1165 2966 1487
rect 3026 2103 3092 2257
rect 3026 2039 3027 2103
rect 3091 2039 3092 2103
rect 3026 2023 3092 2039
rect 3026 1959 3027 2023
rect 3091 1959 3092 2023
rect 3026 1943 3092 1959
rect 3026 1879 3027 1943
rect 3091 1879 3092 1943
rect 3026 1863 3092 1879
rect 3026 1799 3027 1863
rect 3091 1799 3092 1863
rect 3026 1783 3092 1799
rect 3026 1719 3027 1783
rect 3091 1719 3092 1783
rect 3026 1703 3092 1719
rect 3026 1639 3027 1703
rect 3091 1639 3092 1703
rect 3026 1623 3092 1639
rect 3026 1559 3027 1623
rect 3091 1559 3092 1623
rect 3026 1543 3092 1559
rect 3026 1479 3027 1543
rect 3091 1479 3092 1543
rect 3026 1463 3092 1479
rect 3026 1399 3027 1463
rect 3091 1399 3092 1463
rect 3026 1383 3092 1399
rect 3026 1319 3027 1383
rect 3091 1319 3092 1383
rect 3026 1229 3092 1319
rect 3152 1563 3212 2195
rect 3272 1563 3332 2257
rect 3152 1487 3332 1563
rect 3152 1165 3212 1487
rect 3272 1225 3332 1487
rect 3392 1165 3452 2195
rect 3512 1225 3572 2257
rect 3632 2103 3698 2257
rect 3632 2039 3633 2103
rect 3697 2039 3698 2103
rect 3632 2023 3698 2039
rect 3632 1959 3633 2023
rect 3697 1959 3698 2023
rect 3632 1943 3698 1959
rect 3632 1879 3633 1943
rect 3697 1879 3698 1943
rect 3632 1863 3698 1879
rect 3632 1799 3633 1863
rect 3697 1799 3698 1863
rect 3632 1783 3698 1799
rect 3632 1719 3633 1783
rect 3697 1719 3698 1783
rect 3632 1703 3698 1719
rect 3632 1639 3633 1703
rect 3697 1639 3698 1703
rect 3632 1623 3698 1639
rect 3632 1559 3633 1623
rect 3697 1559 3698 1623
rect 3632 1543 3698 1559
rect 3632 1479 3633 1543
rect 3697 1479 3698 1543
rect 3632 1463 3698 1479
rect 3632 1399 3633 1463
rect 3697 1399 3698 1463
rect 3632 1383 3698 1399
rect 3632 1319 3633 1383
rect 3697 1319 3698 1383
rect 3632 1229 3698 1319
rect 3758 1225 3818 2257
rect 3878 1165 3938 2195
rect 3998 1563 4058 2257
rect 4118 1563 4178 2195
rect 3998 1487 4178 1563
rect 3998 1225 4058 1487
rect 4118 1165 4178 1487
rect 4238 2103 4304 2257
rect 4238 2039 4239 2103
rect 4303 2039 4304 2103
rect 4238 2023 4304 2039
rect 4238 1959 4239 2023
rect 4303 1959 4304 2023
rect 4238 1943 4304 1959
rect 4238 1879 4239 1943
rect 4303 1879 4304 1943
rect 4238 1863 4304 1879
rect 4238 1799 4239 1863
rect 4303 1799 4304 1863
rect 4238 1783 4304 1799
rect 4238 1719 4239 1783
rect 4303 1719 4304 1783
rect 4238 1703 4304 1719
rect 4238 1639 4239 1703
rect 4303 1639 4304 1703
rect 4238 1623 4304 1639
rect 4238 1559 4239 1623
rect 4303 1559 4304 1623
rect 4238 1543 4304 1559
rect 4238 1479 4239 1543
rect 4303 1479 4304 1543
rect 4238 1463 4304 1479
rect 4238 1399 4239 1463
rect 4303 1399 4304 1463
rect 4238 1383 4304 1399
rect 4238 1319 4239 1383
rect 4303 1319 4304 1383
rect 4238 1229 4304 1319
rect 4364 2323 5642 2325
rect 4364 2259 4468 2323
rect 4532 2259 4548 2323
rect 4612 2259 4628 2323
rect 4692 2259 4708 2323
rect 4772 2259 4788 2323
rect 4852 2259 4868 2323
rect 4932 2259 5074 2323
rect 5138 2259 5154 2323
rect 5218 2259 5234 2323
rect 5298 2259 5314 2323
rect 5378 2259 5394 2323
rect 5458 2259 5474 2323
rect 5538 2259 5642 2323
rect 4364 2257 5642 2259
rect 4364 2103 4430 2257
rect 4364 2039 4365 2103
rect 4429 2039 4430 2103
rect 4364 2023 4430 2039
rect 4364 1959 4365 2023
rect 4429 1959 4430 2023
rect 4364 1943 4430 1959
rect 4364 1879 4365 1943
rect 4429 1879 4430 1943
rect 4364 1863 4430 1879
rect 4364 1799 4365 1863
rect 4429 1799 4430 1863
rect 4364 1783 4430 1799
rect 4364 1719 4365 1783
rect 4429 1719 4430 1783
rect 4364 1703 4430 1719
rect 4364 1639 4365 1703
rect 4429 1639 4430 1703
rect 4364 1623 4430 1639
rect 4364 1559 4365 1623
rect 4429 1559 4430 1623
rect 4364 1543 4430 1559
rect 4364 1479 4365 1543
rect 4429 1479 4430 1543
rect 4364 1463 4430 1479
rect 4364 1399 4365 1463
rect 4429 1399 4430 1463
rect 4364 1383 4430 1399
rect 4364 1319 4365 1383
rect 4429 1319 4430 1383
rect 4364 1229 4430 1319
rect 4490 1563 4550 2195
rect 4610 1563 4670 2257
rect 4490 1487 4670 1563
rect 4490 1165 4550 1487
rect 4610 1225 4670 1487
rect 4730 1165 4790 2195
rect 4850 1225 4910 2257
rect 4970 2103 5036 2257
rect 4970 2039 4971 2103
rect 5035 2039 5036 2103
rect 4970 2023 5036 2039
rect 4970 1959 4971 2023
rect 5035 1959 5036 2023
rect 4970 1943 5036 1959
rect 4970 1879 4971 1943
rect 5035 1879 5036 1943
rect 4970 1863 5036 1879
rect 4970 1799 4971 1863
rect 5035 1799 5036 1863
rect 4970 1783 5036 1799
rect 4970 1719 4971 1783
rect 5035 1719 5036 1783
rect 4970 1703 5036 1719
rect 4970 1639 4971 1703
rect 5035 1639 5036 1703
rect 4970 1623 5036 1639
rect 4970 1559 4971 1623
rect 5035 1559 5036 1623
rect 4970 1543 5036 1559
rect 4970 1479 4971 1543
rect 5035 1479 5036 1543
rect 4970 1463 5036 1479
rect 4970 1399 4971 1463
rect 5035 1399 5036 1463
rect 4970 1383 5036 1399
rect 4970 1319 4971 1383
rect 5035 1319 5036 1383
rect 4970 1229 5036 1319
rect 5096 1225 5156 2257
rect 5216 1165 5276 2195
rect 5336 1563 5396 2257
rect 5456 1563 5516 2195
rect 5336 1487 5516 1563
rect 5336 1225 5396 1487
rect 5456 1165 5516 1487
rect 5576 2103 5642 2257
rect 5576 2039 5577 2103
rect 5641 2039 5642 2103
rect 5576 2023 5642 2039
rect 5576 1959 5577 2023
rect 5641 1959 5642 2023
rect 5576 1943 5642 1959
rect 5576 1879 5577 1943
rect 5641 1879 5642 1943
rect 5576 1863 5642 1879
rect 5576 1799 5577 1863
rect 5641 1799 5642 1863
rect 5576 1783 5642 1799
rect 5576 1719 5577 1783
rect 5641 1719 5642 1783
rect 5576 1703 5642 1719
rect 5576 1639 5577 1703
rect 5641 1639 5642 1703
rect 5576 1623 5642 1639
rect 5576 1559 5577 1623
rect 5641 1559 5642 1623
rect 5576 1543 5642 1559
rect 5576 1479 5577 1543
rect 5641 1479 5642 1543
rect 5576 1463 5642 1479
rect 5576 1399 5577 1463
rect 5641 1399 5642 1463
rect 5576 1383 5642 1399
rect 5576 1319 5577 1383
rect 5641 1319 5642 1383
rect 5576 1229 5642 1319
rect 5704 2323 6376 2325
rect 5704 2259 5808 2323
rect 5872 2259 5888 2323
rect 5952 2259 5968 2323
rect 6032 2259 6048 2323
rect 6112 2259 6128 2323
rect 6192 2259 6208 2323
rect 6272 2259 6376 2323
rect 5704 2257 6376 2259
rect 5704 2103 5770 2257
rect 5704 2039 5705 2103
rect 5769 2039 5770 2103
rect 5704 2023 5770 2039
rect 5704 1959 5705 2023
rect 5769 1959 5770 2023
rect 5704 1943 5770 1959
rect 5704 1879 5705 1943
rect 5769 1879 5770 1943
rect 5704 1863 5770 1879
rect 5704 1799 5705 1863
rect 5769 1799 5770 1863
rect 5704 1783 5770 1799
rect 5704 1719 5705 1783
rect 5769 1719 5770 1783
rect 5704 1703 5770 1719
rect 5704 1639 5705 1703
rect 5769 1639 5770 1703
rect 5704 1623 5770 1639
rect 5704 1559 5705 1623
rect 5769 1559 5770 1623
rect 5704 1543 5770 1559
rect 5704 1479 5705 1543
rect 5769 1479 5770 1543
rect 5704 1463 5770 1479
rect 5704 1399 5705 1463
rect 5769 1399 5770 1463
rect 5704 1383 5770 1399
rect 5704 1319 5705 1383
rect 5769 1319 5770 1383
rect 5704 1229 5770 1319
rect 5830 1225 5890 2257
rect 5950 1165 6010 2195
rect 6070 1563 6130 2257
rect 6190 1563 6250 2195
rect 6070 1487 6250 1563
rect 6070 1225 6130 1487
rect 6190 1165 6250 1487
rect 6310 2103 6376 2257
rect 6310 2039 6311 2103
rect 6375 2039 6376 2103
rect 6310 2023 6376 2039
rect 6310 1959 6311 2023
rect 6375 1959 6376 2023
rect 6310 1943 6376 1959
rect 6310 1879 6311 1943
rect 6375 1879 6376 1943
rect 6310 1863 6376 1879
rect 6310 1799 6311 1863
rect 6375 1799 6376 1863
rect 6310 1783 6376 1799
rect 6310 1719 6311 1783
rect 6375 1719 6376 1783
rect 6310 1703 6376 1719
rect 6310 1639 6311 1703
rect 6375 1639 6376 1703
rect 6310 1623 6376 1639
rect 6310 1559 6311 1623
rect 6375 1559 6376 1623
rect 6310 1543 6376 1559
rect 6310 1479 6311 1543
rect 6375 1479 6376 1543
rect 6310 1463 6376 1479
rect 6310 1399 6311 1463
rect 6375 1399 6376 1463
rect 6310 1383 6376 1399
rect 6310 1319 6311 1383
rect 6375 1319 6376 1383
rect 6310 1229 6376 1319
rect 6437 2095 6497 2476
rect 6695 2357 6755 2735
rect 7440 3044 7441 3108
rect 7505 3044 7506 3108
rect 7440 3028 7506 3044
rect 7440 2964 7441 3028
rect 7505 2964 7506 3028
rect 7440 2948 7506 2964
rect 7440 2884 7441 2948
rect 7505 2884 7506 2948
rect 7440 2868 7506 2884
rect 7440 2804 7441 2868
rect 7505 2804 7506 2868
rect 7440 2788 7506 2804
rect 7440 2724 7441 2788
rect 7505 2724 7506 2788
rect 6841 2587 7218 2602
rect 6841 2523 6848 2587
rect 6912 2523 6968 2587
rect 7032 2523 7111 2587
rect 7175 2523 7218 2587
rect 7440 2570 7506 2724
rect 7566 3197 7626 3662
rect 7686 3197 7746 3602
rect 7566 3137 7746 3197
rect 7566 2632 7626 3137
rect 7686 2570 7746 3137
rect 7806 2632 7866 3662
rect 7926 2570 7986 3602
rect 8046 3508 8112 3598
rect 8046 3444 8047 3508
rect 8111 3444 8112 3508
rect 8046 3428 8112 3444
rect 8046 3364 8047 3428
rect 8111 3364 8112 3428
rect 8046 3348 8112 3364
rect 8046 3284 8047 3348
rect 8111 3284 8112 3348
rect 8046 3268 8112 3284
rect 8046 3204 8047 3268
rect 8111 3204 8112 3268
rect 8046 3188 8112 3204
rect 8046 3124 8047 3188
rect 8111 3124 8112 3188
rect 8046 3108 8112 3124
rect 8046 3044 8047 3108
rect 8111 3044 8112 3108
rect 8046 3028 8112 3044
rect 8046 2964 8047 3028
rect 8111 2964 8112 3028
rect 8046 2948 8112 2964
rect 8046 2884 8047 2948
rect 8111 2884 8112 2948
rect 8046 2868 8112 2884
rect 8046 2804 8047 2868
rect 8111 2804 8112 2868
rect 8046 2788 8112 2804
rect 8046 2724 8047 2788
rect 8111 2724 8112 2788
rect 8046 2570 8112 2724
rect 7440 2568 8112 2570
rect 6557 2347 6755 2357
rect 6557 2283 6558 2347
rect 6622 2283 6755 2347
rect 6557 2273 6755 2283
rect 6437 2085 6755 2095
rect 6437 2021 6467 2085
rect 6531 2021 6755 2085
rect 1082 1164 1754 1165
rect 1814 1164 4304 1165
rect 4364 1164 5642 1165
rect 5704 1164 6376 1165
rect 6437 1164 6755 2021
rect 3 1163 6755 1164
rect 3 1160 1266 1163
rect 3 1096 724 1160
rect 788 1099 1266 1160
rect 1330 1099 1346 1163
rect 1410 1099 1426 1163
rect 1490 1099 1506 1163
rect 1570 1099 1998 1163
rect 2062 1099 2078 1163
rect 2142 1099 2158 1163
rect 2222 1099 2238 1163
rect 2302 1099 2604 1163
rect 2668 1099 2684 1163
rect 2748 1099 2764 1163
rect 2828 1099 2844 1163
rect 2908 1099 3210 1163
rect 3274 1099 3290 1163
rect 3354 1099 3370 1163
rect 3434 1099 3450 1163
rect 3514 1099 3816 1163
rect 3880 1099 3896 1163
rect 3960 1099 3976 1163
rect 4040 1099 4056 1163
rect 4120 1099 4548 1163
rect 4612 1099 4628 1163
rect 4692 1099 4708 1163
rect 4772 1099 4788 1163
rect 4852 1099 5154 1163
rect 5218 1099 5234 1163
rect 5298 1099 5314 1163
rect 5378 1099 5394 1163
rect 5458 1099 5888 1163
rect 5952 1099 5968 1163
rect 6032 1099 6048 1163
rect 6112 1099 6128 1163
rect 6192 1150 6755 1163
rect 6843 1164 7219 2523
rect 7440 2504 7544 2568
rect 7608 2504 7624 2568
rect 7688 2504 7704 2568
rect 7768 2504 7784 2568
rect 7848 2504 7864 2568
rect 7928 2504 7944 2568
rect 8008 2504 8112 2568
rect 8172 3511 8238 3601
rect 8172 3447 8173 3511
rect 8237 3447 8238 3511
rect 8172 3431 8238 3447
rect 8172 3367 8173 3431
rect 8237 3367 8238 3431
rect 8172 3351 8238 3367
rect 8172 3287 8173 3351
rect 8237 3287 8238 3351
rect 8172 3271 8238 3287
rect 8172 3207 8173 3271
rect 8237 3207 8238 3271
rect 8172 3191 8238 3207
rect 8172 3127 8173 3191
rect 8237 3127 8238 3191
rect 8172 3111 8238 3127
rect 8172 3047 8173 3111
rect 8237 3047 8238 3111
rect 8172 3031 8238 3047
rect 8172 2967 8173 3031
rect 8237 2967 8238 3031
rect 8172 2951 8238 2967
rect 8172 2887 8173 2951
rect 8237 2887 8238 2951
rect 8172 2871 8238 2887
rect 8172 2807 8173 2871
rect 8237 2807 8238 2871
rect 8172 2791 8238 2807
rect 8172 2727 8173 2791
rect 8237 2727 8238 2791
rect 8172 2573 8238 2727
rect 8298 3200 8358 3665
rect 8418 3200 8478 3605
rect 8298 3140 8478 3200
rect 8298 2635 8358 3140
rect 8418 2573 8478 3140
rect 8538 2635 8598 3665
rect 8658 2573 8718 3605
rect 8778 3511 8844 3601
rect 8778 3447 8779 3511
rect 8843 3447 8844 3511
rect 8778 3431 8844 3447
rect 8778 3367 8779 3431
rect 8843 3367 8844 3431
rect 8778 3351 8844 3367
rect 8778 3287 8779 3351
rect 8843 3287 8844 3351
rect 8778 3271 8844 3287
rect 8778 3207 8779 3271
rect 8843 3207 8844 3271
rect 8778 3191 8844 3207
rect 8778 3127 8779 3191
rect 8843 3127 8844 3191
rect 8778 3111 8844 3127
rect 8778 3047 8779 3111
rect 8843 3047 8844 3111
rect 8778 3031 8844 3047
rect 8778 2967 8779 3031
rect 8843 2967 8844 3031
rect 8778 2951 8844 2967
rect 8778 2887 8779 2951
rect 8843 2887 8844 2951
rect 8778 2871 8844 2887
rect 8778 2807 8779 2871
rect 8843 2807 8844 2871
rect 8778 2791 8844 2807
rect 8778 2727 8779 2791
rect 8843 2727 8844 2791
rect 8778 2573 8844 2727
rect 8904 2573 8964 3605
rect 9024 2635 9084 3665
rect 9144 3200 9204 3605
rect 9264 3200 9324 3665
rect 9144 3140 9324 3200
rect 9144 2573 9204 3140
rect 9264 2635 9324 3140
rect 9384 3511 9450 3601
rect 9384 3447 9385 3511
rect 9449 3447 9450 3511
rect 9384 3431 9450 3447
rect 9384 3367 9385 3431
rect 9449 3367 9450 3431
rect 9384 3351 9450 3367
rect 9384 3287 9385 3351
rect 9449 3287 9450 3351
rect 9384 3271 9450 3287
rect 9384 3207 9385 3271
rect 9449 3207 9450 3271
rect 9384 3191 9450 3207
rect 9384 3127 9385 3191
rect 9449 3127 9450 3191
rect 9384 3111 9450 3127
rect 9384 3047 9385 3111
rect 9449 3047 9450 3111
rect 9384 3031 9450 3047
rect 9384 2967 9385 3031
rect 9449 2967 9450 3031
rect 9384 2951 9450 2967
rect 9384 2887 9385 2951
rect 9449 2887 9450 2951
rect 9384 2871 9450 2887
rect 9384 2807 9385 2871
rect 9449 2807 9450 2871
rect 9384 2791 9450 2807
rect 9384 2727 9385 2791
rect 9449 2727 9450 2791
rect 9384 2573 9450 2727
rect 9510 3200 9570 3665
rect 9630 3200 9690 3605
rect 9510 3140 9690 3200
rect 9510 2635 9570 3140
rect 9630 2573 9690 3140
rect 9750 2635 9810 3665
rect 9870 2573 9930 3605
rect 9990 3511 10056 3601
rect 9990 3447 9991 3511
rect 10055 3447 10056 3511
rect 9990 3431 10056 3447
rect 9990 3367 9991 3431
rect 10055 3367 10056 3431
rect 9990 3351 10056 3367
rect 9990 3287 9991 3351
rect 10055 3287 10056 3351
rect 9990 3271 10056 3287
rect 9990 3207 9991 3271
rect 10055 3207 10056 3271
rect 9990 3191 10056 3207
rect 9990 3127 9991 3191
rect 10055 3127 10056 3191
rect 9990 3111 10056 3127
rect 9990 3047 9991 3111
rect 10055 3047 10056 3111
rect 9990 3031 10056 3047
rect 9990 2967 9991 3031
rect 10055 2967 10056 3031
rect 9990 2951 10056 2967
rect 9990 2887 9991 2951
rect 10055 2887 10056 2951
rect 9990 2871 10056 2887
rect 9990 2807 9991 2871
rect 10055 2807 10056 2871
rect 9990 2791 10056 2807
rect 9990 2727 9991 2791
rect 10055 2727 10056 2791
rect 9990 2573 10056 2727
rect 10116 2573 10176 3605
rect 10236 2635 10296 3665
rect 10356 3200 10416 3605
rect 10476 3200 10536 3665
rect 10356 3140 10536 3200
rect 10356 2573 10416 3140
rect 10476 2635 10536 3140
rect 10596 3511 10662 3601
rect 10596 3447 10597 3511
rect 10661 3447 10662 3511
rect 10596 3431 10662 3447
rect 10596 3367 10597 3431
rect 10661 3367 10662 3431
rect 10596 3351 10662 3367
rect 10596 3287 10597 3351
rect 10661 3287 10662 3351
rect 10596 3271 10662 3287
rect 10596 3207 10597 3271
rect 10661 3207 10662 3271
rect 10596 3191 10662 3207
rect 10596 3127 10597 3191
rect 10661 3127 10662 3191
rect 10596 3111 10662 3127
rect 10596 3047 10597 3111
rect 10661 3047 10662 3111
rect 10596 3031 10662 3047
rect 10596 2967 10597 3031
rect 10661 2967 10662 3031
rect 10596 2951 10662 2967
rect 10596 2887 10597 2951
rect 10661 2887 10662 2951
rect 10596 2871 10662 2887
rect 10596 2807 10597 2871
rect 10661 2807 10662 2871
rect 10596 2791 10662 2807
rect 10596 2727 10597 2791
rect 10661 2727 10662 2791
rect 10596 2573 10662 2727
rect 10722 3200 10782 3665
rect 10842 3200 10902 3605
rect 10722 3140 10902 3200
rect 10722 2635 10782 3140
rect 10842 2573 10902 3140
rect 10962 2635 11022 3665
rect 11082 2573 11142 3605
rect 11202 3511 11268 3601
rect 11202 3447 11203 3511
rect 11267 3447 11268 3511
rect 11202 3431 11268 3447
rect 11202 3367 11203 3431
rect 11267 3367 11268 3431
rect 11202 3351 11268 3367
rect 11202 3287 11203 3351
rect 11267 3287 11268 3351
rect 11202 3271 11268 3287
rect 11202 3207 11203 3271
rect 11267 3207 11268 3271
rect 11202 3191 11268 3207
rect 11202 3127 11203 3191
rect 11267 3127 11268 3191
rect 11202 3111 11268 3127
rect 11202 3047 11203 3111
rect 11267 3047 11268 3111
rect 11202 3031 11268 3047
rect 11202 2967 11203 3031
rect 11267 2967 11268 3031
rect 11202 2951 11268 2967
rect 11202 2887 11203 2951
rect 11267 2887 11268 2951
rect 11202 2871 11268 2887
rect 11202 2807 11203 2871
rect 11267 2807 11268 2871
rect 11202 2791 11268 2807
rect 11202 2727 11203 2791
rect 11267 2727 11268 2791
rect 11202 2573 11268 2727
rect 11328 2573 11388 3605
rect 11448 2635 11508 3665
rect 11568 3200 11628 3605
rect 11688 3200 11748 3665
rect 11568 3140 11748 3200
rect 11568 2573 11628 3140
rect 11688 2635 11748 3140
rect 11808 3511 11874 3601
rect 11808 3447 11809 3511
rect 11873 3447 11874 3511
rect 11808 3431 11874 3447
rect 11808 3367 11809 3431
rect 11873 3367 11874 3431
rect 11808 3351 11874 3367
rect 11808 3287 11809 3351
rect 11873 3287 11874 3351
rect 11808 3271 11874 3287
rect 11808 3207 11809 3271
rect 11873 3207 11874 3271
rect 11808 3191 11874 3207
rect 11808 3127 11809 3191
rect 11873 3127 11874 3191
rect 11808 3111 11874 3127
rect 11808 3047 11809 3111
rect 11873 3047 11874 3111
rect 11808 3031 11874 3047
rect 11808 2967 11809 3031
rect 11873 2967 11874 3031
rect 11808 2951 11874 2967
rect 11808 2887 11809 2951
rect 11873 2887 11874 2951
rect 11808 2871 11874 2887
rect 11808 2807 11809 2871
rect 11873 2807 11874 2871
rect 11808 2791 11874 2807
rect 11808 2727 11809 2791
rect 11873 2727 11874 2791
rect 11808 2573 11874 2727
rect 11934 3200 11994 3665
rect 12054 3200 12114 3605
rect 11934 3140 12114 3200
rect 11934 2635 11994 3140
rect 12054 2573 12114 3140
rect 12174 2635 12234 3665
rect 12294 2573 12354 3605
rect 12414 3511 12480 3601
rect 12414 3447 12415 3511
rect 12479 3447 12480 3511
rect 12414 3431 12480 3447
rect 12414 3367 12415 3431
rect 12479 3367 12480 3431
rect 12414 3351 12480 3367
rect 12414 3287 12415 3351
rect 12479 3287 12480 3351
rect 12414 3271 12480 3287
rect 12414 3207 12415 3271
rect 12479 3207 12480 3271
rect 12414 3191 12480 3207
rect 12414 3127 12415 3191
rect 12479 3127 12480 3191
rect 12414 3111 12480 3127
rect 12414 3047 12415 3111
rect 12479 3047 12480 3111
rect 12414 3031 12480 3047
rect 12414 2967 12415 3031
rect 12479 2967 12480 3031
rect 12414 2951 12480 2967
rect 12414 2887 12415 2951
rect 12479 2887 12480 2951
rect 12414 2871 12480 2887
rect 12414 2807 12415 2871
rect 12479 2807 12480 2871
rect 12414 2791 12480 2807
rect 12414 2727 12415 2791
rect 12479 2727 12480 2791
rect 12414 2573 12480 2727
rect 12540 2573 12600 3605
rect 12660 2635 12720 3665
rect 12780 3200 12840 3605
rect 12900 3200 12960 3665
rect 13146 3612 13256 3665
rect 13320 3612 13464 3676
rect 12780 3140 12960 3200
rect 12780 2573 12840 3140
rect 12900 2635 12960 3140
rect 13020 3511 13086 3601
rect 13020 3447 13021 3511
rect 13085 3447 13086 3511
rect 13020 3431 13086 3447
rect 13020 3367 13021 3431
rect 13085 3367 13086 3431
rect 13020 3351 13086 3367
rect 13020 3287 13021 3351
rect 13085 3287 13086 3351
rect 13020 3271 13086 3287
rect 13020 3207 13021 3271
rect 13085 3207 13086 3271
rect 13020 3191 13086 3207
rect 13020 3127 13021 3191
rect 13085 3127 13086 3191
rect 13020 3111 13086 3127
rect 13020 3047 13021 3111
rect 13085 3047 13086 3111
rect 13020 3031 13086 3047
rect 13020 2967 13021 3031
rect 13085 2967 13086 3031
rect 13020 2951 13086 2967
rect 13020 2887 13021 2951
rect 13085 2887 13086 2951
rect 13020 2871 13086 2887
rect 13020 2807 13021 2871
rect 13085 2807 13086 2871
rect 13020 2791 13086 2807
rect 13020 2727 13021 2791
rect 13085 2727 13086 2791
rect 13146 3532 13464 3612
rect 13146 3468 13261 3532
rect 13325 3468 13464 3532
rect 13146 3380 13464 3468
rect 13146 3316 13262 3380
rect 13326 3316 13464 3380
rect 13146 3210 13464 3316
rect 13146 3146 13262 3210
rect 13326 3146 13464 3210
rect 13146 3053 13464 3146
rect 13146 2989 13261 3053
rect 13325 2989 13464 3053
rect 13146 2811 13464 2989
rect 13146 2747 13179 2811
rect 13243 2747 13464 2811
rect 13146 2735 13464 2747
rect 13020 2573 13086 2727
rect 8172 2571 13086 2573
rect 8172 2507 8276 2571
rect 8340 2507 8356 2571
rect 8420 2507 8436 2571
rect 8500 2507 8516 2571
rect 8580 2507 8596 2571
rect 8660 2507 8676 2571
rect 8740 2507 8882 2571
rect 8946 2507 8962 2571
rect 9026 2507 9042 2571
rect 9106 2507 9122 2571
rect 9186 2507 9202 2571
rect 9266 2507 9282 2571
rect 9346 2507 9488 2571
rect 9552 2507 9568 2571
rect 9632 2507 9648 2571
rect 9712 2507 9728 2571
rect 9792 2507 9808 2571
rect 9872 2507 9888 2571
rect 9952 2507 10094 2571
rect 10158 2507 10174 2571
rect 10238 2507 10254 2571
rect 10318 2507 10334 2571
rect 10398 2507 10414 2571
rect 10478 2507 10494 2571
rect 10558 2507 10700 2571
rect 10764 2507 10780 2571
rect 10844 2507 10860 2571
rect 10924 2507 10940 2571
rect 11004 2507 11020 2571
rect 11084 2507 11100 2571
rect 11164 2507 11306 2571
rect 11370 2507 11386 2571
rect 11450 2507 11466 2571
rect 11530 2507 11546 2571
rect 11610 2507 11626 2571
rect 11690 2507 11706 2571
rect 11770 2507 11912 2571
rect 11976 2507 11992 2571
rect 12056 2507 12072 2571
rect 12136 2507 12152 2571
rect 12216 2507 12232 2571
rect 12296 2507 12312 2571
rect 12376 2507 12518 2571
rect 12582 2507 12598 2571
rect 12662 2507 12678 2571
rect 12742 2507 12758 2571
rect 12822 2507 12838 2571
rect 12902 2507 12918 2571
rect 12982 2507 13086 2571
rect 8172 2505 13086 2507
rect 13146 2550 13344 2560
rect 7440 2502 8112 2504
rect 13146 2486 13267 2550
rect 13331 2486 13344 2550
rect 13146 2476 13344 2486
rect 7791 2323 8463 2325
rect 7791 2259 7895 2323
rect 7959 2259 7975 2323
rect 8039 2259 8055 2323
rect 8119 2259 8135 2323
rect 8199 2259 8215 2323
rect 8279 2259 8295 2323
rect 8359 2259 8463 2323
rect 7791 2257 8463 2259
rect 7791 2103 7857 2257
rect 7791 2039 7792 2103
rect 7856 2039 7857 2103
rect 7791 2023 7857 2039
rect 7791 1959 7792 2023
rect 7856 1959 7857 2023
rect 7791 1943 7857 1959
rect 7791 1879 7792 1943
rect 7856 1879 7857 1943
rect 7791 1863 7857 1879
rect 7791 1799 7792 1863
rect 7856 1799 7857 1863
rect 7791 1783 7857 1799
rect 7791 1719 7792 1783
rect 7856 1719 7857 1783
rect 7791 1703 7857 1719
rect 7791 1639 7792 1703
rect 7856 1639 7857 1703
rect 7791 1623 7857 1639
rect 7791 1559 7792 1623
rect 7856 1559 7857 1623
rect 7791 1543 7857 1559
rect 7791 1479 7792 1543
rect 7856 1479 7857 1543
rect 7791 1463 7857 1479
rect 7791 1399 7792 1463
rect 7856 1399 7857 1463
rect 7791 1383 7857 1399
rect 7791 1319 7792 1383
rect 7856 1319 7857 1383
rect 7791 1229 7857 1319
rect 7917 1563 7977 2195
rect 8037 1563 8097 2257
rect 7917 1487 8097 1563
rect 7403 1164 7528 1170
rect 7917 1165 7977 1487
rect 8037 1225 8097 1487
rect 8157 1165 8217 2195
rect 8277 1225 8337 2257
rect 8397 2103 8463 2257
rect 8397 2039 8398 2103
rect 8462 2039 8463 2103
rect 8397 2023 8463 2039
rect 8397 1959 8398 2023
rect 8462 1959 8463 2023
rect 8397 1943 8463 1959
rect 8397 1879 8398 1943
rect 8462 1879 8463 1943
rect 8397 1863 8463 1879
rect 8397 1799 8398 1863
rect 8462 1799 8463 1863
rect 8397 1783 8463 1799
rect 8397 1719 8398 1783
rect 8462 1719 8463 1783
rect 8397 1703 8463 1719
rect 8397 1639 8398 1703
rect 8462 1639 8463 1703
rect 8397 1623 8463 1639
rect 8397 1559 8398 1623
rect 8462 1559 8463 1623
rect 8397 1543 8463 1559
rect 8397 1479 8398 1543
rect 8462 1479 8463 1543
rect 8397 1463 8463 1479
rect 8397 1399 8398 1463
rect 8462 1399 8463 1463
rect 8397 1383 8463 1399
rect 8397 1319 8398 1383
rect 8462 1319 8463 1383
rect 8397 1229 8463 1319
rect 8523 2323 11013 2325
rect 8523 2259 8627 2323
rect 8691 2259 8707 2323
rect 8771 2259 8787 2323
rect 8851 2259 8867 2323
rect 8931 2259 8947 2323
rect 9011 2259 9027 2323
rect 9091 2259 9233 2323
rect 9297 2259 9313 2323
rect 9377 2259 9393 2323
rect 9457 2259 9473 2323
rect 9537 2259 9553 2323
rect 9617 2259 9633 2323
rect 9697 2259 9839 2323
rect 9903 2259 9919 2323
rect 9983 2259 9999 2323
rect 10063 2259 10079 2323
rect 10143 2259 10159 2323
rect 10223 2259 10239 2323
rect 10303 2259 10445 2323
rect 10509 2259 10525 2323
rect 10589 2259 10605 2323
rect 10669 2259 10685 2323
rect 10749 2259 10765 2323
rect 10829 2259 10845 2323
rect 10909 2259 11013 2323
rect 8523 2257 11013 2259
rect 8523 2103 8589 2257
rect 8523 2039 8524 2103
rect 8588 2039 8589 2103
rect 8523 2023 8589 2039
rect 8523 1959 8524 2023
rect 8588 1959 8589 2023
rect 8523 1943 8589 1959
rect 8523 1879 8524 1943
rect 8588 1879 8589 1943
rect 8523 1863 8589 1879
rect 8523 1799 8524 1863
rect 8588 1799 8589 1863
rect 8523 1783 8589 1799
rect 8523 1719 8524 1783
rect 8588 1719 8589 1783
rect 8523 1703 8589 1719
rect 8523 1639 8524 1703
rect 8588 1639 8589 1703
rect 8523 1623 8589 1639
rect 8523 1559 8524 1623
rect 8588 1559 8589 1623
rect 8523 1543 8589 1559
rect 8523 1479 8524 1543
rect 8588 1479 8589 1543
rect 8523 1463 8589 1479
rect 8523 1399 8524 1463
rect 8588 1399 8589 1463
rect 8523 1383 8589 1399
rect 8523 1319 8524 1383
rect 8588 1319 8589 1383
rect 8523 1229 8589 1319
rect 8649 1563 8709 2195
rect 8769 1563 8829 2257
rect 8649 1487 8829 1563
rect 8649 1165 8709 1487
rect 8769 1225 8829 1487
rect 8889 1165 8949 2195
rect 9009 1225 9069 2257
rect 9129 2103 9195 2257
rect 9129 2039 9130 2103
rect 9194 2039 9195 2103
rect 9129 2023 9195 2039
rect 9129 1959 9130 2023
rect 9194 1959 9195 2023
rect 9129 1943 9195 1959
rect 9129 1879 9130 1943
rect 9194 1879 9195 1943
rect 9129 1863 9195 1879
rect 9129 1799 9130 1863
rect 9194 1799 9195 1863
rect 9129 1783 9195 1799
rect 9129 1719 9130 1783
rect 9194 1719 9195 1783
rect 9129 1703 9195 1719
rect 9129 1639 9130 1703
rect 9194 1639 9195 1703
rect 9129 1623 9195 1639
rect 9129 1559 9130 1623
rect 9194 1559 9195 1623
rect 9129 1543 9195 1559
rect 9129 1479 9130 1543
rect 9194 1479 9195 1543
rect 9129 1463 9195 1479
rect 9129 1399 9130 1463
rect 9194 1399 9195 1463
rect 9129 1383 9195 1399
rect 9129 1319 9130 1383
rect 9194 1319 9195 1383
rect 9129 1229 9195 1319
rect 9255 1225 9315 2257
rect 9375 1165 9435 2195
rect 9495 1563 9555 2257
rect 9615 1563 9675 2195
rect 9495 1487 9675 1563
rect 9495 1225 9555 1487
rect 9615 1165 9675 1487
rect 9735 2103 9801 2257
rect 9735 2039 9736 2103
rect 9800 2039 9801 2103
rect 9735 2023 9801 2039
rect 9735 1959 9736 2023
rect 9800 1959 9801 2023
rect 9735 1943 9801 1959
rect 9735 1879 9736 1943
rect 9800 1879 9801 1943
rect 9735 1863 9801 1879
rect 9735 1799 9736 1863
rect 9800 1799 9801 1863
rect 9735 1783 9801 1799
rect 9735 1719 9736 1783
rect 9800 1719 9801 1783
rect 9735 1703 9801 1719
rect 9735 1639 9736 1703
rect 9800 1639 9801 1703
rect 9735 1623 9801 1639
rect 9735 1559 9736 1623
rect 9800 1559 9801 1623
rect 9735 1543 9801 1559
rect 9735 1479 9736 1543
rect 9800 1479 9801 1543
rect 9735 1463 9801 1479
rect 9735 1399 9736 1463
rect 9800 1399 9801 1463
rect 9735 1383 9801 1399
rect 9735 1319 9736 1383
rect 9800 1319 9801 1383
rect 9735 1229 9801 1319
rect 9861 1563 9921 2195
rect 9981 1563 10041 2257
rect 9861 1487 10041 1563
rect 9861 1165 9921 1487
rect 9981 1225 10041 1487
rect 10101 1165 10161 2195
rect 10221 1225 10281 2257
rect 10341 2103 10407 2257
rect 10341 2039 10342 2103
rect 10406 2039 10407 2103
rect 10341 2023 10407 2039
rect 10341 1959 10342 2023
rect 10406 1959 10407 2023
rect 10341 1943 10407 1959
rect 10341 1879 10342 1943
rect 10406 1879 10407 1943
rect 10341 1863 10407 1879
rect 10341 1799 10342 1863
rect 10406 1799 10407 1863
rect 10341 1783 10407 1799
rect 10341 1719 10342 1783
rect 10406 1719 10407 1783
rect 10341 1703 10407 1719
rect 10341 1639 10342 1703
rect 10406 1639 10407 1703
rect 10341 1623 10407 1639
rect 10341 1559 10342 1623
rect 10406 1559 10407 1623
rect 10341 1543 10407 1559
rect 10341 1479 10342 1543
rect 10406 1479 10407 1543
rect 10341 1463 10407 1479
rect 10341 1399 10342 1463
rect 10406 1399 10407 1463
rect 10341 1383 10407 1399
rect 10341 1319 10342 1383
rect 10406 1319 10407 1383
rect 10341 1229 10407 1319
rect 10467 1225 10527 2257
rect 10587 1165 10647 2195
rect 10707 1563 10767 2257
rect 10827 1563 10887 2195
rect 10707 1487 10887 1563
rect 10707 1225 10767 1487
rect 10827 1165 10887 1487
rect 10947 2103 11013 2257
rect 10947 2039 10948 2103
rect 11012 2039 11013 2103
rect 10947 2023 11013 2039
rect 10947 1959 10948 2023
rect 11012 1959 11013 2023
rect 10947 1943 11013 1959
rect 10947 1879 10948 1943
rect 11012 1879 11013 1943
rect 10947 1863 11013 1879
rect 10947 1799 10948 1863
rect 11012 1799 11013 1863
rect 10947 1783 11013 1799
rect 10947 1719 10948 1783
rect 11012 1719 11013 1783
rect 10947 1703 11013 1719
rect 10947 1639 10948 1703
rect 11012 1639 11013 1703
rect 10947 1623 11013 1639
rect 10947 1559 10948 1623
rect 11012 1559 11013 1623
rect 10947 1543 11013 1559
rect 10947 1479 10948 1543
rect 11012 1479 11013 1543
rect 10947 1463 11013 1479
rect 10947 1399 10948 1463
rect 11012 1399 11013 1463
rect 10947 1383 11013 1399
rect 10947 1319 10948 1383
rect 11012 1319 11013 1383
rect 10947 1229 11013 1319
rect 11073 2323 12351 2325
rect 11073 2259 11177 2323
rect 11241 2259 11257 2323
rect 11321 2259 11337 2323
rect 11401 2259 11417 2323
rect 11481 2259 11497 2323
rect 11561 2259 11577 2323
rect 11641 2259 11783 2323
rect 11847 2259 11863 2323
rect 11927 2259 11943 2323
rect 12007 2259 12023 2323
rect 12087 2259 12103 2323
rect 12167 2259 12183 2323
rect 12247 2259 12351 2323
rect 11073 2257 12351 2259
rect 11073 2103 11139 2257
rect 11073 2039 11074 2103
rect 11138 2039 11139 2103
rect 11073 2023 11139 2039
rect 11073 1959 11074 2023
rect 11138 1959 11139 2023
rect 11073 1943 11139 1959
rect 11073 1879 11074 1943
rect 11138 1879 11139 1943
rect 11073 1863 11139 1879
rect 11073 1799 11074 1863
rect 11138 1799 11139 1863
rect 11073 1783 11139 1799
rect 11073 1719 11074 1783
rect 11138 1719 11139 1783
rect 11073 1703 11139 1719
rect 11073 1639 11074 1703
rect 11138 1639 11139 1703
rect 11073 1623 11139 1639
rect 11073 1559 11074 1623
rect 11138 1559 11139 1623
rect 11073 1543 11139 1559
rect 11073 1479 11074 1543
rect 11138 1479 11139 1543
rect 11073 1463 11139 1479
rect 11073 1399 11074 1463
rect 11138 1399 11139 1463
rect 11073 1383 11139 1399
rect 11073 1319 11074 1383
rect 11138 1319 11139 1383
rect 11073 1229 11139 1319
rect 11199 1563 11259 2195
rect 11319 1563 11379 2257
rect 11199 1487 11379 1563
rect 11199 1165 11259 1487
rect 11319 1225 11379 1487
rect 11439 1165 11499 2195
rect 11559 1225 11619 2257
rect 11679 2103 11745 2257
rect 11679 2039 11680 2103
rect 11744 2039 11745 2103
rect 11679 2023 11745 2039
rect 11679 1959 11680 2023
rect 11744 1959 11745 2023
rect 11679 1943 11745 1959
rect 11679 1879 11680 1943
rect 11744 1879 11745 1943
rect 11679 1863 11745 1879
rect 11679 1799 11680 1863
rect 11744 1799 11745 1863
rect 11679 1783 11745 1799
rect 11679 1719 11680 1783
rect 11744 1719 11745 1783
rect 11679 1703 11745 1719
rect 11679 1639 11680 1703
rect 11744 1639 11745 1703
rect 11679 1623 11745 1639
rect 11679 1559 11680 1623
rect 11744 1559 11745 1623
rect 11679 1543 11745 1559
rect 11679 1479 11680 1543
rect 11744 1479 11745 1543
rect 11679 1463 11745 1479
rect 11679 1399 11680 1463
rect 11744 1399 11745 1463
rect 11679 1383 11745 1399
rect 11679 1319 11680 1383
rect 11744 1319 11745 1383
rect 11679 1229 11745 1319
rect 11805 1225 11865 2257
rect 11925 1165 11985 2195
rect 12045 1563 12105 2257
rect 12165 1563 12225 2195
rect 12045 1487 12225 1563
rect 12045 1225 12105 1487
rect 12165 1165 12225 1487
rect 12285 2103 12351 2257
rect 12285 2039 12286 2103
rect 12350 2039 12351 2103
rect 12285 2023 12351 2039
rect 12285 1959 12286 2023
rect 12350 1959 12351 2023
rect 12285 1943 12351 1959
rect 12285 1879 12286 1943
rect 12350 1879 12351 1943
rect 12285 1863 12351 1879
rect 12285 1799 12286 1863
rect 12350 1799 12351 1863
rect 12285 1783 12351 1799
rect 12285 1719 12286 1783
rect 12350 1719 12351 1783
rect 12285 1703 12351 1719
rect 12285 1639 12286 1703
rect 12350 1639 12351 1703
rect 12285 1623 12351 1639
rect 12285 1559 12286 1623
rect 12350 1559 12351 1623
rect 12285 1543 12351 1559
rect 12285 1479 12286 1543
rect 12350 1479 12351 1543
rect 12285 1463 12351 1479
rect 12285 1399 12286 1463
rect 12350 1399 12351 1463
rect 12285 1383 12351 1399
rect 12285 1319 12286 1383
rect 12350 1319 12351 1383
rect 12285 1229 12351 1319
rect 12413 2323 13085 2325
rect 12413 2259 12517 2323
rect 12581 2259 12597 2323
rect 12661 2259 12677 2323
rect 12741 2259 12757 2323
rect 12821 2259 12837 2323
rect 12901 2259 12917 2323
rect 12981 2259 13085 2323
rect 12413 2257 13085 2259
rect 12413 2103 12479 2257
rect 12413 2039 12414 2103
rect 12478 2039 12479 2103
rect 12413 2023 12479 2039
rect 12413 1959 12414 2023
rect 12478 1959 12479 2023
rect 12413 1943 12479 1959
rect 12413 1879 12414 1943
rect 12478 1879 12479 1943
rect 12413 1863 12479 1879
rect 12413 1799 12414 1863
rect 12478 1799 12479 1863
rect 12413 1783 12479 1799
rect 12413 1719 12414 1783
rect 12478 1719 12479 1783
rect 12413 1703 12479 1719
rect 12413 1639 12414 1703
rect 12478 1639 12479 1703
rect 12413 1623 12479 1639
rect 12413 1559 12414 1623
rect 12478 1559 12479 1623
rect 12413 1543 12479 1559
rect 12413 1479 12414 1543
rect 12478 1479 12479 1543
rect 12413 1463 12479 1479
rect 12413 1399 12414 1463
rect 12478 1399 12479 1463
rect 12413 1383 12479 1399
rect 12413 1319 12414 1383
rect 12478 1319 12479 1383
rect 12413 1229 12479 1319
rect 12539 1225 12599 2257
rect 12659 1165 12719 2195
rect 12779 1563 12839 2257
rect 12899 1563 12959 2195
rect 12779 1487 12959 1563
rect 12779 1225 12839 1487
rect 12899 1165 12959 1487
rect 13019 2103 13085 2257
rect 13019 2039 13020 2103
rect 13084 2039 13085 2103
rect 13019 2023 13085 2039
rect 13019 1959 13020 2023
rect 13084 1959 13085 2023
rect 13019 1943 13085 1959
rect 13019 1879 13020 1943
rect 13084 1879 13085 1943
rect 13019 1863 13085 1879
rect 13019 1799 13020 1863
rect 13084 1799 13085 1863
rect 13019 1783 13085 1799
rect 13019 1719 13020 1783
rect 13084 1719 13085 1783
rect 13019 1703 13085 1719
rect 13019 1639 13020 1703
rect 13084 1639 13085 1703
rect 13019 1623 13085 1639
rect 13019 1559 13020 1623
rect 13084 1559 13085 1623
rect 13019 1543 13085 1559
rect 13019 1479 13020 1543
rect 13084 1479 13085 1543
rect 13019 1463 13085 1479
rect 13019 1399 13020 1463
rect 13084 1399 13085 1463
rect 13019 1383 13085 1399
rect 13019 1319 13020 1383
rect 13084 1319 13085 1383
rect 13019 1229 13085 1319
rect 13146 2095 13206 2476
rect 13404 2357 13464 2735
rect 13266 2347 13464 2357
rect 13266 2283 13267 2347
rect 13331 2283 13464 2347
rect 13266 2273 13464 2283
rect 13146 2085 13464 2095
rect 13146 2021 13176 2085
rect 13240 2021 13464 2085
rect 7791 1164 8463 1165
rect 8523 1164 11013 1165
rect 11073 1164 12351 1165
rect 12413 1164 13085 1165
rect 13146 1164 13464 2021
rect 6843 1163 13464 1164
rect 6843 1160 7975 1163
rect 6843 1150 7433 1160
rect 6192 1099 7433 1150
rect 788 1096 7433 1099
rect 7497 1099 7975 1160
rect 8039 1099 8055 1163
rect 8119 1099 8135 1163
rect 8199 1099 8215 1163
rect 8279 1099 8707 1163
rect 8771 1099 8787 1163
rect 8851 1099 8867 1163
rect 8931 1099 8947 1163
rect 9011 1099 9313 1163
rect 9377 1099 9393 1163
rect 9457 1099 9473 1163
rect 9537 1099 9553 1163
rect 9617 1099 9919 1163
rect 9983 1099 9999 1163
rect 10063 1099 10079 1163
rect 10143 1099 10159 1163
rect 10223 1099 10525 1163
rect 10589 1099 10605 1163
rect 10669 1099 10685 1163
rect 10749 1099 10765 1163
rect 10829 1099 11257 1163
rect 11321 1099 11337 1163
rect 11401 1099 11417 1163
rect 11481 1099 11497 1163
rect 11561 1099 11863 1163
rect 11927 1099 11943 1163
rect 12007 1099 12023 1163
rect 12087 1099 12103 1163
rect 12167 1099 12597 1163
rect 12661 1099 12677 1163
rect 12741 1099 12757 1163
rect 12821 1099 12837 1163
rect 12901 1099 13464 1163
rect 7497 1096 13464 1099
rect 3 1047 13464 1096
rect 4 867 13464 1047
rect 4 483 933 867
rect 2237 483 2772 867
rect 3884 483 4284 867
rect 5779 866 13464 867
rect 5779 503 7001 866
rect 8138 503 8727 866
rect 9605 503 10116 866
rect 11111 503 11641 866
rect 12555 503 13464 866
rect 5779 483 13464 503
rect 4 256 13464 483
rect 3 235 13464 256
rect 0 225 13464 235
rect 0 222 5967 225
rect 0 158 563 222
rect 627 158 643 222
rect 707 158 723 222
rect 787 158 803 222
rect 867 158 1297 222
rect 1361 158 1377 222
rect 1441 158 1457 222
rect 1521 158 1537 222
rect 1601 158 1903 222
rect 1967 158 1983 222
rect 2047 158 2063 222
rect 2127 158 2143 222
rect 2207 158 2635 222
rect 2699 158 2715 222
rect 2779 158 2795 222
rect 2859 158 2875 222
rect 2939 158 3241 222
rect 3305 158 3321 222
rect 3385 158 3401 222
rect 3465 158 3481 222
rect 3545 158 3847 222
rect 3911 158 3927 222
rect 3991 158 4007 222
rect 4071 158 4087 222
rect 4151 158 4453 222
rect 4517 158 4533 222
rect 4597 158 4613 222
rect 4677 158 4693 222
rect 4757 158 5185 222
rect 5249 158 5265 222
rect 5329 158 5345 222
rect 5409 158 5425 222
rect 5489 161 5967 222
rect 6031 222 12676 225
rect 6031 217 7272 222
rect 6031 161 6621 217
rect 5489 158 6621 161
rect 0 157 6621 158
rect 0 -700 318 157
rect 379 156 1051 157
rect 1113 156 2391 157
rect 2451 156 4941 157
rect 5001 156 5673 157
rect 0 -764 224 -700
rect 288 -764 318 -700
rect 0 -774 318 -764
rect 0 -962 198 -952
rect 0 -1026 133 -962
rect 197 -1026 198 -962
rect 0 -1036 198 -1026
rect 0 -1414 60 -1036
rect 258 -1155 318 -774
rect 379 2 445 92
rect 379 -62 380 2
rect 444 -62 445 2
rect 379 -78 445 -62
rect 379 -142 380 -78
rect 444 -142 445 -78
rect 379 -158 445 -142
rect 379 -222 380 -158
rect 444 -222 445 -158
rect 379 -238 445 -222
rect 379 -302 380 -238
rect 444 -302 445 -238
rect 379 -318 445 -302
rect 379 -382 380 -318
rect 444 -382 445 -318
rect 379 -398 445 -382
rect 379 -462 380 -398
rect 444 -462 445 -398
rect 379 -478 445 -462
rect 379 -542 380 -478
rect 444 -542 445 -478
rect 379 -558 445 -542
rect 379 -622 380 -558
rect 444 -622 445 -558
rect 379 -638 445 -622
rect 379 -702 380 -638
rect 444 -702 445 -638
rect 379 -718 445 -702
rect 379 -782 380 -718
rect 444 -782 445 -718
rect 379 -936 445 -782
rect 505 -166 565 156
rect 625 -166 685 96
rect 505 -242 685 -166
rect 505 -874 565 -242
rect 625 -936 685 -242
rect 745 -874 805 156
rect 865 -936 925 96
rect 985 2 1051 92
rect 985 -62 986 2
rect 1050 -62 1051 2
rect 985 -78 1051 -62
rect 985 -142 986 -78
rect 1050 -142 1051 -78
rect 985 -158 1051 -142
rect 985 -222 986 -158
rect 1050 -222 1051 -158
rect 985 -238 1051 -222
rect 985 -302 986 -238
rect 1050 -302 1051 -238
rect 985 -318 1051 -302
rect 985 -382 986 -318
rect 1050 -382 1051 -318
rect 985 -398 1051 -382
rect 985 -462 986 -398
rect 1050 -462 1051 -398
rect 985 -478 1051 -462
rect 985 -542 986 -478
rect 1050 -542 1051 -478
rect 985 -558 1051 -542
rect 985 -622 986 -558
rect 1050 -622 1051 -558
rect 985 -638 1051 -622
rect 985 -702 986 -638
rect 1050 -702 1051 -638
rect 985 -718 1051 -702
rect 985 -782 986 -718
rect 1050 -782 1051 -718
rect 985 -936 1051 -782
rect 379 -938 1051 -936
rect 379 -1002 483 -938
rect 547 -1002 563 -938
rect 627 -1002 643 -938
rect 707 -1002 723 -938
rect 787 -1002 803 -938
rect 867 -1002 883 -938
rect 947 -1002 1051 -938
rect 379 -1004 1051 -1002
rect 1113 2 1179 92
rect 1113 -62 1114 2
rect 1178 -62 1179 2
rect 1113 -78 1179 -62
rect 1113 -142 1114 -78
rect 1178 -142 1179 -78
rect 1113 -158 1179 -142
rect 1113 -222 1114 -158
rect 1178 -222 1179 -158
rect 1113 -238 1179 -222
rect 1113 -302 1114 -238
rect 1178 -302 1179 -238
rect 1113 -318 1179 -302
rect 1113 -382 1114 -318
rect 1178 -382 1179 -318
rect 1113 -398 1179 -382
rect 1113 -462 1114 -398
rect 1178 -462 1179 -398
rect 1113 -478 1179 -462
rect 1113 -542 1114 -478
rect 1178 -542 1179 -478
rect 1113 -558 1179 -542
rect 1113 -622 1114 -558
rect 1178 -622 1179 -558
rect 1113 -638 1179 -622
rect 1113 -702 1114 -638
rect 1178 -702 1179 -638
rect 1113 -718 1179 -702
rect 1113 -782 1114 -718
rect 1178 -782 1179 -718
rect 1113 -936 1179 -782
rect 1239 -166 1299 156
rect 1359 -166 1419 96
rect 1239 -242 1419 -166
rect 1239 -874 1299 -242
rect 1359 -936 1419 -242
rect 1479 -874 1539 156
rect 1599 -936 1659 96
rect 1719 2 1785 92
rect 1719 -62 1720 2
rect 1784 -62 1785 2
rect 1719 -78 1785 -62
rect 1719 -142 1720 -78
rect 1784 -142 1785 -78
rect 1719 -158 1785 -142
rect 1719 -222 1720 -158
rect 1784 -222 1785 -158
rect 1719 -238 1785 -222
rect 1719 -302 1720 -238
rect 1784 -302 1785 -238
rect 1719 -318 1785 -302
rect 1719 -382 1720 -318
rect 1784 -382 1785 -318
rect 1719 -398 1785 -382
rect 1719 -462 1720 -398
rect 1784 -462 1785 -398
rect 1719 -478 1785 -462
rect 1719 -542 1720 -478
rect 1784 -542 1785 -478
rect 1719 -558 1785 -542
rect 1719 -622 1720 -558
rect 1784 -622 1785 -558
rect 1719 -638 1785 -622
rect 1719 -702 1720 -638
rect 1784 -702 1785 -638
rect 1719 -718 1785 -702
rect 1719 -782 1720 -718
rect 1784 -782 1785 -718
rect 1719 -936 1785 -782
rect 1845 -936 1905 96
rect 1965 -874 2025 156
rect 2085 -166 2145 96
rect 2205 -166 2265 156
rect 2085 -242 2265 -166
rect 2085 -936 2145 -242
rect 2205 -874 2265 -242
rect 2325 2 2391 92
rect 2325 -62 2326 2
rect 2390 -62 2391 2
rect 2325 -78 2391 -62
rect 2325 -142 2326 -78
rect 2390 -142 2391 -78
rect 2325 -158 2391 -142
rect 2325 -222 2326 -158
rect 2390 -222 2391 -158
rect 2325 -238 2391 -222
rect 2325 -302 2326 -238
rect 2390 -302 2391 -238
rect 2325 -318 2391 -302
rect 2325 -382 2326 -318
rect 2390 -382 2391 -318
rect 2325 -398 2391 -382
rect 2325 -462 2326 -398
rect 2390 -462 2391 -398
rect 2325 -478 2391 -462
rect 2325 -542 2326 -478
rect 2390 -542 2391 -478
rect 2325 -558 2391 -542
rect 2325 -622 2326 -558
rect 2390 -622 2391 -558
rect 2325 -638 2391 -622
rect 2325 -702 2326 -638
rect 2390 -702 2391 -638
rect 2325 -718 2391 -702
rect 2325 -782 2326 -718
rect 2390 -782 2391 -718
rect 2325 -936 2391 -782
rect 1113 -938 2391 -936
rect 1113 -1002 1217 -938
rect 1281 -1002 1297 -938
rect 1361 -1002 1377 -938
rect 1441 -1002 1457 -938
rect 1521 -1002 1537 -938
rect 1601 -1002 1617 -938
rect 1681 -1002 1823 -938
rect 1887 -1002 1903 -938
rect 1967 -1002 1983 -938
rect 2047 -1002 2063 -938
rect 2127 -1002 2143 -938
rect 2207 -1002 2223 -938
rect 2287 -1002 2391 -938
rect 1113 -1004 2391 -1002
rect 2451 2 2517 92
rect 2451 -62 2452 2
rect 2516 -62 2517 2
rect 2451 -78 2517 -62
rect 2451 -142 2452 -78
rect 2516 -142 2517 -78
rect 2451 -158 2517 -142
rect 2451 -222 2452 -158
rect 2516 -222 2517 -158
rect 2451 -238 2517 -222
rect 2451 -302 2452 -238
rect 2516 -302 2517 -238
rect 2451 -318 2517 -302
rect 2451 -382 2452 -318
rect 2516 -382 2517 -318
rect 2451 -398 2517 -382
rect 2451 -462 2452 -398
rect 2516 -462 2517 -398
rect 2451 -478 2517 -462
rect 2451 -542 2452 -478
rect 2516 -542 2517 -478
rect 2451 -558 2517 -542
rect 2451 -622 2452 -558
rect 2516 -622 2517 -558
rect 2451 -638 2517 -622
rect 2451 -702 2452 -638
rect 2516 -702 2517 -638
rect 2451 -718 2517 -702
rect 2451 -782 2452 -718
rect 2516 -782 2517 -718
rect 2451 -936 2517 -782
rect 2577 -166 2637 156
rect 2697 -166 2757 96
rect 2577 -242 2757 -166
rect 2577 -874 2637 -242
rect 2697 -936 2757 -242
rect 2817 -874 2877 156
rect 2937 -936 2997 96
rect 3057 2 3123 92
rect 3057 -62 3058 2
rect 3122 -62 3123 2
rect 3057 -78 3123 -62
rect 3057 -142 3058 -78
rect 3122 -142 3123 -78
rect 3057 -158 3123 -142
rect 3057 -222 3058 -158
rect 3122 -222 3123 -158
rect 3057 -238 3123 -222
rect 3057 -302 3058 -238
rect 3122 -302 3123 -238
rect 3057 -318 3123 -302
rect 3057 -382 3058 -318
rect 3122 -382 3123 -318
rect 3057 -398 3123 -382
rect 3057 -462 3058 -398
rect 3122 -462 3123 -398
rect 3057 -478 3123 -462
rect 3057 -542 3058 -478
rect 3122 -542 3123 -478
rect 3057 -558 3123 -542
rect 3057 -622 3058 -558
rect 3122 -622 3123 -558
rect 3057 -638 3123 -622
rect 3057 -702 3058 -638
rect 3122 -702 3123 -638
rect 3057 -718 3123 -702
rect 3057 -782 3058 -718
rect 3122 -782 3123 -718
rect 3057 -936 3123 -782
rect 3183 -936 3243 96
rect 3303 -874 3363 156
rect 3423 -166 3483 96
rect 3543 -166 3603 156
rect 3423 -242 3603 -166
rect 3423 -936 3483 -242
rect 3543 -874 3603 -242
rect 3663 2 3729 92
rect 3663 -62 3664 2
rect 3728 -62 3729 2
rect 3663 -78 3729 -62
rect 3663 -142 3664 -78
rect 3728 -142 3729 -78
rect 3663 -158 3729 -142
rect 3663 -222 3664 -158
rect 3728 -222 3729 -158
rect 3663 -238 3729 -222
rect 3663 -302 3664 -238
rect 3728 -302 3729 -238
rect 3663 -318 3729 -302
rect 3663 -382 3664 -318
rect 3728 -382 3729 -318
rect 3663 -398 3729 -382
rect 3663 -462 3664 -398
rect 3728 -462 3729 -398
rect 3663 -478 3729 -462
rect 3663 -542 3664 -478
rect 3728 -542 3729 -478
rect 3663 -558 3729 -542
rect 3663 -622 3664 -558
rect 3728 -622 3729 -558
rect 3663 -638 3729 -622
rect 3663 -702 3664 -638
rect 3728 -702 3729 -638
rect 3663 -718 3729 -702
rect 3663 -782 3664 -718
rect 3728 -782 3729 -718
rect 3663 -936 3729 -782
rect 3789 -166 3849 156
rect 3909 -166 3969 96
rect 3789 -242 3969 -166
rect 3789 -874 3849 -242
rect 3909 -936 3969 -242
rect 4029 -874 4089 156
rect 4149 -936 4209 96
rect 4269 2 4335 92
rect 4269 -62 4270 2
rect 4334 -62 4335 2
rect 4269 -78 4335 -62
rect 4269 -142 4270 -78
rect 4334 -142 4335 -78
rect 4269 -158 4335 -142
rect 4269 -222 4270 -158
rect 4334 -222 4335 -158
rect 4269 -238 4335 -222
rect 4269 -302 4270 -238
rect 4334 -302 4335 -238
rect 4269 -318 4335 -302
rect 4269 -382 4270 -318
rect 4334 -382 4335 -318
rect 4269 -398 4335 -382
rect 4269 -462 4270 -398
rect 4334 -462 4335 -398
rect 4269 -478 4335 -462
rect 4269 -542 4270 -478
rect 4334 -542 4335 -478
rect 4269 -558 4335 -542
rect 4269 -622 4270 -558
rect 4334 -622 4335 -558
rect 4269 -638 4335 -622
rect 4269 -702 4270 -638
rect 4334 -702 4335 -638
rect 4269 -718 4335 -702
rect 4269 -782 4270 -718
rect 4334 -782 4335 -718
rect 4269 -936 4335 -782
rect 4395 -936 4455 96
rect 4515 -874 4575 156
rect 4635 -166 4695 96
rect 4755 -166 4815 156
rect 4635 -242 4815 -166
rect 4635 -936 4695 -242
rect 4755 -874 4815 -242
rect 4875 2 4941 92
rect 4875 -62 4876 2
rect 4940 -62 4941 2
rect 4875 -78 4941 -62
rect 4875 -142 4876 -78
rect 4940 -142 4941 -78
rect 4875 -158 4941 -142
rect 4875 -222 4876 -158
rect 4940 -222 4941 -158
rect 4875 -238 4941 -222
rect 4875 -302 4876 -238
rect 4940 -302 4941 -238
rect 4875 -318 4941 -302
rect 4875 -382 4876 -318
rect 4940 -382 4941 -318
rect 4875 -398 4941 -382
rect 4875 -462 4876 -398
rect 4940 -462 4941 -398
rect 4875 -478 4941 -462
rect 4875 -542 4876 -478
rect 4940 -542 4941 -478
rect 4875 -558 4941 -542
rect 4875 -622 4876 -558
rect 4940 -622 4941 -558
rect 4875 -638 4941 -622
rect 4875 -702 4876 -638
rect 4940 -702 4941 -638
rect 4875 -718 4941 -702
rect 4875 -782 4876 -718
rect 4940 -782 4941 -718
rect 4875 -936 4941 -782
rect 2451 -938 4941 -936
rect 2451 -1002 2555 -938
rect 2619 -1002 2635 -938
rect 2699 -1002 2715 -938
rect 2779 -1002 2795 -938
rect 2859 -1002 2875 -938
rect 2939 -1002 2955 -938
rect 3019 -1002 3161 -938
rect 3225 -1002 3241 -938
rect 3305 -1002 3321 -938
rect 3385 -1002 3401 -938
rect 3465 -1002 3481 -938
rect 3545 -1002 3561 -938
rect 3625 -1002 3767 -938
rect 3831 -1002 3847 -938
rect 3911 -1002 3927 -938
rect 3991 -1002 4007 -938
rect 4071 -1002 4087 -938
rect 4151 -1002 4167 -938
rect 4231 -1002 4373 -938
rect 4437 -1002 4453 -938
rect 4517 -1002 4533 -938
rect 4597 -1002 4613 -938
rect 4677 -1002 4693 -938
rect 4757 -1002 4773 -938
rect 4837 -1002 4941 -938
rect 2451 -1004 4941 -1002
rect 5001 2 5067 92
rect 5001 -62 5002 2
rect 5066 -62 5067 2
rect 5001 -78 5067 -62
rect 5001 -142 5002 -78
rect 5066 -142 5067 -78
rect 5001 -158 5067 -142
rect 5001 -222 5002 -158
rect 5066 -222 5067 -158
rect 5001 -238 5067 -222
rect 5001 -302 5002 -238
rect 5066 -302 5067 -238
rect 5001 -318 5067 -302
rect 5001 -382 5002 -318
rect 5066 -382 5067 -318
rect 5001 -398 5067 -382
rect 5001 -462 5002 -398
rect 5066 -462 5067 -398
rect 5001 -478 5067 -462
rect 5001 -542 5002 -478
rect 5066 -542 5067 -478
rect 5001 -558 5067 -542
rect 5001 -622 5002 -558
rect 5066 -622 5067 -558
rect 5001 -638 5067 -622
rect 5001 -702 5002 -638
rect 5066 -702 5067 -638
rect 5001 -718 5067 -702
rect 5001 -782 5002 -718
rect 5066 -782 5067 -718
rect 5001 -936 5067 -782
rect 5127 -936 5187 96
rect 5247 -874 5307 156
rect 5367 -166 5427 96
rect 5487 -166 5547 156
rect 5936 151 6061 157
rect 5367 -242 5547 -166
rect 5367 -936 5427 -242
rect 5487 -874 5547 -242
rect 5607 2 5673 92
rect 5607 -62 5608 2
rect 5672 -62 5673 2
rect 5607 -78 5673 -62
rect 5607 -142 5608 -78
rect 5672 -142 5673 -78
rect 5607 -158 5673 -142
rect 5607 -222 5608 -158
rect 5672 -222 5673 -158
rect 5607 -238 5673 -222
rect 5607 -302 5608 -238
rect 5672 -302 5673 -238
rect 5607 -318 5673 -302
rect 5607 -382 5608 -318
rect 5672 -382 5673 -318
rect 5607 -398 5673 -382
rect 5607 -462 5608 -398
rect 5672 -462 5673 -398
rect 5607 -478 5673 -462
rect 5607 -542 5608 -478
rect 5672 -542 5673 -478
rect 5607 -558 5673 -542
rect 5607 -622 5608 -558
rect 5672 -622 5673 -558
rect 5607 -638 5673 -622
rect 5607 -702 5608 -638
rect 5672 -702 5673 -638
rect 5607 -718 5673 -702
rect 5607 -782 5608 -718
rect 5672 -782 5673 -718
rect 5607 -936 5673 -782
rect 5001 -938 5673 -936
rect 5001 -1002 5105 -938
rect 5169 -1002 5185 -938
rect 5249 -1002 5265 -938
rect 5329 -1002 5345 -938
rect 5409 -1002 5425 -938
rect 5489 -1002 5505 -938
rect 5569 -1002 5673 -938
rect 5001 -1004 5673 -1002
rect 120 -1165 318 -1155
rect 120 -1229 133 -1165
rect 197 -1229 318 -1165
rect 5352 -1183 6024 -1181
rect 120 -1239 318 -1229
rect 378 -1186 5292 -1184
rect 378 -1250 482 -1186
rect 546 -1250 562 -1186
rect 626 -1250 642 -1186
rect 706 -1250 722 -1186
rect 786 -1250 802 -1186
rect 866 -1250 882 -1186
rect 946 -1250 1088 -1186
rect 1152 -1250 1168 -1186
rect 1232 -1250 1248 -1186
rect 1312 -1250 1328 -1186
rect 1392 -1250 1408 -1186
rect 1472 -1250 1488 -1186
rect 1552 -1250 1694 -1186
rect 1758 -1250 1774 -1186
rect 1838 -1250 1854 -1186
rect 1918 -1250 1934 -1186
rect 1998 -1250 2014 -1186
rect 2078 -1250 2094 -1186
rect 2158 -1250 2300 -1186
rect 2364 -1250 2380 -1186
rect 2444 -1250 2460 -1186
rect 2524 -1250 2540 -1186
rect 2604 -1250 2620 -1186
rect 2684 -1250 2700 -1186
rect 2764 -1250 2906 -1186
rect 2970 -1250 2986 -1186
rect 3050 -1250 3066 -1186
rect 3130 -1250 3146 -1186
rect 3210 -1250 3226 -1186
rect 3290 -1250 3306 -1186
rect 3370 -1250 3512 -1186
rect 3576 -1250 3592 -1186
rect 3656 -1250 3672 -1186
rect 3736 -1250 3752 -1186
rect 3816 -1250 3832 -1186
rect 3896 -1250 3912 -1186
rect 3976 -1250 4118 -1186
rect 4182 -1250 4198 -1186
rect 4262 -1250 4278 -1186
rect 4342 -1250 4358 -1186
rect 4422 -1250 4438 -1186
rect 4502 -1250 4518 -1186
rect 4582 -1250 4724 -1186
rect 4788 -1250 4804 -1186
rect 4868 -1250 4884 -1186
rect 4948 -1250 4964 -1186
rect 5028 -1250 5044 -1186
rect 5108 -1250 5124 -1186
rect 5188 -1250 5292 -1186
rect 378 -1252 5292 -1250
rect 378 -1406 444 -1252
rect 0 -1426 318 -1414
rect 0 -1490 221 -1426
rect 285 -1490 318 -1426
rect 0 -1668 318 -1490
rect 0 -1732 139 -1668
rect 203 -1732 318 -1668
rect 0 -1825 318 -1732
rect 0 -1889 138 -1825
rect 202 -1889 318 -1825
rect 0 -1995 318 -1889
rect 0 -2059 138 -1995
rect 202 -2059 318 -1995
rect 0 -2147 318 -2059
rect 0 -2211 139 -2147
rect 203 -2211 318 -2147
rect 0 -2291 318 -2211
rect 378 -1470 379 -1406
rect 443 -1470 444 -1406
rect 378 -1486 444 -1470
rect 378 -1550 379 -1486
rect 443 -1550 444 -1486
rect 378 -1566 444 -1550
rect 378 -1630 379 -1566
rect 443 -1630 444 -1566
rect 378 -1646 444 -1630
rect 378 -1710 379 -1646
rect 443 -1710 444 -1646
rect 378 -1726 444 -1710
rect 378 -1790 379 -1726
rect 443 -1790 444 -1726
rect 378 -1806 444 -1790
rect 378 -1870 379 -1806
rect 443 -1870 444 -1806
rect 378 -1886 444 -1870
rect 378 -1950 379 -1886
rect 443 -1950 444 -1886
rect 378 -1966 444 -1950
rect 378 -2030 379 -1966
rect 443 -2030 444 -1966
rect 378 -2046 444 -2030
rect 378 -2110 379 -2046
rect 443 -2110 444 -2046
rect 378 -2126 444 -2110
rect 378 -2190 379 -2126
rect 443 -2190 444 -2126
rect 378 -2280 444 -2190
rect 504 -1819 564 -1314
rect 624 -1819 684 -1252
rect 504 -1879 684 -1819
rect 0 -2355 144 -2291
rect 208 -2344 318 -2291
rect 504 -2344 564 -1879
rect 624 -2284 684 -1879
rect 744 -2344 804 -1314
rect 864 -2284 924 -1252
rect 984 -1406 1050 -1252
rect 984 -1470 985 -1406
rect 1049 -1470 1050 -1406
rect 984 -1486 1050 -1470
rect 984 -1550 985 -1486
rect 1049 -1550 1050 -1486
rect 984 -1566 1050 -1550
rect 984 -1630 985 -1566
rect 1049 -1630 1050 -1566
rect 984 -1646 1050 -1630
rect 984 -1710 985 -1646
rect 1049 -1710 1050 -1646
rect 984 -1726 1050 -1710
rect 984 -1790 985 -1726
rect 1049 -1790 1050 -1726
rect 984 -1806 1050 -1790
rect 984 -1870 985 -1806
rect 1049 -1870 1050 -1806
rect 984 -1886 1050 -1870
rect 984 -1950 985 -1886
rect 1049 -1950 1050 -1886
rect 984 -1966 1050 -1950
rect 984 -2030 985 -1966
rect 1049 -2030 1050 -1966
rect 984 -2046 1050 -2030
rect 984 -2110 985 -2046
rect 1049 -2110 1050 -2046
rect 984 -2126 1050 -2110
rect 984 -2190 985 -2126
rect 1049 -2190 1050 -2126
rect 984 -2280 1050 -2190
rect 1110 -2284 1170 -1252
rect 1230 -2344 1290 -1314
rect 1350 -1819 1410 -1252
rect 1470 -1819 1530 -1314
rect 1350 -1879 1530 -1819
rect 1350 -2284 1410 -1879
rect 1470 -2344 1530 -1879
rect 1590 -1406 1656 -1252
rect 1590 -1470 1591 -1406
rect 1655 -1470 1656 -1406
rect 1590 -1486 1656 -1470
rect 1590 -1550 1591 -1486
rect 1655 -1550 1656 -1486
rect 1590 -1566 1656 -1550
rect 1590 -1630 1591 -1566
rect 1655 -1630 1656 -1566
rect 1590 -1646 1656 -1630
rect 1590 -1710 1591 -1646
rect 1655 -1710 1656 -1646
rect 1590 -1726 1656 -1710
rect 1590 -1790 1591 -1726
rect 1655 -1790 1656 -1726
rect 1590 -1806 1656 -1790
rect 1590 -1870 1591 -1806
rect 1655 -1870 1656 -1806
rect 1590 -1886 1656 -1870
rect 1590 -1950 1591 -1886
rect 1655 -1950 1656 -1886
rect 1590 -1966 1656 -1950
rect 1590 -2030 1591 -1966
rect 1655 -2030 1656 -1966
rect 1590 -2046 1656 -2030
rect 1590 -2110 1591 -2046
rect 1655 -2110 1656 -2046
rect 1590 -2126 1656 -2110
rect 1590 -2190 1591 -2126
rect 1655 -2190 1656 -2126
rect 1590 -2280 1656 -2190
rect 1716 -1819 1776 -1314
rect 1836 -1819 1896 -1252
rect 1716 -1879 1896 -1819
rect 1716 -2344 1776 -1879
rect 1836 -2284 1896 -1879
rect 1956 -2344 2016 -1314
rect 2076 -2284 2136 -1252
rect 2196 -1406 2262 -1252
rect 2196 -1470 2197 -1406
rect 2261 -1470 2262 -1406
rect 2196 -1486 2262 -1470
rect 2196 -1550 2197 -1486
rect 2261 -1550 2262 -1486
rect 2196 -1566 2262 -1550
rect 2196 -1630 2197 -1566
rect 2261 -1630 2262 -1566
rect 2196 -1646 2262 -1630
rect 2196 -1710 2197 -1646
rect 2261 -1710 2262 -1646
rect 2196 -1726 2262 -1710
rect 2196 -1790 2197 -1726
rect 2261 -1790 2262 -1726
rect 2196 -1806 2262 -1790
rect 2196 -1870 2197 -1806
rect 2261 -1870 2262 -1806
rect 2196 -1886 2262 -1870
rect 2196 -1950 2197 -1886
rect 2261 -1950 2262 -1886
rect 2196 -1966 2262 -1950
rect 2196 -2030 2197 -1966
rect 2261 -2030 2262 -1966
rect 2196 -2046 2262 -2030
rect 2196 -2110 2197 -2046
rect 2261 -2110 2262 -2046
rect 2196 -2126 2262 -2110
rect 2196 -2190 2197 -2126
rect 2261 -2190 2262 -2126
rect 2196 -2280 2262 -2190
rect 2322 -2284 2382 -1252
rect 2442 -2344 2502 -1314
rect 2562 -1819 2622 -1252
rect 2682 -1819 2742 -1314
rect 2562 -1879 2742 -1819
rect 2562 -2284 2622 -1879
rect 2682 -2344 2742 -1879
rect 2802 -1406 2868 -1252
rect 2802 -1470 2803 -1406
rect 2867 -1470 2868 -1406
rect 2802 -1486 2868 -1470
rect 2802 -1550 2803 -1486
rect 2867 -1550 2868 -1486
rect 2802 -1566 2868 -1550
rect 2802 -1630 2803 -1566
rect 2867 -1630 2868 -1566
rect 2802 -1646 2868 -1630
rect 2802 -1710 2803 -1646
rect 2867 -1710 2868 -1646
rect 2802 -1726 2868 -1710
rect 2802 -1790 2803 -1726
rect 2867 -1790 2868 -1726
rect 2802 -1806 2868 -1790
rect 2802 -1870 2803 -1806
rect 2867 -1870 2868 -1806
rect 2802 -1886 2868 -1870
rect 2802 -1950 2803 -1886
rect 2867 -1950 2868 -1886
rect 2802 -1966 2868 -1950
rect 2802 -2030 2803 -1966
rect 2867 -2030 2868 -1966
rect 2802 -2046 2868 -2030
rect 2802 -2110 2803 -2046
rect 2867 -2110 2868 -2046
rect 2802 -2126 2868 -2110
rect 2802 -2190 2803 -2126
rect 2867 -2190 2868 -2126
rect 2802 -2280 2868 -2190
rect 2928 -1819 2988 -1314
rect 3048 -1819 3108 -1252
rect 2928 -1879 3108 -1819
rect 2928 -2344 2988 -1879
rect 3048 -2284 3108 -1879
rect 3168 -2344 3228 -1314
rect 3288 -2284 3348 -1252
rect 3408 -1406 3474 -1252
rect 3408 -1470 3409 -1406
rect 3473 -1470 3474 -1406
rect 3408 -1486 3474 -1470
rect 3408 -1550 3409 -1486
rect 3473 -1550 3474 -1486
rect 3408 -1566 3474 -1550
rect 3408 -1630 3409 -1566
rect 3473 -1630 3474 -1566
rect 3408 -1646 3474 -1630
rect 3408 -1710 3409 -1646
rect 3473 -1710 3474 -1646
rect 3408 -1726 3474 -1710
rect 3408 -1790 3409 -1726
rect 3473 -1790 3474 -1726
rect 3408 -1806 3474 -1790
rect 3408 -1870 3409 -1806
rect 3473 -1870 3474 -1806
rect 3408 -1886 3474 -1870
rect 3408 -1950 3409 -1886
rect 3473 -1950 3474 -1886
rect 3408 -1966 3474 -1950
rect 3408 -2030 3409 -1966
rect 3473 -2030 3474 -1966
rect 3408 -2046 3474 -2030
rect 3408 -2110 3409 -2046
rect 3473 -2110 3474 -2046
rect 3408 -2126 3474 -2110
rect 3408 -2190 3409 -2126
rect 3473 -2190 3474 -2126
rect 3408 -2280 3474 -2190
rect 3534 -2284 3594 -1252
rect 3654 -2344 3714 -1314
rect 3774 -1819 3834 -1252
rect 3894 -1819 3954 -1314
rect 3774 -1879 3954 -1819
rect 3774 -2284 3834 -1879
rect 3894 -2344 3954 -1879
rect 4014 -1406 4080 -1252
rect 4014 -1470 4015 -1406
rect 4079 -1470 4080 -1406
rect 4014 -1486 4080 -1470
rect 4014 -1550 4015 -1486
rect 4079 -1550 4080 -1486
rect 4014 -1566 4080 -1550
rect 4014 -1630 4015 -1566
rect 4079 -1630 4080 -1566
rect 4014 -1646 4080 -1630
rect 4014 -1710 4015 -1646
rect 4079 -1710 4080 -1646
rect 4014 -1726 4080 -1710
rect 4014 -1790 4015 -1726
rect 4079 -1790 4080 -1726
rect 4014 -1806 4080 -1790
rect 4014 -1870 4015 -1806
rect 4079 -1870 4080 -1806
rect 4014 -1886 4080 -1870
rect 4014 -1950 4015 -1886
rect 4079 -1950 4080 -1886
rect 4014 -1966 4080 -1950
rect 4014 -2030 4015 -1966
rect 4079 -2030 4080 -1966
rect 4014 -2046 4080 -2030
rect 4014 -2110 4015 -2046
rect 4079 -2110 4080 -2046
rect 4014 -2126 4080 -2110
rect 4014 -2190 4015 -2126
rect 4079 -2190 4080 -2126
rect 4014 -2280 4080 -2190
rect 4140 -1819 4200 -1314
rect 4260 -1819 4320 -1252
rect 4140 -1879 4320 -1819
rect 4140 -2344 4200 -1879
rect 4260 -2284 4320 -1879
rect 4380 -2344 4440 -1314
rect 4500 -2284 4560 -1252
rect 4620 -1406 4686 -1252
rect 4620 -1470 4621 -1406
rect 4685 -1470 4686 -1406
rect 4620 -1486 4686 -1470
rect 4620 -1550 4621 -1486
rect 4685 -1550 4686 -1486
rect 4620 -1566 4686 -1550
rect 4620 -1630 4621 -1566
rect 4685 -1630 4686 -1566
rect 4620 -1646 4686 -1630
rect 4620 -1710 4621 -1646
rect 4685 -1710 4686 -1646
rect 4620 -1726 4686 -1710
rect 4620 -1790 4621 -1726
rect 4685 -1790 4686 -1726
rect 4620 -1806 4686 -1790
rect 4620 -1870 4621 -1806
rect 4685 -1870 4686 -1806
rect 4620 -1886 4686 -1870
rect 4620 -1950 4621 -1886
rect 4685 -1950 4686 -1886
rect 4620 -1966 4686 -1950
rect 4620 -2030 4621 -1966
rect 4685 -2030 4686 -1966
rect 4620 -2046 4686 -2030
rect 4620 -2110 4621 -2046
rect 4685 -2110 4686 -2046
rect 4620 -2126 4686 -2110
rect 4620 -2190 4621 -2126
rect 4685 -2190 4686 -2126
rect 4620 -2280 4686 -2190
rect 4746 -2284 4806 -1252
rect 4866 -2344 4926 -1314
rect 4986 -1819 5046 -1252
rect 5106 -1819 5166 -1314
rect 4986 -1879 5166 -1819
rect 4986 -2284 5046 -1879
rect 5106 -2344 5166 -1879
rect 5226 -1406 5292 -1252
rect 5226 -1470 5227 -1406
rect 5291 -1470 5292 -1406
rect 5226 -1486 5292 -1470
rect 5226 -1550 5227 -1486
rect 5291 -1550 5292 -1486
rect 5226 -1566 5292 -1550
rect 5226 -1630 5227 -1566
rect 5291 -1630 5292 -1566
rect 5226 -1646 5292 -1630
rect 5226 -1710 5227 -1646
rect 5291 -1710 5292 -1646
rect 5226 -1726 5292 -1710
rect 5226 -1790 5227 -1726
rect 5291 -1790 5292 -1726
rect 5226 -1806 5292 -1790
rect 5226 -1870 5227 -1806
rect 5291 -1870 5292 -1806
rect 5226 -1886 5292 -1870
rect 5226 -1950 5227 -1886
rect 5291 -1950 5292 -1886
rect 5226 -1966 5292 -1950
rect 5226 -2030 5227 -1966
rect 5291 -2030 5292 -1966
rect 5226 -2046 5292 -2030
rect 5226 -2110 5227 -2046
rect 5291 -2110 5292 -2046
rect 5226 -2126 5292 -2110
rect 5226 -2190 5227 -2126
rect 5291 -2190 5292 -2126
rect 5226 -2280 5292 -2190
rect 5352 -1247 5456 -1183
rect 5520 -1247 5536 -1183
rect 5600 -1247 5616 -1183
rect 5680 -1247 5696 -1183
rect 5760 -1247 5776 -1183
rect 5840 -1247 5856 -1183
rect 5920 -1247 6024 -1183
rect 6245 -1202 6621 157
rect 6709 158 7272 217
rect 7336 158 7352 222
rect 7416 158 7432 222
rect 7496 158 7512 222
rect 7576 158 8006 222
rect 8070 158 8086 222
rect 8150 158 8166 222
rect 8230 158 8246 222
rect 8310 158 8612 222
rect 8676 158 8692 222
rect 8756 158 8772 222
rect 8836 158 8852 222
rect 8916 158 9344 222
rect 9408 158 9424 222
rect 9488 158 9504 222
rect 9568 158 9584 222
rect 9648 158 9950 222
rect 10014 158 10030 222
rect 10094 158 10110 222
rect 10174 158 10190 222
rect 10254 158 10556 222
rect 10620 158 10636 222
rect 10700 158 10716 222
rect 10780 158 10796 222
rect 10860 158 11162 222
rect 11226 158 11242 222
rect 11306 158 11322 222
rect 11386 158 11402 222
rect 11466 158 11894 222
rect 11958 158 11974 222
rect 12038 158 12054 222
rect 12118 158 12134 222
rect 12198 161 12676 222
rect 12740 161 13464 225
rect 12198 158 13464 161
rect 6709 157 13464 158
rect 6709 -700 7027 157
rect 7088 156 7760 157
rect 7822 156 9100 157
rect 9160 156 11650 157
rect 11710 156 12382 157
rect 6709 -764 6933 -700
rect 6997 -764 7027 -700
rect 6709 -774 7027 -764
rect 6709 -962 6907 -952
rect 6709 -1026 6842 -962
rect 6906 -1026 6907 -962
rect 6709 -1036 6907 -1026
rect 5352 -1249 6024 -1247
rect 5352 -1403 5418 -1249
rect 5352 -1467 5353 -1403
rect 5417 -1467 5418 -1403
rect 5352 -1483 5418 -1467
rect 5352 -1547 5353 -1483
rect 5417 -1547 5418 -1483
rect 5352 -1563 5418 -1547
rect 5352 -1627 5353 -1563
rect 5417 -1627 5418 -1563
rect 5352 -1643 5418 -1627
rect 5352 -1707 5353 -1643
rect 5417 -1707 5418 -1643
rect 5352 -1723 5418 -1707
rect 5352 -1787 5353 -1723
rect 5417 -1787 5418 -1723
rect 5352 -1803 5418 -1787
rect 5352 -1867 5353 -1803
rect 5417 -1867 5418 -1803
rect 5352 -1883 5418 -1867
rect 5352 -1947 5353 -1883
rect 5417 -1947 5418 -1883
rect 5352 -1963 5418 -1947
rect 5352 -2027 5353 -1963
rect 5417 -2027 5418 -1963
rect 5352 -2043 5418 -2027
rect 5352 -2107 5353 -2043
rect 5417 -2107 5418 -2043
rect 5352 -2123 5418 -2107
rect 5352 -2187 5353 -2123
rect 5417 -2187 5418 -2123
rect 5352 -2277 5418 -2187
rect 5478 -2281 5538 -1249
rect 5598 -2341 5658 -1311
rect 5718 -1816 5778 -1249
rect 5838 -1816 5898 -1311
rect 5718 -1876 5898 -1816
rect 5718 -2281 5778 -1876
rect 5838 -2341 5898 -1876
rect 5958 -1403 6024 -1249
rect 6246 -1266 6289 -1202
rect 6353 -1266 6432 -1202
rect 6496 -1266 6552 -1202
rect 6616 -1266 6623 -1202
rect 6246 -1281 6623 -1266
rect 5958 -1467 5959 -1403
rect 6023 -1467 6024 -1403
rect 5958 -1483 6024 -1467
rect 5958 -1547 5959 -1483
rect 6023 -1547 6024 -1483
rect 5958 -1563 6024 -1547
rect 5958 -1627 5959 -1563
rect 6023 -1627 6024 -1563
rect 5958 -1643 6024 -1627
rect 5958 -1707 5959 -1643
rect 6023 -1707 6024 -1643
rect 5958 -1723 6024 -1707
rect 5958 -1787 5959 -1723
rect 6023 -1787 6024 -1723
rect 6709 -1414 6769 -1036
rect 6967 -1155 7027 -774
rect 7088 2 7154 92
rect 7088 -62 7089 2
rect 7153 -62 7154 2
rect 7088 -78 7154 -62
rect 7088 -142 7089 -78
rect 7153 -142 7154 -78
rect 7088 -158 7154 -142
rect 7088 -222 7089 -158
rect 7153 -222 7154 -158
rect 7088 -238 7154 -222
rect 7088 -302 7089 -238
rect 7153 -302 7154 -238
rect 7088 -318 7154 -302
rect 7088 -382 7089 -318
rect 7153 -382 7154 -318
rect 7088 -398 7154 -382
rect 7088 -462 7089 -398
rect 7153 -462 7154 -398
rect 7088 -478 7154 -462
rect 7088 -542 7089 -478
rect 7153 -542 7154 -478
rect 7088 -558 7154 -542
rect 7088 -622 7089 -558
rect 7153 -622 7154 -558
rect 7088 -638 7154 -622
rect 7088 -702 7089 -638
rect 7153 -702 7154 -638
rect 7088 -718 7154 -702
rect 7088 -782 7089 -718
rect 7153 -782 7154 -718
rect 7088 -936 7154 -782
rect 7214 -166 7274 156
rect 7334 -166 7394 96
rect 7214 -242 7394 -166
rect 7214 -874 7274 -242
rect 7334 -936 7394 -242
rect 7454 -874 7514 156
rect 7574 -936 7634 96
rect 7694 2 7760 92
rect 7694 -62 7695 2
rect 7759 -62 7760 2
rect 7694 -78 7760 -62
rect 7694 -142 7695 -78
rect 7759 -142 7760 -78
rect 7694 -158 7760 -142
rect 7694 -222 7695 -158
rect 7759 -222 7760 -158
rect 7694 -238 7760 -222
rect 7694 -302 7695 -238
rect 7759 -302 7760 -238
rect 7694 -318 7760 -302
rect 7694 -382 7695 -318
rect 7759 -382 7760 -318
rect 7694 -398 7760 -382
rect 7694 -462 7695 -398
rect 7759 -462 7760 -398
rect 7694 -478 7760 -462
rect 7694 -542 7695 -478
rect 7759 -542 7760 -478
rect 7694 -558 7760 -542
rect 7694 -622 7695 -558
rect 7759 -622 7760 -558
rect 7694 -638 7760 -622
rect 7694 -702 7695 -638
rect 7759 -702 7760 -638
rect 7694 -718 7760 -702
rect 7694 -782 7695 -718
rect 7759 -782 7760 -718
rect 7694 -936 7760 -782
rect 7088 -938 7760 -936
rect 7088 -1002 7192 -938
rect 7256 -1002 7272 -938
rect 7336 -1002 7352 -938
rect 7416 -1002 7432 -938
rect 7496 -1002 7512 -938
rect 7576 -1002 7592 -938
rect 7656 -1002 7760 -938
rect 7088 -1004 7760 -1002
rect 7822 2 7888 92
rect 7822 -62 7823 2
rect 7887 -62 7888 2
rect 7822 -78 7888 -62
rect 7822 -142 7823 -78
rect 7887 -142 7888 -78
rect 7822 -158 7888 -142
rect 7822 -222 7823 -158
rect 7887 -222 7888 -158
rect 7822 -238 7888 -222
rect 7822 -302 7823 -238
rect 7887 -302 7888 -238
rect 7822 -318 7888 -302
rect 7822 -382 7823 -318
rect 7887 -382 7888 -318
rect 7822 -398 7888 -382
rect 7822 -462 7823 -398
rect 7887 -462 7888 -398
rect 7822 -478 7888 -462
rect 7822 -542 7823 -478
rect 7887 -542 7888 -478
rect 7822 -558 7888 -542
rect 7822 -622 7823 -558
rect 7887 -622 7888 -558
rect 7822 -638 7888 -622
rect 7822 -702 7823 -638
rect 7887 -702 7888 -638
rect 7822 -718 7888 -702
rect 7822 -782 7823 -718
rect 7887 -782 7888 -718
rect 7822 -936 7888 -782
rect 7948 -166 8008 156
rect 8068 -166 8128 96
rect 7948 -242 8128 -166
rect 7948 -874 8008 -242
rect 8068 -936 8128 -242
rect 8188 -874 8248 156
rect 8308 -936 8368 96
rect 8428 2 8494 92
rect 8428 -62 8429 2
rect 8493 -62 8494 2
rect 8428 -78 8494 -62
rect 8428 -142 8429 -78
rect 8493 -142 8494 -78
rect 8428 -158 8494 -142
rect 8428 -222 8429 -158
rect 8493 -222 8494 -158
rect 8428 -238 8494 -222
rect 8428 -302 8429 -238
rect 8493 -302 8494 -238
rect 8428 -318 8494 -302
rect 8428 -382 8429 -318
rect 8493 -382 8494 -318
rect 8428 -398 8494 -382
rect 8428 -462 8429 -398
rect 8493 -462 8494 -398
rect 8428 -478 8494 -462
rect 8428 -542 8429 -478
rect 8493 -542 8494 -478
rect 8428 -558 8494 -542
rect 8428 -622 8429 -558
rect 8493 -622 8494 -558
rect 8428 -638 8494 -622
rect 8428 -702 8429 -638
rect 8493 -702 8494 -638
rect 8428 -718 8494 -702
rect 8428 -782 8429 -718
rect 8493 -782 8494 -718
rect 8428 -936 8494 -782
rect 8554 -936 8614 96
rect 8674 -874 8734 156
rect 8794 -166 8854 96
rect 8914 -166 8974 156
rect 8794 -242 8974 -166
rect 8794 -936 8854 -242
rect 8914 -874 8974 -242
rect 9034 2 9100 92
rect 9034 -62 9035 2
rect 9099 -62 9100 2
rect 9034 -78 9100 -62
rect 9034 -142 9035 -78
rect 9099 -142 9100 -78
rect 9034 -158 9100 -142
rect 9034 -222 9035 -158
rect 9099 -222 9100 -158
rect 9034 -238 9100 -222
rect 9034 -302 9035 -238
rect 9099 -302 9100 -238
rect 9034 -318 9100 -302
rect 9034 -382 9035 -318
rect 9099 -382 9100 -318
rect 9034 -398 9100 -382
rect 9034 -462 9035 -398
rect 9099 -462 9100 -398
rect 9034 -478 9100 -462
rect 9034 -542 9035 -478
rect 9099 -542 9100 -478
rect 9034 -558 9100 -542
rect 9034 -622 9035 -558
rect 9099 -622 9100 -558
rect 9034 -638 9100 -622
rect 9034 -702 9035 -638
rect 9099 -702 9100 -638
rect 9034 -718 9100 -702
rect 9034 -782 9035 -718
rect 9099 -782 9100 -718
rect 9034 -936 9100 -782
rect 7822 -938 9100 -936
rect 7822 -1002 7926 -938
rect 7990 -1002 8006 -938
rect 8070 -1002 8086 -938
rect 8150 -1002 8166 -938
rect 8230 -1002 8246 -938
rect 8310 -1002 8326 -938
rect 8390 -1002 8532 -938
rect 8596 -1002 8612 -938
rect 8676 -1002 8692 -938
rect 8756 -1002 8772 -938
rect 8836 -1002 8852 -938
rect 8916 -1002 8932 -938
rect 8996 -1002 9100 -938
rect 7822 -1004 9100 -1002
rect 9160 2 9226 92
rect 9160 -62 9161 2
rect 9225 -62 9226 2
rect 9160 -78 9226 -62
rect 9160 -142 9161 -78
rect 9225 -142 9226 -78
rect 9160 -158 9226 -142
rect 9160 -222 9161 -158
rect 9225 -222 9226 -158
rect 9160 -238 9226 -222
rect 9160 -302 9161 -238
rect 9225 -302 9226 -238
rect 9160 -318 9226 -302
rect 9160 -382 9161 -318
rect 9225 -382 9226 -318
rect 9160 -398 9226 -382
rect 9160 -462 9161 -398
rect 9225 -462 9226 -398
rect 9160 -478 9226 -462
rect 9160 -542 9161 -478
rect 9225 -542 9226 -478
rect 9160 -558 9226 -542
rect 9160 -622 9161 -558
rect 9225 -622 9226 -558
rect 9160 -638 9226 -622
rect 9160 -702 9161 -638
rect 9225 -702 9226 -638
rect 9160 -718 9226 -702
rect 9160 -782 9161 -718
rect 9225 -782 9226 -718
rect 9160 -936 9226 -782
rect 9286 -166 9346 156
rect 9406 -166 9466 96
rect 9286 -242 9466 -166
rect 9286 -874 9346 -242
rect 9406 -936 9466 -242
rect 9526 -874 9586 156
rect 9646 -936 9706 96
rect 9766 2 9832 92
rect 9766 -62 9767 2
rect 9831 -62 9832 2
rect 9766 -78 9832 -62
rect 9766 -142 9767 -78
rect 9831 -142 9832 -78
rect 9766 -158 9832 -142
rect 9766 -222 9767 -158
rect 9831 -222 9832 -158
rect 9766 -238 9832 -222
rect 9766 -302 9767 -238
rect 9831 -302 9832 -238
rect 9766 -318 9832 -302
rect 9766 -382 9767 -318
rect 9831 -382 9832 -318
rect 9766 -398 9832 -382
rect 9766 -462 9767 -398
rect 9831 -462 9832 -398
rect 9766 -478 9832 -462
rect 9766 -542 9767 -478
rect 9831 -542 9832 -478
rect 9766 -558 9832 -542
rect 9766 -622 9767 -558
rect 9831 -622 9832 -558
rect 9766 -638 9832 -622
rect 9766 -702 9767 -638
rect 9831 -702 9832 -638
rect 9766 -718 9832 -702
rect 9766 -782 9767 -718
rect 9831 -782 9832 -718
rect 9766 -936 9832 -782
rect 9892 -936 9952 96
rect 10012 -874 10072 156
rect 10132 -166 10192 96
rect 10252 -166 10312 156
rect 10132 -242 10312 -166
rect 10132 -936 10192 -242
rect 10252 -874 10312 -242
rect 10372 2 10438 92
rect 10372 -62 10373 2
rect 10437 -62 10438 2
rect 10372 -78 10438 -62
rect 10372 -142 10373 -78
rect 10437 -142 10438 -78
rect 10372 -158 10438 -142
rect 10372 -222 10373 -158
rect 10437 -222 10438 -158
rect 10372 -238 10438 -222
rect 10372 -302 10373 -238
rect 10437 -302 10438 -238
rect 10372 -318 10438 -302
rect 10372 -382 10373 -318
rect 10437 -382 10438 -318
rect 10372 -398 10438 -382
rect 10372 -462 10373 -398
rect 10437 -462 10438 -398
rect 10372 -478 10438 -462
rect 10372 -542 10373 -478
rect 10437 -542 10438 -478
rect 10372 -558 10438 -542
rect 10372 -622 10373 -558
rect 10437 -622 10438 -558
rect 10372 -638 10438 -622
rect 10372 -702 10373 -638
rect 10437 -702 10438 -638
rect 10372 -718 10438 -702
rect 10372 -782 10373 -718
rect 10437 -782 10438 -718
rect 10372 -936 10438 -782
rect 10498 -166 10558 156
rect 10618 -166 10678 96
rect 10498 -242 10678 -166
rect 10498 -874 10558 -242
rect 10618 -936 10678 -242
rect 10738 -874 10798 156
rect 10858 -936 10918 96
rect 10978 2 11044 92
rect 10978 -62 10979 2
rect 11043 -62 11044 2
rect 10978 -78 11044 -62
rect 10978 -142 10979 -78
rect 11043 -142 11044 -78
rect 10978 -158 11044 -142
rect 10978 -222 10979 -158
rect 11043 -222 11044 -158
rect 10978 -238 11044 -222
rect 10978 -302 10979 -238
rect 11043 -302 11044 -238
rect 10978 -318 11044 -302
rect 10978 -382 10979 -318
rect 11043 -382 11044 -318
rect 10978 -398 11044 -382
rect 10978 -462 10979 -398
rect 11043 -462 11044 -398
rect 10978 -478 11044 -462
rect 10978 -542 10979 -478
rect 11043 -542 11044 -478
rect 10978 -558 11044 -542
rect 10978 -622 10979 -558
rect 11043 -622 11044 -558
rect 10978 -638 11044 -622
rect 10978 -702 10979 -638
rect 11043 -702 11044 -638
rect 10978 -718 11044 -702
rect 10978 -782 10979 -718
rect 11043 -782 11044 -718
rect 10978 -936 11044 -782
rect 11104 -936 11164 96
rect 11224 -874 11284 156
rect 11344 -166 11404 96
rect 11464 -166 11524 156
rect 11344 -242 11524 -166
rect 11344 -936 11404 -242
rect 11464 -874 11524 -242
rect 11584 2 11650 92
rect 11584 -62 11585 2
rect 11649 -62 11650 2
rect 11584 -78 11650 -62
rect 11584 -142 11585 -78
rect 11649 -142 11650 -78
rect 11584 -158 11650 -142
rect 11584 -222 11585 -158
rect 11649 -222 11650 -158
rect 11584 -238 11650 -222
rect 11584 -302 11585 -238
rect 11649 -302 11650 -238
rect 11584 -318 11650 -302
rect 11584 -382 11585 -318
rect 11649 -382 11650 -318
rect 11584 -398 11650 -382
rect 11584 -462 11585 -398
rect 11649 -462 11650 -398
rect 11584 -478 11650 -462
rect 11584 -542 11585 -478
rect 11649 -542 11650 -478
rect 11584 -558 11650 -542
rect 11584 -622 11585 -558
rect 11649 -622 11650 -558
rect 11584 -638 11650 -622
rect 11584 -702 11585 -638
rect 11649 -702 11650 -638
rect 11584 -718 11650 -702
rect 11584 -782 11585 -718
rect 11649 -782 11650 -718
rect 11584 -936 11650 -782
rect 9160 -938 11650 -936
rect 9160 -1002 9264 -938
rect 9328 -1002 9344 -938
rect 9408 -1002 9424 -938
rect 9488 -1002 9504 -938
rect 9568 -1002 9584 -938
rect 9648 -1002 9664 -938
rect 9728 -1002 9870 -938
rect 9934 -1002 9950 -938
rect 10014 -1002 10030 -938
rect 10094 -1002 10110 -938
rect 10174 -1002 10190 -938
rect 10254 -1002 10270 -938
rect 10334 -1002 10476 -938
rect 10540 -1002 10556 -938
rect 10620 -1002 10636 -938
rect 10700 -1002 10716 -938
rect 10780 -1002 10796 -938
rect 10860 -1002 10876 -938
rect 10940 -1002 11082 -938
rect 11146 -1002 11162 -938
rect 11226 -1002 11242 -938
rect 11306 -1002 11322 -938
rect 11386 -1002 11402 -938
rect 11466 -1002 11482 -938
rect 11546 -1002 11650 -938
rect 9160 -1004 11650 -1002
rect 11710 2 11776 92
rect 11710 -62 11711 2
rect 11775 -62 11776 2
rect 11710 -78 11776 -62
rect 11710 -142 11711 -78
rect 11775 -142 11776 -78
rect 11710 -158 11776 -142
rect 11710 -222 11711 -158
rect 11775 -222 11776 -158
rect 11710 -238 11776 -222
rect 11710 -302 11711 -238
rect 11775 -302 11776 -238
rect 11710 -318 11776 -302
rect 11710 -382 11711 -318
rect 11775 -382 11776 -318
rect 11710 -398 11776 -382
rect 11710 -462 11711 -398
rect 11775 -462 11776 -398
rect 11710 -478 11776 -462
rect 11710 -542 11711 -478
rect 11775 -542 11776 -478
rect 11710 -558 11776 -542
rect 11710 -622 11711 -558
rect 11775 -622 11776 -558
rect 11710 -638 11776 -622
rect 11710 -702 11711 -638
rect 11775 -702 11776 -638
rect 11710 -718 11776 -702
rect 11710 -782 11711 -718
rect 11775 -782 11776 -718
rect 11710 -936 11776 -782
rect 11836 -936 11896 96
rect 11956 -874 12016 156
rect 12076 -166 12136 96
rect 12196 -166 12256 156
rect 12645 151 12770 157
rect 12076 -242 12256 -166
rect 12076 -936 12136 -242
rect 12196 -874 12256 -242
rect 12316 2 12382 92
rect 12316 -62 12317 2
rect 12381 -62 12382 2
rect 12316 -78 12382 -62
rect 12316 -142 12317 -78
rect 12381 -142 12382 -78
rect 12316 -158 12382 -142
rect 12316 -222 12317 -158
rect 12381 -222 12382 -158
rect 12316 -238 12382 -222
rect 12316 -302 12317 -238
rect 12381 -302 12382 -238
rect 12316 -318 12382 -302
rect 12316 -382 12317 -318
rect 12381 -382 12382 -318
rect 12316 -398 12382 -382
rect 12316 -462 12317 -398
rect 12381 -462 12382 -398
rect 12316 -478 12382 -462
rect 12316 -542 12317 -478
rect 12381 -542 12382 -478
rect 12316 -558 12382 -542
rect 12316 -622 12317 -558
rect 12381 -622 12382 -558
rect 12316 -638 12382 -622
rect 12316 -702 12317 -638
rect 12381 -702 12382 -638
rect 12316 -718 12382 -702
rect 12316 -782 12317 -718
rect 12381 -782 12382 -718
rect 12316 -936 12382 -782
rect 11710 -938 12382 -936
rect 11710 -1002 11814 -938
rect 11878 -1002 11894 -938
rect 11958 -1002 11974 -938
rect 12038 -1002 12054 -938
rect 12118 -1002 12134 -938
rect 12198 -1002 12214 -938
rect 12278 -1002 12382 -938
rect 11710 -1004 12382 -1002
rect 6829 -1165 7027 -1155
rect 6829 -1229 6842 -1165
rect 6906 -1229 7027 -1165
rect 12061 -1183 12733 -1181
rect 6829 -1239 7027 -1229
rect 7087 -1186 12001 -1184
rect 7087 -1250 7191 -1186
rect 7255 -1250 7271 -1186
rect 7335 -1250 7351 -1186
rect 7415 -1250 7431 -1186
rect 7495 -1250 7511 -1186
rect 7575 -1250 7591 -1186
rect 7655 -1250 7797 -1186
rect 7861 -1250 7877 -1186
rect 7941 -1250 7957 -1186
rect 8021 -1250 8037 -1186
rect 8101 -1250 8117 -1186
rect 8181 -1250 8197 -1186
rect 8261 -1250 8403 -1186
rect 8467 -1250 8483 -1186
rect 8547 -1250 8563 -1186
rect 8627 -1250 8643 -1186
rect 8707 -1250 8723 -1186
rect 8787 -1250 8803 -1186
rect 8867 -1250 9009 -1186
rect 9073 -1250 9089 -1186
rect 9153 -1250 9169 -1186
rect 9233 -1250 9249 -1186
rect 9313 -1250 9329 -1186
rect 9393 -1250 9409 -1186
rect 9473 -1250 9615 -1186
rect 9679 -1250 9695 -1186
rect 9759 -1250 9775 -1186
rect 9839 -1250 9855 -1186
rect 9919 -1250 9935 -1186
rect 9999 -1250 10015 -1186
rect 10079 -1250 10221 -1186
rect 10285 -1250 10301 -1186
rect 10365 -1250 10381 -1186
rect 10445 -1250 10461 -1186
rect 10525 -1250 10541 -1186
rect 10605 -1250 10621 -1186
rect 10685 -1250 10827 -1186
rect 10891 -1250 10907 -1186
rect 10971 -1250 10987 -1186
rect 11051 -1250 11067 -1186
rect 11131 -1250 11147 -1186
rect 11211 -1250 11227 -1186
rect 11291 -1250 11433 -1186
rect 11497 -1250 11513 -1186
rect 11577 -1250 11593 -1186
rect 11657 -1250 11673 -1186
rect 11737 -1250 11753 -1186
rect 11817 -1250 11833 -1186
rect 11897 -1250 12001 -1186
rect 7087 -1252 12001 -1250
rect 7087 -1406 7153 -1252
rect 6709 -1426 7027 -1414
rect 6709 -1490 6930 -1426
rect 6994 -1490 7027 -1426
rect 6709 -1668 7027 -1490
rect 5958 -1803 6024 -1787
rect 5958 -1867 5959 -1803
rect 6023 -1867 6024 -1803
rect 6232 -1747 6649 -1729
rect 6232 -1748 6439 -1747
rect 6232 -1806 6295 -1748
rect 5958 -1883 6024 -1867
rect 5958 -1947 5959 -1883
rect 6023 -1947 6024 -1883
rect 5958 -1963 6024 -1947
rect 5958 -2027 5959 -1963
rect 6023 -2027 6024 -1963
rect 5958 -2043 6024 -2027
rect 5958 -2107 5959 -2043
rect 6023 -2107 6024 -2043
rect 5958 -2123 6024 -2107
rect 5958 -2187 5959 -2123
rect 6023 -2187 6024 -2123
rect 5958 -2277 6024 -2187
rect 6231 -1812 6295 -1806
rect 6359 -1811 6439 -1748
rect 6503 -1748 6649 -1747
rect 6503 -1811 6570 -1748
rect 6359 -1812 6570 -1811
rect 6634 -1812 6649 -1748
rect 6231 -1897 6649 -1812
rect 6231 -1961 6425 -1897
rect 6489 -1961 6649 -1897
rect 6231 -2093 6649 -1961
rect 6231 -2157 6425 -2093
rect 6489 -2157 6649 -2093
rect 6231 -2268 6649 -2157
rect 6231 -2332 6425 -2268
rect 6489 -2332 6649 -2268
rect 5352 -2342 6024 -2341
rect 5351 -2343 6024 -2342
rect 5351 -2344 5456 -2343
rect 208 -2346 5456 -2344
rect 208 -2355 482 -2346
rect 0 -2392 482 -2355
rect -2 -2410 482 -2392
rect 546 -2410 562 -2346
rect 626 -2410 642 -2346
rect 706 -2410 722 -2346
rect 786 -2410 802 -2346
rect 866 -2410 882 -2346
rect 946 -2410 1088 -2346
rect 1152 -2410 1168 -2346
rect 1232 -2410 1248 -2346
rect 1312 -2410 1328 -2346
rect 1392 -2410 1408 -2346
rect 1472 -2410 1488 -2346
rect 1552 -2410 1694 -2346
rect 1758 -2410 1774 -2346
rect 1838 -2410 1854 -2346
rect 1918 -2410 1934 -2346
rect 1998 -2410 2014 -2346
rect 2078 -2410 2094 -2346
rect 2158 -2410 2300 -2346
rect 2364 -2410 2380 -2346
rect 2444 -2410 2460 -2346
rect 2524 -2410 2540 -2346
rect 2604 -2410 2620 -2346
rect 2684 -2410 2700 -2346
rect 2764 -2410 2906 -2346
rect 2970 -2410 2986 -2346
rect 3050 -2410 3066 -2346
rect 3130 -2410 3146 -2346
rect 3210 -2410 3226 -2346
rect 3290 -2410 3306 -2346
rect 3370 -2410 3512 -2346
rect 3576 -2410 3592 -2346
rect 3656 -2410 3672 -2346
rect 3736 -2410 3752 -2346
rect 3816 -2410 3832 -2346
rect 3896 -2410 3912 -2346
rect 3976 -2410 4118 -2346
rect 4182 -2410 4198 -2346
rect 4262 -2410 4278 -2346
rect 4342 -2410 4358 -2346
rect 4422 -2410 4438 -2346
rect 4502 -2410 4518 -2346
rect 4582 -2410 4724 -2346
rect 4788 -2410 4804 -2346
rect 4868 -2410 4884 -2346
rect 4948 -2410 4964 -2346
rect 5028 -2410 5044 -2346
rect 5108 -2410 5124 -2346
rect 5188 -2407 5456 -2346
rect 5520 -2407 5536 -2343
rect 5600 -2407 5616 -2343
rect 5680 -2407 5696 -2343
rect 5760 -2407 5776 -2343
rect 5840 -2407 5856 -2343
rect 5920 -2344 6024 -2343
rect 6231 -2344 6649 -2332
rect 5920 -2353 6649 -2344
rect 5920 -2407 5953 -2353
rect 5188 -2410 5953 -2407
rect -2 -2417 5953 -2410
rect 6017 -2392 6649 -2353
rect 6709 -1732 6848 -1668
rect 6912 -1732 7027 -1668
rect 6709 -1825 7027 -1732
rect 6709 -1889 6847 -1825
rect 6911 -1889 7027 -1825
rect 6709 -1995 7027 -1889
rect 6709 -2059 6847 -1995
rect 6911 -2059 7027 -1995
rect 6709 -2147 7027 -2059
rect 6709 -2211 6848 -2147
rect 6912 -2211 7027 -2147
rect 6709 -2291 7027 -2211
rect 7087 -1470 7088 -1406
rect 7152 -1470 7153 -1406
rect 7087 -1486 7153 -1470
rect 7087 -1550 7088 -1486
rect 7152 -1550 7153 -1486
rect 7087 -1566 7153 -1550
rect 7087 -1630 7088 -1566
rect 7152 -1630 7153 -1566
rect 7087 -1646 7153 -1630
rect 7087 -1710 7088 -1646
rect 7152 -1710 7153 -1646
rect 7087 -1726 7153 -1710
rect 7087 -1790 7088 -1726
rect 7152 -1790 7153 -1726
rect 7087 -1806 7153 -1790
rect 7087 -1870 7088 -1806
rect 7152 -1870 7153 -1806
rect 7087 -1886 7153 -1870
rect 7087 -1950 7088 -1886
rect 7152 -1950 7153 -1886
rect 7087 -1966 7153 -1950
rect 7087 -2030 7088 -1966
rect 7152 -2030 7153 -1966
rect 7087 -2046 7153 -2030
rect 7087 -2110 7088 -2046
rect 7152 -2110 7153 -2046
rect 7087 -2126 7153 -2110
rect 7087 -2190 7088 -2126
rect 7152 -2190 7153 -2126
rect 7087 -2280 7153 -2190
rect 7213 -1819 7273 -1314
rect 7333 -1819 7393 -1252
rect 7213 -1879 7393 -1819
rect 6709 -2355 6853 -2291
rect 6917 -2344 7027 -2291
rect 7213 -2344 7273 -1879
rect 7333 -2284 7393 -1879
rect 7453 -2344 7513 -1314
rect 7573 -2284 7633 -1252
rect 7693 -1406 7759 -1252
rect 7693 -1470 7694 -1406
rect 7758 -1470 7759 -1406
rect 7693 -1486 7759 -1470
rect 7693 -1550 7694 -1486
rect 7758 -1550 7759 -1486
rect 7693 -1566 7759 -1550
rect 7693 -1630 7694 -1566
rect 7758 -1630 7759 -1566
rect 7693 -1646 7759 -1630
rect 7693 -1710 7694 -1646
rect 7758 -1710 7759 -1646
rect 7693 -1726 7759 -1710
rect 7693 -1790 7694 -1726
rect 7758 -1790 7759 -1726
rect 7693 -1806 7759 -1790
rect 7693 -1870 7694 -1806
rect 7758 -1870 7759 -1806
rect 7693 -1886 7759 -1870
rect 7693 -1950 7694 -1886
rect 7758 -1950 7759 -1886
rect 7693 -1966 7759 -1950
rect 7693 -2030 7694 -1966
rect 7758 -2030 7759 -1966
rect 7693 -2046 7759 -2030
rect 7693 -2110 7694 -2046
rect 7758 -2110 7759 -2046
rect 7693 -2126 7759 -2110
rect 7693 -2190 7694 -2126
rect 7758 -2190 7759 -2126
rect 7693 -2280 7759 -2190
rect 7819 -2284 7879 -1252
rect 7939 -2344 7999 -1314
rect 8059 -1819 8119 -1252
rect 8179 -1819 8239 -1314
rect 8059 -1879 8239 -1819
rect 8059 -2284 8119 -1879
rect 8179 -2344 8239 -1879
rect 8299 -1406 8365 -1252
rect 8299 -1470 8300 -1406
rect 8364 -1470 8365 -1406
rect 8299 -1486 8365 -1470
rect 8299 -1550 8300 -1486
rect 8364 -1550 8365 -1486
rect 8299 -1566 8365 -1550
rect 8299 -1630 8300 -1566
rect 8364 -1630 8365 -1566
rect 8299 -1646 8365 -1630
rect 8299 -1710 8300 -1646
rect 8364 -1710 8365 -1646
rect 8299 -1726 8365 -1710
rect 8299 -1790 8300 -1726
rect 8364 -1790 8365 -1726
rect 8299 -1806 8365 -1790
rect 8299 -1870 8300 -1806
rect 8364 -1870 8365 -1806
rect 8299 -1886 8365 -1870
rect 8299 -1950 8300 -1886
rect 8364 -1950 8365 -1886
rect 8299 -1966 8365 -1950
rect 8299 -2030 8300 -1966
rect 8364 -2030 8365 -1966
rect 8299 -2046 8365 -2030
rect 8299 -2110 8300 -2046
rect 8364 -2110 8365 -2046
rect 8299 -2126 8365 -2110
rect 8299 -2190 8300 -2126
rect 8364 -2190 8365 -2126
rect 8299 -2280 8365 -2190
rect 8425 -1819 8485 -1314
rect 8545 -1819 8605 -1252
rect 8425 -1879 8605 -1819
rect 8425 -2344 8485 -1879
rect 8545 -2284 8605 -1879
rect 8665 -2344 8725 -1314
rect 8785 -2284 8845 -1252
rect 8905 -1406 8971 -1252
rect 8905 -1470 8906 -1406
rect 8970 -1470 8971 -1406
rect 8905 -1486 8971 -1470
rect 8905 -1550 8906 -1486
rect 8970 -1550 8971 -1486
rect 8905 -1566 8971 -1550
rect 8905 -1630 8906 -1566
rect 8970 -1630 8971 -1566
rect 8905 -1646 8971 -1630
rect 8905 -1710 8906 -1646
rect 8970 -1710 8971 -1646
rect 8905 -1726 8971 -1710
rect 8905 -1790 8906 -1726
rect 8970 -1790 8971 -1726
rect 8905 -1806 8971 -1790
rect 8905 -1870 8906 -1806
rect 8970 -1870 8971 -1806
rect 8905 -1886 8971 -1870
rect 8905 -1950 8906 -1886
rect 8970 -1950 8971 -1886
rect 8905 -1966 8971 -1950
rect 8905 -2030 8906 -1966
rect 8970 -2030 8971 -1966
rect 8905 -2046 8971 -2030
rect 8905 -2110 8906 -2046
rect 8970 -2110 8971 -2046
rect 8905 -2126 8971 -2110
rect 8905 -2190 8906 -2126
rect 8970 -2190 8971 -2126
rect 8905 -2280 8971 -2190
rect 9031 -2284 9091 -1252
rect 9151 -2344 9211 -1314
rect 9271 -1819 9331 -1252
rect 9391 -1819 9451 -1314
rect 9271 -1879 9451 -1819
rect 9271 -2284 9331 -1879
rect 9391 -2344 9451 -1879
rect 9511 -1406 9577 -1252
rect 9511 -1470 9512 -1406
rect 9576 -1470 9577 -1406
rect 9511 -1486 9577 -1470
rect 9511 -1550 9512 -1486
rect 9576 -1550 9577 -1486
rect 9511 -1566 9577 -1550
rect 9511 -1630 9512 -1566
rect 9576 -1630 9577 -1566
rect 9511 -1646 9577 -1630
rect 9511 -1710 9512 -1646
rect 9576 -1710 9577 -1646
rect 9511 -1726 9577 -1710
rect 9511 -1790 9512 -1726
rect 9576 -1790 9577 -1726
rect 9511 -1806 9577 -1790
rect 9511 -1870 9512 -1806
rect 9576 -1870 9577 -1806
rect 9511 -1886 9577 -1870
rect 9511 -1950 9512 -1886
rect 9576 -1950 9577 -1886
rect 9511 -1966 9577 -1950
rect 9511 -2030 9512 -1966
rect 9576 -2030 9577 -1966
rect 9511 -2046 9577 -2030
rect 9511 -2110 9512 -2046
rect 9576 -2110 9577 -2046
rect 9511 -2126 9577 -2110
rect 9511 -2190 9512 -2126
rect 9576 -2190 9577 -2126
rect 9511 -2280 9577 -2190
rect 9637 -1819 9697 -1314
rect 9757 -1819 9817 -1252
rect 9637 -1879 9817 -1819
rect 9637 -2344 9697 -1879
rect 9757 -2284 9817 -1879
rect 9877 -2344 9937 -1314
rect 9997 -2284 10057 -1252
rect 10117 -1406 10183 -1252
rect 10117 -1470 10118 -1406
rect 10182 -1470 10183 -1406
rect 10117 -1486 10183 -1470
rect 10117 -1550 10118 -1486
rect 10182 -1550 10183 -1486
rect 10117 -1566 10183 -1550
rect 10117 -1630 10118 -1566
rect 10182 -1630 10183 -1566
rect 10117 -1646 10183 -1630
rect 10117 -1710 10118 -1646
rect 10182 -1710 10183 -1646
rect 10117 -1726 10183 -1710
rect 10117 -1790 10118 -1726
rect 10182 -1790 10183 -1726
rect 10117 -1806 10183 -1790
rect 10117 -1870 10118 -1806
rect 10182 -1870 10183 -1806
rect 10117 -1886 10183 -1870
rect 10117 -1950 10118 -1886
rect 10182 -1950 10183 -1886
rect 10117 -1966 10183 -1950
rect 10117 -2030 10118 -1966
rect 10182 -2030 10183 -1966
rect 10117 -2046 10183 -2030
rect 10117 -2110 10118 -2046
rect 10182 -2110 10183 -2046
rect 10117 -2126 10183 -2110
rect 10117 -2190 10118 -2126
rect 10182 -2190 10183 -2126
rect 10117 -2280 10183 -2190
rect 10243 -2284 10303 -1252
rect 10363 -2344 10423 -1314
rect 10483 -1819 10543 -1252
rect 10603 -1819 10663 -1314
rect 10483 -1879 10663 -1819
rect 10483 -2284 10543 -1879
rect 10603 -2344 10663 -1879
rect 10723 -1406 10789 -1252
rect 10723 -1470 10724 -1406
rect 10788 -1470 10789 -1406
rect 10723 -1486 10789 -1470
rect 10723 -1550 10724 -1486
rect 10788 -1550 10789 -1486
rect 10723 -1566 10789 -1550
rect 10723 -1630 10724 -1566
rect 10788 -1630 10789 -1566
rect 10723 -1646 10789 -1630
rect 10723 -1710 10724 -1646
rect 10788 -1710 10789 -1646
rect 10723 -1726 10789 -1710
rect 10723 -1790 10724 -1726
rect 10788 -1790 10789 -1726
rect 10723 -1806 10789 -1790
rect 10723 -1870 10724 -1806
rect 10788 -1870 10789 -1806
rect 10723 -1886 10789 -1870
rect 10723 -1950 10724 -1886
rect 10788 -1950 10789 -1886
rect 10723 -1966 10789 -1950
rect 10723 -2030 10724 -1966
rect 10788 -2030 10789 -1966
rect 10723 -2046 10789 -2030
rect 10723 -2110 10724 -2046
rect 10788 -2110 10789 -2046
rect 10723 -2126 10789 -2110
rect 10723 -2190 10724 -2126
rect 10788 -2190 10789 -2126
rect 10723 -2280 10789 -2190
rect 10849 -1819 10909 -1314
rect 10969 -1819 11029 -1252
rect 10849 -1879 11029 -1819
rect 10849 -2344 10909 -1879
rect 10969 -2284 11029 -1879
rect 11089 -2344 11149 -1314
rect 11209 -2284 11269 -1252
rect 11329 -1406 11395 -1252
rect 11329 -1470 11330 -1406
rect 11394 -1470 11395 -1406
rect 11329 -1486 11395 -1470
rect 11329 -1550 11330 -1486
rect 11394 -1550 11395 -1486
rect 11329 -1566 11395 -1550
rect 11329 -1630 11330 -1566
rect 11394 -1630 11395 -1566
rect 11329 -1646 11395 -1630
rect 11329 -1710 11330 -1646
rect 11394 -1710 11395 -1646
rect 11329 -1726 11395 -1710
rect 11329 -1790 11330 -1726
rect 11394 -1790 11395 -1726
rect 11329 -1806 11395 -1790
rect 11329 -1870 11330 -1806
rect 11394 -1870 11395 -1806
rect 11329 -1886 11395 -1870
rect 11329 -1950 11330 -1886
rect 11394 -1950 11395 -1886
rect 11329 -1966 11395 -1950
rect 11329 -2030 11330 -1966
rect 11394 -2030 11395 -1966
rect 11329 -2046 11395 -2030
rect 11329 -2110 11330 -2046
rect 11394 -2110 11395 -2046
rect 11329 -2126 11395 -2110
rect 11329 -2190 11330 -2126
rect 11394 -2190 11395 -2126
rect 11329 -2280 11395 -2190
rect 11455 -2284 11515 -1252
rect 11575 -2344 11635 -1314
rect 11695 -1819 11755 -1252
rect 11815 -1819 11875 -1314
rect 11695 -1879 11875 -1819
rect 11695 -2284 11755 -1879
rect 11815 -2344 11875 -1879
rect 11935 -1406 12001 -1252
rect 11935 -1470 11936 -1406
rect 12000 -1470 12001 -1406
rect 11935 -1486 12001 -1470
rect 11935 -1550 11936 -1486
rect 12000 -1550 12001 -1486
rect 11935 -1566 12001 -1550
rect 11935 -1630 11936 -1566
rect 12000 -1630 12001 -1566
rect 11935 -1646 12001 -1630
rect 11935 -1710 11936 -1646
rect 12000 -1710 12001 -1646
rect 11935 -1726 12001 -1710
rect 11935 -1790 11936 -1726
rect 12000 -1790 12001 -1726
rect 11935 -1806 12001 -1790
rect 11935 -1870 11936 -1806
rect 12000 -1870 12001 -1806
rect 11935 -1886 12001 -1870
rect 11935 -1950 11936 -1886
rect 12000 -1950 12001 -1886
rect 11935 -1966 12001 -1950
rect 11935 -2030 11936 -1966
rect 12000 -2030 12001 -1966
rect 11935 -2046 12001 -2030
rect 11935 -2110 11936 -2046
rect 12000 -2110 12001 -2046
rect 11935 -2126 12001 -2110
rect 11935 -2190 11936 -2126
rect 12000 -2190 12001 -2126
rect 11935 -2280 12001 -2190
rect 12061 -1247 12165 -1183
rect 12229 -1247 12245 -1183
rect 12309 -1247 12325 -1183
rect 12389 -1247 12405 -1183
rect 12469 -1247 12485 -1183
rect 12549 -1247 12565 -1183
rect 12629 -1247 12733 -1183
rect 12954 -1202 13464 157
rect 12061 -1249 12733 -1247
rect 12061 -1403 12127 -1249
rect 12061 -1467 12062 -1403
rect 12126 -1467 12127 -1403
rect 12061 -1483 12127 -1467
rect 12061 -1547 12062 -1483
rect 12126 -1547 12127 -1483
rect 12061 -1563 12127 -1547
rect 12061 -1627 12062 -1563
rect 12126 -1627 12127 -1563
rect 12061 -1643 12127 -1627
rect 12061 -1707 12062 -1643
rect 12126 -1707 12127 -1643
rect 12061 -1723 12127 -1707
rect 12061 -1787 12062 -1723
rect 12126 -1787 12127 -1723
rect 12061 -1803 12127 -1787
rect 12061 -1867 12062 -1803
rect 12126 -1867 12127 -1803
rect 12061 -1883 12127 -1867
rect 12061 -1947 12062 -1883
rect 12126 -1947 12127 -1883
rect 12061 -1963 12127 -1947
rect 12061 -2027 12062 -1963
rect 12126 -2027 12127 -1963
rect 12061 -2043 12127 -2027
rect 12061 -2107 12062 -2043
rect 12126 -2107 12127 -2043
rect 12061 -2123 12127 -2107
rect 12061 -2187 12062 -2123
rect 12126 -2187 12127 -2123
rect 12061 -2277 12127 -2187
rect 12187 -2281 12247 -1249
rect 12307 -2341 12367 -1311
rect 12427 -1816 12487 -1249
rect 12547 -1816 12607 -1311
rect 12427 -1876 12607 -1816
rect 12427 -2281 12487 -1876
rect 12547 -2341 12607 -1876
rect 12667 -1403 12733 -1249
rect 12955 -1266 12998 -1202
rect 13062 -1266 13141 -1202
rect 13205 -1266 13261 -1202
rect 13325 -1205 13464 -1202
rect 13325 -1266 13332 -1205
rect 12955 -1281 13332 -1266
rect 12667 -1467 12668 -1403
rect 12732 -1467 12733 -1403
rect 12667 -1483 12733 -1467
rect 12667 -1547 12668 -1483
rect 12732 -1547 12733 -1483
rect 12667 -1563 12733 -1547
rect 12667 -1627 12668 -1563
rect 12732 -1627 12733 -1563
rect 12667 -1643 12733 -1627
rect 12667 -1707 12668 -1643
rect 12732 -1707 12733 -1643
rect 12667 -1723 12733 -1707
rect 12667 -1787 12668 -1723
rect 12732 -1787 12733 -1723
rect 12667 -1803 12733 -1787
rect 12667 -1867 12668 -1803
rect 12732 -1867 12733 -1803
rect 12941 -1747 13358 -1729
rect 12941 -1748 13148 -1747
rect 12941 -1806 13004 -1748
rect 12667 -1883 12733 -1867
rect 12667 -1947 12668 -1883
rect 12732 -1947 12733 -1883
rect 12667 -1963 12733 -1947
rect 12667 -2027 12668 -1963
rect 12732 -2027 12733 -1963
rect 12667 -2043 12733 -2027
rect 12667 -2107 12668 -2043
rect 12732 -2107 12733 -2043
rect 12667 -2123 12733 -2107
rect 12667 -2187 12668 -2123
rect 12732 -2187 12733 -2123
rect 12667 -2277 12733 -2187
rect 12940 -1812 13004 -1806
rect 13068 -1811 13148 -1748
rect 13212 -1748 13358 -1747
rect 13212 -1811 13279 -1748
rect 13068 -1812 13279 -1811
rect 13343 -1812 13358 -1748
rect 12061 -2342 12733 -2341
rect 12060 -2343 12733 -2342
rect 12060 -2344 12165 -2343
rect 6917 -2346 12165 -2344
rect 6917 -2355 7191 -2346
rect 6709 -2392 7191 -2355
rect 6017 -2410 7191 -2392
rect 7255 -2410 7271 -2346
rect 7335 -2410 7351 -2346
rect 7415 -2410 7431 -2346
rect 7495 -2410 7511 -2346
rect 7575 -2410 7591 -2346
rect 7655 -2410 7797 -2346
rect 7861 -2410 7877 -2346
rect 7941 -2410 7957 -2346
rect 8021 -2410 8037 -2346
rect 8101 -2410 8117 -2346
rect 8181 -2410 8197 -2346
rect 8261 -2410 8403 -2346
rect 8467 -2410 8483 -2346
rect 8547 -2410 8563 -2346
rect 8627 -2410 8643 -2346
rect 8707 -2410 8723 -2346
rect 8787 -2410 8803 -2346
rect 8867 -2410 9009 -2346
rect 9073 -2410 9089 -2346
rect 9153 -2410 9169 -2346
rect 9233 -2410 9249 -2346
rect 9313 -2410 9329 -2346
rect 9393 -2410 9409 -2346
rect 9473 -2410 9615 -2346
rect 9679 -2410 9695 -2346
rect 9759 -2410 9775 -2346
rect 9839 -2410 9855 -2346
rect 9919 -2410 9935 -2346
rect 9999 -2410 10015 -2346
rect 10079 -2410 10221 -2346
rect 10285 -2410 10301 -2346
rect 10365 -2410 10381 -2346
rect 10445 -2410 10461 -2346
rect 10525 -2410 10541 -2346
rect 10605 -2410 10621 -2346
rect 10685 -2410 10827 -2346
rect 10891 -2410 10907 -2346
rect 10971 -2410 10987 -2346
rect 11051 -2410 11067 -2346
rect 11131 -2410 11147 -2346
rect 11211 -2410 11227 -2346
rect 11291 -2410 11433 -2346
rect 11497 -2410 11513 -2346
rect 11577 -2410 11593 -2346
rect 11657 -2410 11673 -2346
rect 11737 -2410 11753 -2346
rect 11817 -2410 11833 -2346
rect 11897 -2407 12165 -2346
rect 12229 -2407 12245 -2343
rect 12309 -2407 12325 -2343
rect 12389 -2407 12405 -2343
rect 12469 -2407 12485 -2343
rect 12549 -2407 12565 -2343
rect 12629 -2344 12733 -2343
rect 12940 -2344 13358 -1812
rect 12629 -2353 13358 -2344
rect 12629 -2407 12662 -2353
rect 11897 -2410 12662 -2407
rect 6017 -2417 12662 -2410
rect 12726 -2392 13358 -2353
rect 13544 -2392 13943 3731
rect 12726 -2417 13943 -2392
rect -2 -2536 13943 -2417
<< labels >>
flabel metal1 24 -1114 78 -1068 0 FreeSans 320 0 0 0 out
port 1 nsew
flabel metal4 106 3732 13465 3796 0 FreeSans 320 0 0 0 VDD
port 2 nsew
flabel metal1 283 599 900 711 0 FreeSans 320 0 0 0 sample_delay_offset
port 4 nsew
flabel metal1 37 2391 705 2438 0 FreeSans 320 0 0 0 in
port 5 nsew
flabel metal1 0 2774 138 2808 0 FreeSans 320 0 0 0 sample_code0[3]
port 6 nsew
flabel metal1 6709 2774 6847 2808 0 FreeSans 320 0 0 0 sample_code1[3]
port 7 nsew
flabel metal1 13326 -1487 13464 -1453 0 FreeSans 320 0 0 0 sample_code2[3]
port 8 nsew
flabel metal1 6617 -1487 6755 -1453 0 FreeSans 320 0 0 0 sample_code3[3]
port 9 nsew
flabel metal1 283 795 11682 823 0 FreeSans 320 0 0 0 sample_code1[1]
port 14 nsew
flabel metal1 283 739 12538 767 0 FreeSans 320 0 0 0 sample_code1[0]
port 15 nsew
flabel metal1 283 263 984 291 0 FreeSans 320 0 0 0 sample_code3[0]
port 16 nsew
flabel metal1 283 319 1840 347 0 FreeSans 320 0 0 0 sample_code3[1]
port 17 nsew
flabel metal1 283 375 4266 403 0 FreeSans 320 0 0 0 sample_code3[2]
port 18 nsew
flabel metal1 283 431 7693 459 0 FreeSans 320 0 0 0 sample_code2[0]
port 19 nsew
flabel metal1 283 487 8549 515 0 FreeSans 320 0 0 0 sample_code2[1]
port 20 nsew
flabel metal1 283 543 10975 571 0 FreeSans 320 0 0 0 sample_code2[2]
port 22 nsew
flabel metal1 283 851 9256 879 0 FreeSans 320 0 0 0 sample_code1[2]
port 28 nsew
flabel metal4 12555 217 13464 1150 0 FreeSans 320 0 0 0 VSS
port 30 nsew
flabel metal1 283 1019 2547 1047 0 FreeSans 320 0 0 0 sample_code0[2]
port 31 nsew
flabel metal1 283 963 4973 991 0 FreeSans 320 0 0 0 sample_code0[1]
port 32 nsew
flabel metal1 283 907 5829 935 0 FreeSans 320 0 0 0 sample_code0[0]
port 34 nsew
flabel metal1 6746 2391 7414 2438 0 FreeSans 320 0 0 0 x1.IN
flabel metal1 13222 2389 13404 2435 0 FreeSans 320 0 0 0 x1.OUT
flabel metal1 6709 2774 6847 2808 0 FreeSans 320 0 0 0 x1.code[3]
flabel metal1 11624 1063 11682 2240 0 FreeSans 320 0 0 0 x1.code[1]
flabel metal1 9198 1063 9256 2240 0 FreeSans 320 0 0 0 x1.code[2]
flabel metal4 6815 3133 7233 3743 0 FreeSans 320 0 0 0 x1.VDD
flabel metal4 6843 1086 7219 2523 0 FreeSans 320 0 0 0 x1.VSS
flabel metal2 7173 2189 7609 2235 0 FreeSans 320 0 0 0 x1.code_offset
flabel metal1 12480 1062 12539 2243 0 FreeSans 320 0 0 0 x1.code[0]
flabel metal1 7357 2844 7391 2878 0 FreeSans 320 0 0 0 x1.x8.input_stack
flabel nwell 7401 3627 7435 3687 0 FreeSans 320 0 0 0 x1.x8.vdd
flabel metal1 7395 2925 7441 2937 0 FreeSans 320 0 0 0 x1.x8.output_stack
flabel poly 7334 2187 7436 2217 0 FreeSans 320 0 0 0 x1.x9.input_stack
flabel metal1 7448 1134 7482 1194 0 FreeSans 320 0 0 0 x1.x9.vss
flabel metal1 7442 2160 7488 2172 0 FreeSans 320 0 0 0 x1.x9.output_stack
flabel locali 6935 2844 6969 2878 0 FreeSans 340 0 0 0 x1.x10.Y
flabel locali 6935 2776 6969 2810 0 FreeSans 340 0 0 0 x1.x10.Y
flabel locali 6843 2776 6877 2810 0 FreeSans 340 0 0 0 x1.x10.A
flabel metal1 6800 2538 6834 2572 0 FreeSans 200 0 0 0 x1.x10.VGND
flabel metal1 6800 3082 6834 3116 0 FreeSans 200 0 0 0 x1.x10.VPWR
rlabel comment 6771 2555 6771 2555 4 x1.x10.inv_1
rlabel metal1 6771 2507 7047 2603 1 x1.x10.VGND
rlabel metal1 6771 3051 7047 3147 1 x1.x10.VPWR
flabel pwell 6800 2538 6834 2572 0 FreeSans 200 0 0 0 x1.x10.VNB
flabel nwell 6800 3082 6834 3116 0 FreeSans 200 0 0 0 x1.x10.VPB
flabel locali 7033 2844 7067 2878 0 FreeSans 340 0 0 0 x1.x11.Y
flabel locali 7033 2776 7067 2810 0 FreeSans 340 0 0 0 x1.x11.Y
flabel locali 7125 2776 7159 2810 0 FreeSans 340 0 0 0 x1.x11.A
flabel metal1 7168 2538 7202 2572 0 FreeSans 200 0 0 0 x1.x11.VGND
flabel metal1 7168 3082 7202 3116 0 FreeSans 200 0 0 0 x1.x11.VPWR
rlabel comment 7231 2555 7231 2555 6 x1.x11.inv_1
rlabel metal1 6955 2507 7231 2603 1 x1.x11.VGND
rlabel metal1 6955 3051 7231 3147 1 x1.x11.VPWR
flabel pwell 7168 2538 7202 2572 0 FreeSans 200 0 0 0 x1.x11.VNB
flabel nwell 7168 3082 7202 3116 0 FreeSans 200 0 0 0 x1.x11.VPB
flabel metal1 7999 2601 8033 2635 0 FreeSans 320 0 0 0 x1.x6.SW
flabel nwell 7443 3663 8113 3731 0 FreeSans 320 0 0 0 x1.x6.VDD
flabel pdiff 8031 2470 8089 2554 0 FreeSans 320 0 0 0 x1.x6.delay_signal
flabel metal4 7443 3662 7544 3731 0 FreeSans 320 0 0 0 x1.x6.VDD
flabel metal1 8352 2200 8386 2234 0 FreeSans 320 0 0 0 x1.x7.SW
flabel ndiff 8384 2272 8442 2356 0 FreeSans 320 0 0 0 x1.x7.delay_signal
flabel metal4 7791 1095 8463 1163 0 FreeSans 320 0 0 0 x1.x7.VSS
flabel metal1 9084 2200 9118 2234 0 FreeSans 320 0 0 0 x1.x4[3].SW
flabel ndiff 9116 2272 9174 2356 0 FreeSans 320 0 0 0 x1.x4[3].delay_signal
flabel metal4 8523 1095 9195 1163 0 FreeSans 320 0 0 0 x1.x4[3].VSS
flabel metal1 8857 2604 8891 2638 0 FreeSans 320 0 0 0 x1.x5[6].SW
flabel nwell 8777 3666 9447 3734 0 FreeSans 320 0 0 0 x1.x5[6].VDD
flabel pdiff 8801 2473 8859 2557 0 FreeSans 320 0 0 0 x1.x5[6].delay_signal
flabel metal4 9346 3665 9447 3734 0 FreeSans 320 0 0 0 x1.x5[6].VDD
flabel metal1 8731 2604 8765 2638 0 FreeSans 320 0 0 0 x1.x5[7].SW
flabel nwell 8175 3666 8845 3734 0 FreeSans 320 0 0 0 x1.x5[7].VDD
flabel pdiff 8763 2473 8821 2557 0 FreeSans 320 0 0 0 x1.x5[7].delay_signal
flabel metal4 8175 3665 8276 3734 0 FreeSans 320 0 0 0 x1.x5[7].VDD
flabel metal1 9206 2200 9240 2234 0 FreeSans 320 0 0 0 x1.x4[2].SW
flabel ndiff 9150 2272 9208 2356 0 FreeSans 320 0 0 0 x1.x4[2].delay_signal
flabel metal4 9129 1095 9801 1163 0 FreeSans 320 0 0 0 x1.x4[2].VSS
flabel metal1 9943 2604 9977 2638 0 FreeSans 320 0 0 0 x1.x5[5].SW
flabel nwell 9387 3666 10057 3734 0 FreeSans 320 0 0 0 x1.x5[5].VDD
flabel pdiff 9975 2473 10033 2557 0 FreeSans 320 0 0 0 x1.x5[5].delay_signal
flabel metal4 9387 3665 9488 3734 0 FreeSans 320 0 0 0 x1.x5[5].VDD
flabel metal1 10296 2200 10330 2234 0 FreeSans 320 0 0 0 x1.x4[1].SW
flabel ndiff 10328 2272 10386 2356 0 FreeSans 320 0 0 0 x1.x4[1].delay_signal
flabel metal4 9735 1095 10407 1163 0 FreeSans 320 0 0 0 x1.x4[1].VSS
flabel metal1 10069 2604 10103 2638 0 FreeSans 320 0 0 0 x1.x5[4].SW
flabel nwell 9989 3666 10659 3734 0 FreeSans 320 0 0 0 x1.x5[4].VDD
flabel pdiff 10013 2473 10071 2557 0 FreeSans 320 0 0 0 x1.x5[4].delay_signal
flabel metal4 10558 3665 10659 3734 0 FreeSans 320 0 0 0 x1.x5[4].VDD
flabel metal1 10418 2200 10452 2234 0 FreeSans 320 0 0 0 x1.x4[0].SW
flabel ndiff 10362 2272 10420 2356 0 FreeSans 320 0 0 0 x1.x4[0].delay_signal
flabel metal4 10341 1095 11013 1163 0 FreeSans 320 0 0 0 x1.x4[0].VSS
flabel metal1 11155 2604 11189 2638 0 FreeSans 320 0 0 0 x1.x5[3].SW
flabel nwell 10599 3666 11269 3734 0 FreeSans 320 0 0 0 x1.x5[3].VDD
flabel pdiff 11187 2473 11245 2557 0 FreeSans 320 0 0 0 x1.x5[3].delay_signal
flabel metal4 10599 3665 10700 3734 0 FreeSans 320 0 0 0 x1.x5[3].VDD
flabel metal1 11634 2200 11668 2234 0 FreeSans 320 0 0 0 x1.x3[1].SW
flabel ndiff 11666 2272 11724 2356 0 FreeSans 320 0 0 0 x1.x3[1].delay_signal
flabel metal4 11073 1095 11745 1163 0 FreeSans 320 0 0 0 x1.x3[1].VSS
flabel metal1 11281 2604 11315 2638 0 FreeSans 320 0 0 0 x1.x5[2].SW
flabel nwell 11201 3666 11871 3734 0 FreeSans 320 0 0 0 x1.x5[2].VDD
flabel pdiff 11225 2473 11283 2557 0 FreeSans 320 0 0 0 x1.x5[2].delay_signal
flabel metal4 11770 3665 11871 3734 0 FreeSans 320 0 0 0 x1.x5[2].VDD
flabel metal1 11756 2200 11790 2234 0 FreeSans 320 0 0 0 x1.x3[0].SW
flabel ndiff 11700 2272 11758 2356 0 FreeSans 320 0 0 0 x1.x3[0].delay_signal
flabel metal4 11679 1095 12351 1163 0 FreeSans 320 0 0 0 x1.x3[0].VSS
flabel metal1 12367 2604 12401 2638 0 FreeSans 320 0 0 0 x1.x5[1].SW
flabel nwell 11811 3666 12481 3734 0 FreeSans 320 0 0 0 x1.x5[1].VDD
flabel pdiff 12399 2473 12457 2557 0 FreeSans 320 0 0 0 x1.x5[1].delay_signal
flabel metal4 11811 3665 11912 3734 0 FreeSans 320 0 0 0 x1.x5[1].VDD
flabel metal1 12490 2200 12524 2234 0 FreeSans 320 0 0 0 x1.x2.SW
flabel ndiff 12434 2272 12492 2356 0 FreeSans 320 0 0 0 x1.x2.delay_signal
flabel metal4 12413 1095 13085 1163 0 FreeSans 320 0 0 0 x1.x2.VSS
flabel metal1 12493 2604 12527 2638 0 FreeSans 320 0 0 0 x1.x5[0].SW
flabel nwell 12413 3666 13083 3734 0 FreeSans 320 0 0 0 x1.x5[0].VDD
flabel pdiff 12437 2473 12495 2557 0 FreeSans 320 0 0 0 x1.x5[0].delay_signal
flabel metal4 12982 3665 13083 3734 0 FreeSans 320 0 0 0 x1.x5[0].VDD
flabel metal1 12759 -1117 13427 -1070 0 FreeSans 320 0 0 0 x2.IN
flabel metal1 6769 -1114 6951 -1068 0 FreeSans 320 0 0 0 x2.OUT
flabel metal1 13326 -1487 13464 -1453 0 FreeSans 320 0 0 0 x2.code[3]
flabel metal1 8491 -919 8549 258 0 FreeSans 320 0 0 0 x2.code[1]
flabel metal1 10917 -919 10975 258 0 FreeSans 320 0 0 0 x2.code[2]
flabel metal4 12940 -2422 13358 -1812 0 FreeSans 320 0 0 0 x2.VDD
flabel metal4 12954 -1202 13330 235 0 FreeSans 320 0 0 0 x2.VSS
flabel metal2 12564 -914 13000 -868 0 FreeSans 320 0 0 0 x2.code_offset
flabel metal1 7634 -922 7693 259 0 FreeSans 320 0 0 0 x2.code[0]
flabel metal1 12782 -1557 12816 -1523 0 FreeSans 320 0 0 0 x2.x8.input_stack
flabel nwell 12738 -2366 12772 -2306 0 FreeSans 320 0 0 0 x2.x8.vdd
flabel metal1 12732 -1616 12778 -1604 0 FreeSans 320 0 0 0 x2.x8.output_stack
flabel poly 12737 -896 12839 -866 0 FreeSans 320 0 0 0 x2.x9.input_stack
flabel metal1 12691 127 12725 187 0 FreeSans 320 0 0 0 x2.x9.vss
flabel metal1 12685 -851 12731 -839 0 FreeSans 320 0 0 0 x2.x9.output_stack
flabel locali 13204 -1557 13238 -1523 0 FreeSans 340 0 0 0 x2.x10.Y
flabel locali 13204 -1489 13238 -1455 0 FreeSans 340 0 0 0 x2.x10.Y
flabel locali 13296 -1489 13330 -1455 0 FreeSans 340 0 0 0 x2.x10.A
flabel metal1 13339 -1251 13373 -1217 0 FreeSans 200 0 0 0 x2.x10.VGND
flabel metal1 13339 -1795 13373 -1761 0 FreeSans 200 0 0 0 x2.x10.VPWR
rlabel comment 13402 -1234 13402 -1234 8 x2.x10.inv_1
rlabel metal1 13126 -1282 13402 -1186 5 x2.x10.VGND
rlabel metal1 13126 -1826 13402 -1730 5 x2.x10.VPWR
flabel pwell 13339 -1251 13373 -1217 0 FreeSans 200 0 0 0 x2.x10.VNB
flabel nwell 13339 -1795 13373 -1761 0 FreeSans 200 0 0 0 x2.x10.VPB
flabel locali 13106 -1557 13140 -1523 0 FreeSans 340 0 0 0 x2.x11.Y
flabel locali 13106 -1489 13140 -1455 0 FreeSans 340 0 0 0 x2.x11.Y
flabel locali 13014 -1489 13048 -1455 0 FreeSans 340 0 0 0 x2.x11.A
flabel metal1 12971 -1251 13005 -1217 0 FreeSans 200 0 0 0 x2.x11.VGND
flabel metal1 12971 -1795 13005 -1761 0 FreeSans 200 0 0 0 x2.x11.VPWR
rlabel comment 12942 -1234 12942 -1234 2 x2.x11.inv_1
rlabel metal1 12942 -1282 13218 -1186 5 x2.x11.VGND
rlabel metal1 12942 -1826 13218 -1730 5 x2.x11.VPWR
flabel pwell 12971 -1251 13005 -1217 0 FreeSans 200 0 0 0 x2.x11.VNB
flabel nwell 12971 -1795 13005 -1761 0 FreeSans 200 0 0 0 x2.x11.VPB
flabel metal1 12140 -1314 12174 -1280 0 FreeSans 320 0 0 0 x2.x6.SW
flabel nwell 12060 -2410 12730 -2342 0 FreeSans 320 0 0 0 x2.x6.VDD
flabel pdiff 12084 -1233 12142 -1149 0 FreeSans 320 0 0 0 x2.x6.delay_signal
flabel metal4 12629 -2410 12730 -2341 0 FreeSans 320 0 0 0 x2.x6.VDD
flabel metal1 11787 -913 11821 -879 0 FreeSans 320 0 0 0 x2.x7.SW
flabel ndiff 11731 -1035 11789 -951 0 FreeSans 320 0 0 0 x2.x7.delay_signal
flabel metal4 11710 158 12382 226 0 FreeSans 320 0 0 0 x2.x7.VSS
flabel metal1 11055 -913 11089 -879 0 FreeSans 320 0 0 0 x2.x4[3].SW
flabel ndiff 10999 -1035 11057 -951 0 FreeSans 320 0 0 0 x2.x4[3].delay_signal
flabel metal4 10978 158 11650 226 0 FreeSans 320 0 0 0 x2.x4[3].VSS
flabel metal1 11282 -1317 11316 -1283 0 FreeSans 320 0 0 0 x2.x5[6].SW
flabel nwell 10726 -2413 11396 -2345 0 FreeSans 320 0 0 0 x2.x5[6].VDD
flabel pdiff 11314 -1236 11372 -1152 0 FreeSans 320 0 0 0 x2.x5[6].delay_signal
flabel metal4 10726 -2413 10827 -2344 0 FreeSans 320 0 0 0 x2.x5[6].VDD
flabel metal1 11408 -1317 11442 -1283 0 FreeSans 320 0 0 0 x2.x5[7].SW
flabel nwell 11328 -2413 11998 -2345 0 FreeSans 320 0 0 0 x2.x5[7].VDD
flabel pdiff 11352 -1236 11410 -1152 0 FreeSans 320 0 0 0 x2.x5[7].delay_signal
flabel metal4 11897 -2413 11998 -2344 0 FreeSans 320 0 0 0 x2.x5[7].VDD
flabel metal1 10933 -913 10967 -879 0 FreeSans 320 0 0 0 x2.x4[2].SW
flabel ndiff 10965 -1035 11023 -951 0 FreeSans 320 0 0 0 x2.x4[2].delay_signal
flabel metal4 10372 158 11044 226 0 FreeSans 320 0 0 0 x2.x4[2].VSS
flabel metal1 10196 -1317 10230 -1283 0 FreeSans 320 0 0 0 x2.x5[5].SW
flabel nwell 10116 -2413 10786 -2345 0 FreeSans 320 0 0 0 x2.x5[5].VDD
flabel pdiff 10140 -1236 10198 -1152 0 FreeSans 320 0 0 0 x2.x5[5].delay_signal
flabel metal4 10685 -2413 10786 -2344 0 FreeSans 320 0 0 0 x2.x5[5].VDD
flabel metal1 9843 -913 9877 -879 0 FreeSans 320 0 0 0 x2.x4[1].SW
flabel ndiff 9787 -1035 9845 -951 0 FreeSans 320 0 0 0 x2.x4[1].delay_signal
flabel metal4 9766 158 10438 226 0 FreeSans 320 0 0 0 x2.x4[1].VSS
flabel metal1 10070 -1317 10104 -1283 0 FreeSans 320 0 0 0 x2.x5[4].SW
flabel nwell 9514 -2413 10184 -2345 0 FreeSans 320 0 0 0 x2.x5[4].VDD
flabel pdiff 10102 -1236 10160 -1152 0 FreeSans 320 0 0 0 x2.x5[4].delay_signal
flabel metal4 9514 -2413 9615 -2344 0 FreeSans 320 0 0 0 x2.x5[4].VDD
flabel metal1 9721 -913 9755 -879 0 FreeSans 320 0 0 0 x2.x4[0].SW
flabel ndiff 9753 -1035 9811 -951 0 FreeSans 320 0 0 0 x2.x4[0].delay_signal
flabel metal4 9160 158 9832 226 0 FreeSans 320 0 0 0 x2.x4[0].VSS
flabel metal1 8984 -1317 9018 -1283 0 FreeSans 320 0 0 0 x2.x5[3].SW
flabel nwell 8904 -2413 9574 -2345 0 FreeSans 320 0 0 0 x2.x5[3].VDD
flabel pdiff 8928 -1236 8986 -1152 0 FreeSans 320 0 0 0 x2.x5[3].delay_signal
flabel metal4 9473 -2413 9574 -2344 0 FreeSans 320 0 0 0 x2.x5[3].VDD
flabel metal1 8505 -913 8539 -879 0 FreeSans 320 0 0 0 x2.x3[1].SW
flabel ndiff 8449 -1035 8507 -951 0 FreeSans 320 0 0 0 x2.x3[1].delay_signal
flabel metal4 8428 158 9100 226 0 FreeSans 320 0 0 0 x2.x3[1].VSS
flabel metal1 8858 -1317 8892 -1283 0 FreeSans 320 0 0 0 x2.x5[2].SW
flabel nwell 8302 -2413 8972 -2345 0 FreeSans 320 0 0 0 x2.x5[2].VDD
flabel pdiff 8890 -1236 8948 -1152 0 FreeSans 320 0 0 0 x2.x5[2].delay_signal
flabel metal4 8302 -2413 8403 -2344 0 FreeSans 320 0 0 0 x2.x5[2].VDD
flabel metal1 8383 -913 8417 -879 0 FreeSans 320 0 0 0 x2.x3[0].SW
flabel ndiff 8415 -1035 8473 -951 0 FreeSans 320 0 0 0 x2.x3[0].delay_signal
flabel metal4 7822 158 8494 226 0 FreeSans 320 0 0 0 x2.x3[0].VSS
flabel metal1 7772 -1317 7806 -1283 0 FreeSans 320 0 0 0 x2.x5[1].SW
flabel nwell 7692 -2413 8362 -2345 0 FreeSans 320 0 0 0 x2.x5[1].VDD
flabel pdiff 7716 -1236 7774 -1152 0 FreeSans 320 0 0 0 x2.x5[1].delay_signal
flabel metal4 8261 -2413 8362 -2344 0 FreeSans 320 0 0 0 x2.x5[1].VDD
flabel metal1 7649 -913 7683 -879 0 FreeSans 320 0 0 0 x2.x2.SW
flabel ndiff 7681 -1035 7739 -951 0 FreeSans 320 0 0 0 x2.x2.delay_signal
flabel metal4 7088 158 7760 226 0 FreeSans 320 0 0 0 x2.x2.VSS
flabel metal1 7646 -1317 7680 -1283 0 FreeSans 320 0 0 0 x2.x5[0].SW
flabel nwell 7090 -2413 7760 -2345 0 FreeSans 320 0 0 0 x2.x5[0].VDD
flabel pdiff 7678 -1236 7736 -1152 0 FreeSans 320 0 0 0 x2.x5[0].delay_signal
flabel metal4 7090 -2413 7191 -2344 0 FreeSans 320 0 0 0 x2.x5[0].VDD
flabel metal1 6050 -1117 6718 -1070 0 FreeSans 320 0 0 0 x3.IN
flabel metal1 60 -1114 242 -1068 0 FreeSans 320 0 0 0 x3.OUT
flabel metal1 6617 -1487 6755 -1453 0 FreeSans 320 0 0 0 x3.code[3]
flabel metal1 1782 -919 1840 258 0 FreeSans 320 0 0 0 x3.code[1]
flabel metal1 4208 -919 4266 258 0 FreeSans 320 0 0 0 x3.code[2]
flabel metal4 6231 -2422 6649 -1812 0 FreeSans 320 0 0 0 x3.VDD
flabel metal4 6245 -1202 6621 235 0 FreeSans 320 0 0 0 x3.VSS
flabel metal2 5855 -914 6291 -868 0 FreeSans 320 0 0 0 x3.code_offset
flabel metal1 925 -922 984 259 0 FreeSans 320 0 0 0 x3.code[0]
flabel metal1 6073 -1557 6107 -1523 0 FreeSans 320 0 0 0 x3.x8.input_stack
flabel nwell 6029 -2366 6063 -2306 0 FreeSans 320 0 0 0 x3.x8.vdd
flabel metal1 6023 -1616 6069 -1604 0 FreeSans 320 0 0 0 x3.x8.output_stack
flabel poly 6028 -896 6130 -866 0 FreeSans 320 0 0 0 x3.x9.input_stack
flabel metal1 5982 127 6016 187 0 FreeSans 320 0 0 0 x3.x9.vss
flabel metal1 5976 -851 6022 -839 0 FreeSans 320 0 0 0 x3.x9.output_stack
flabel locali 6495 -1557 6529 -1523 0 FreeSans 340 0 0 0 x3.x10.Y
flabel locali 6495 -1489 6529 -1455 0 FreeSans 340 0 0 0 x3.x10.Y
flabel locali 6587 -1489 6621 -1455 0 FreeSans 340 0 0 0 x3.x10.A
flabel metal1 6630 -1251 6664 -1217 0 FreeSans 200 0 0 0 x3.x10.VGND
flabel metal1 6630 -1795 6664 -1761 0 FreeSans 200 0 0 0 x3.x10.VPWR
rlabel comment 6693 -1234 6693 -1234 8 x3.x10.inv_1
rlabel metal1 6417 -1282 6693 -1186 5 x3.x10.VGND
rlabel metal1 6417 -1826 6693 -1730 5 x3.x10.VPWR
flabel pwell 6630 -1251 6664 -1217 0 FreeSans 200 0 0 0 x3.x10.VNB
flabel nwell 6630 -1795 6664 -1761 0 FreeSans 200 0 0 0 x3.x10.VPB
flabel locali 6397 -1557 6431 -1523 0 FreeSans 340 0 0 0 x3.x11.Y
flabel locali 6397 -1489 6431 -1455 0 FreeSans 340 0 0 0 x3.x11.Y
flabel locali 6305 -1489 6339 -1455 0 FreeSans 340 0 0 0 x3.x11.A
flabel metal1 6262 -1251 6296 -1217 0 FreeSans 200 0 0 0 x3.x11.VGND
flabel metal1 6262 -1795 6296 -1761 0 FreeSans 200 0 0 0 x3.x11.VPWR
rlabel comment 6233 -1234 6233 -1234 2 x3.x11.inv_1
rlabel metal1 6233 -1282 6509 -1186 5 x3.x11.VGND
rlabel metal1 6233 -1826 6509 -1730 5 x3.x11.VPWR
flabel pwell 6262 -1251 6296 -1217 0 FreeSans 200 0 0 0 x3.x11.VNB
flabel nwell 6262 -1795 6296 -1761 0 FreeSans 200 0 0 0 x3.x11.VPB
flabel metal1 5431 -1314 5465 -1280 0 FreeSans 320 0 0 0 x3.x6.SW
flabel nwell 5351 -2410 6021 -2342 0 FreeSans 320 0 0 0 x3.x6.VDD
flabel pdiff 5375 -1233 5433 -1149 0 FreeSans 320 0 0 0 x3.x6.delay_signal
flabel metal4 5920 -2410 6021 -2341 0 FreeSans 320 0 0 0 x3.x6.VDD
flabel metal1 5078 -913 5112 -879 0 FreeSans 320 0 0 0 x3.x7.SW
flabel ndiff 5022 -1035 5080 -951 0 FreeSans 320 0 0 0 x3.x7.delay_signal
flabel metal4 5001 158 5673 226 0 FreeSans 320 0 0 0 x3.x7.VSS
flabel metal1 4346 -913 4380 -879 0 FreeSans 320 0 0 0 x3.x4[3].SW
flabel ndiff 4290 -1035 4348 -951 0 FreeSans 320 0 0 0 x3.x4[3].delay_signal
flabel metal4 4269 158 4941 226 0 FreeSans 320 0 0 0 x3.x4[3].VSS
flabel metal1 4573 -1317 4607 -1283 0 FreeSans 320 0 0 0 x3.x5[6].SW
flabel nwell 4017 -2413 4687 -2345 0 FreeSans 320 0 0 0 x3.x5[6].VDD
flabel pdiff 4605 -1236 4663 -1152 0 FreeSans 320 0 0 0 x3.x5[6].delay_signal
flabel metal4 4017 -2413 4118 -2344 0 FreeSans 320 0 0 0 x3.x5[6].VDD
flabel metal1 4699 -1317 4733 -1283 0 FreeSans 320 0 0 0 x3.x5[7].SW
flabel nwell 4619 -2413 5289 -2345 0 FreeSans 320 0 0 0 x3.x5[7].VDD
flabel pdiff 4643 -1236 4701 -1152 0 FreeSans 320 0 0 0 x3.x5[7].delay_signal
flabel metal4 5188 -2413 5289 -2344 0 FreeSans 320 0 0 0 x3.x5[7].VDD
flabel metal1 4224 -913 4258 -879 0 FreeSans 320 0 0 0 x3.x4[2].SW
flabel ndiff 4256 -1035 4314 -951 0 FreeSans 320 0 0 0 x3.x4[2].delay_signal
flabel metal4 3663 158 4335 226 0 FreeSans 320 0 0 0 x3.x4[2].VSS
flabel metal1 3487 -1317 3521 -1283 0 FreeSans 320 0 0 0 x3.x5[5].SW
flabel nwell 3407 -2413 4077 -2345 0 FreeSans 320 0 0 0 x3.x5[5].VDD
flabel pdiff 3431 -1236 3489 -1152 0 FreeSans 320 0 0 0 x3.x5[5].delay_signal
flabel metal4 3976 -2413 4077 -2344 0 FreeSans 320 0 0 0 x3.x5[5].VDD
flabel metal1 3134 -913 3168 -879 0 FreeSans 320 0 0 0 x3.x4[1].SW
flabel ndiff 3078 -1035 3136 -951 0 FreeSans 320 0 0 0 x3.x4[1].delay_signal
flabel metal4 3057 158 3729 226 0 FreeSans 320 0 0 0 x3.x4[1].VSS
flabel metal1 3361 -1317 3395 -1283 0 FreeSans 320 0 0 0 x3.x5[4].SW
flabel nwell 2805 -2413 3475 -2345 0 FreeSans 320 0 0 0 x3.x5[4].VDD
flabel pdiff 3393 -1236 3451 -1152 0 FreeSans 320 0 0 0 x3.x5[4].delay_signal
flabel metal4 2805 -2413 2906 -2344 0 FreeSans 320 0 0 0 x3.x5[4].VDD
flabel metal1 3012 -913 3046 -879 0 FreeSans 320 0 0 0 x3.x4[0].SW
flabel ndiff 3044 -1035 3102 -951 0 FreeSans 320 0 0 0 x3.x4[0].delay_signal
flabel metal4 2451 158 3123 226 0 FreeSans 320 0 0 0 x3.x4[0].VSS
flabel metal1 2275 -1317 2309 -1283 0 FreeSans 320 0 0 0 x3.x5[3].SW
flabel nwell 2195 -2413 2865 -2345 0 FreeSans 320 0 0 0 x3.x5[3].VDD
flabel pdiff 2219 -1236 2277 -1152 0 FreeSans 320 0 0 0 x3.x5[3].delay_signal
flabel metal4 2764 -2413 2865 -2344 0 FreeSans 320 0 0 0 x3.x5[3].VDD
flabel metal1 1796 -913 1830 -879 0 FreeSans 320 0 0 0 x3.x3[1].SW
flabel ndiff 1740 -1035 1798 -951 0 FreeSans 320 0 0 0 x3.x3[1].delay_signal
flabel metal4 1719 158 2391 226 0 FreeSans 320 0 0 0 x3.x3[1].VSS
flabel metal1 2149 -1317 2183 -1283 0 FreeSans 320 0 0 0 x3.x5[2].SW
flabel nwell 1593 -2413 2263 -2345 0 FreeSans 320 0 0 0 x3.x5[2].VDD
flabel pdiff 2181 -1236 2239 -1152 0 FreeSans 320 0 0 0 x3.x5[2].delay_signal
flabel metal4 1593 -2413 1694 -2344 0 FreeSans 320 0 0 0 x3.x5[2].VDD
flabel metal1 1674 -913 1708 -879 0 FreeSans 320 0 0 0 x3.x3[0].SW
flabel ndiff 1706 -1035 1764 -951 0 FreeSans 320 0 0 0 x3.x3[0].delay_signal
flabel metal4 1113 158 1785 226 0 FreeSans 320 0 0 0 x3.x3[0].VSS
flabel metal1 1063 -1317 1097 -1283 0 FreeSans 320 0 0 0 x3.x5[1].SW
flabel nwell 983 -2413 1653 -2345 0 FreeSans 320 0 0 0 x3.x5[1].VDD
flabel pdiff 1007 -1236 1065 -1152 0 FreeSans 320 0 0 0 x3.x5[1].delay_signal
flabel metal4 1552 -2413 1653 -2344 0 FreeSans 320 0 0 0 x3.x5[1].VDD
flabel metal1 940 -913 974 -879 0 FreeSans 320 0 0 0 x3.x2.SW
flabel ndiff 972 -1035 1030 -951 0 FreeSans 320 0 0 0 x3.x2.delay_signal
flabel metal4 379 158 1051 226 0 FreeSans 320 0 0 0 x3.x2.VSS
flabel metal1 937 -1317 971 -1283 0 FreeSans 320 0 0 0 x3.x5[0].SW
flabel nwell 381 -2413 1051 -2345 0 FreeSans 320 0 0 0 x3.x5[0].VDD
flabel pdiff 969 -1236 1027 -1152 0 FreeSans 320 0 0 0 x3.x5[0].delay_signal
flabel metal4 381 -2413 482 -2344 0 FreeSans 320 0 0 0 x3.x5[0].VDD
flabel metal1 37 2391 705 2438 0 FreeSans 320 0 0 0 x4.IN
flabel metal1 6513 2389 6695 2435 0 FreeSans 320 0 0 0 x4.OUT
flabel metal1 0 2774 138 2808 0 FreeSans 320 0 0 0 x4.code[3]
flabel metal1 4915 1063 4973 2240 0 FreeSans 320 0 0 0 x4.code[1]
flabel metal1 2489 1063 2547 2240 0 FreeSans 320 0 0 0 x4.code[2]
flabel metal4 106 3133 524 3743 0 FreeSans 320 0 0 0 x4.VDD
flabel metal4 134 1086 510 2523 0 FreeSans 320 0 0 0 x4.VSS
flabel metal2 464 2189 900 2235 0 FreeSans 320 0 0 0 x4.code_offset
flabel metal1 5771 1062 5830 2243 0 FreeSans 320 0 0 0 x4.code[0]
flabel metal1 648 2844 682 2878 0 FreeSans 320 0 0 0 x4.x8.input_stack
flabel nwell 692 3627 726 3687 0 FreeSans 320 0 0 0 x4.x8.vdd
flabel metal1 686 2925 732 2937 0 FreeSans 320 0 0 0 x4.x8.output_stack
flabel poly 625 2187 727 2217 0 FreeSans 320 0 0 0 x4.x9.input_stack
flabel metal1 739 1134 773 1194 0 FreeSans 320 0 0 0 x4.x9.vss
flabel metal1 733 2160 779 2172 0 FreeSans 320 0 0 0 x4.x9.output_stack
flabel locali 226 2844 260 2878 0 FreeSans 340 0 0 0 x4.x10.Y
flabel locali 226 2776 260 2810 0 FreeSans 340 0 0 0 x4.x10.Y
flabel locali 134 2776 168 2810 0 FreeSans 340 0 0 0 x4.x10.A
flabel metal1 91 2538 125 2572 0 FreeSans 200 0 0 0 x4.x10.VGND
flabel metal1 91 3082 125 3116 0 FreeSans 200 0 0 0 x4.x10.VPWR
rlabel comment 62 2555 62 2555 4 x4.x10.inv_1
rlabel metal1 62 2507 338 2603 1 x4.x10.VGND
rlabel metal1 62 3051 338 3147 1 x4.x10.VPWR
flabel pwell 91 2538 125 2572 0 FreeSans 200 0 0 0 x4.x10.VNB
flabel nwell 91 3082 125 3116 0 FreeSans 200 0 0 0 x4.x10.VPB
flabel locali 324 2844 358 2878 0 FreeSans 340 0 0 0 x4.x11.Y
flabel locali 324 2776 358 2810 0 FreeSans 340 0 0 0 x4.x11.Y
flabel locali 416 2776 450 2810 0 FreeSans 340 0 0 0 x4.x11.A
flabel metal1 459 2538 493 2572 0 FreeSans 200 0 0 0 x4.x11.VGND
flabel metal1 459 3082 493 3116 0 FreeSans 200 0 0 0 x4.x11.VPWR
rlabel comment 522 2555 522 2555 6 x4.x11.inv_1
rlabel metal1 246 2507 522 2603 1 x4.x11.VGND
rlabel metal1 246 3051 522 3147 1 x4.x11.VPWR
flabel pwell 459 2538 493 2572 0 FreeSans 200 0 0 0 x4.x11.VNB
flabel nwell 459 3082 493 3116 0 FreeSans 200 0 0 0 x4.x11.VPB
flabel metal1 1290 2601 1324 2635 0 FreeSans 320 0 0 0 x4.x6.SW
flabel nwell 734 3663 1404 3731 0 FreeSans 320 0 0 0 x4.x6.VDD
flabel pdiff 1322 2470 1380 2554 0 FreeSans 320 0 0 0 x4.x6.delay_signal
flabel metal4 734 3662 835 3731 0 FreeSans 320 0 0 0 x4.x6.VDD
flabel metal1 1643 2200 1677 2234 0 FreeSans 320 0 0 0 x4.x7.SW
flabel ndiff 1675 2272 1733 2356 0 FreeSans 320 0 0 0 x4.x7.delay_signal
flabel metal4 1082 1095 1754 1163 0 FreeSans 320 0 0 0 x4.x7.VSS
flabel metal1 2375 2200 2409 2234 0 FreeSans 320 0 0 0 x4.x4[3].SW
flabel ndiff 2407 2272 2465 2356 0 FreeSans 320 0 0 0 x4.x4[3].delay_signal
flabel metal4 1814 1095 2486 1163 0 FreeSans 320 0 0 0 x4.x4[3].VSS
flabel metal1 2148 2604 2182 2638 0 FreeSans 320 0 0 0 x4.x5[6].SW
flabel nwell 2068 3666 2738 3734 0 FreeSans 320 0 0 0 x4.x5[6].VDD
flabel pdiff 2092 2473 2150 2557 0 FreeSans 320 0 0 0 x4.x5[6].delay_signal
flabel metal4 2637 3665 2738 3734 0 FreeSans 320 0 0 0 x4.x5[6].VDD
flabel metal1 2022 2604 2056 2638 0 FreeSans 320 0 0 0 x4.x5[7].SW
flabel nwell 1466 3666 2136 3734 0 FreeSans 320 0 0 0 x4.x5[7].VDD
flabel pdiff 2054 2473 2112 2557 0 FreeSans 320 0 0 0 x4.x5[7].delay_signal
flabel metal4 1466 3665 1567 3734 0 FreeSans 320 0 0 0 x4.x5[7].VDD
flabel metal1 2497 2200 2531 2234 0 FreeSans 320 0 0 0 x4.x4[2].SW
flabel ndiff 2441 2272 2499 2356 0 FreeSans 320 0 0 0 x4.x4[2].delay_signal
flabel metal4 2420 1095 3092 1163 0 FreeSans 320 0 0 0 x4.x4[2].VSS
flabel metal1 3234 2604 3268 2638 0 FreeSans 320 0 0 0 x4.x5[5].SW
flabel nwell 2678 3666 3348 3734 0 FreeSans 320 0 0 0 x4.x5[5].VDD
flabel pdiff 3266 2473 3324 2557 0 FreeSans 320 0 0 0 x4.x5[5].delay_signal
flabel metal4 2678 3665 2779 3734 0 FreeSans 320 0 0 0 x4.x5[5].VDD
flabel metal1 3587 2200 3621 2234 0 FreeSans 320 0 0 0 x4.x4[1].SW
flabel ndiff 3619 2272 3677 2356 0 FreeSans 320 0 0 0 x4.x4[1].delay_signal
flabel metal4 3026 1095 3698 1163 0 FreeSans 320 0 0 0 x4.x4[1].VSS
flabel metal1 3360 2604 3394 2638 0 FreeSans 320 0 0 0 x4.x5[4].SW
flabel nwell 3280 3666 3950 3734 0 FreeSans 320 0 0 0 x4.x5[4].VDD
flabel pdiff 3304 2473 3362 2557 0 FreeSans 320 0 0 0 x4.x5[4].delay_signal
flabel metal4 3849 3665 3950 3734 0 FreeSans 320 0 0 0 x4.x5[4].VDD
flabel metal1 3709 2200 3743 2234 0 FreeSans 320 0 0 0 x4.x4[0].SW
flabel ndiff 3653 2272 3711 2356 0 FreeSans 320 0 0 0 x4.x4[0].delay_signal
flabel metal4 3632 1095 4304 1163 0 FreeSans 320 0 0 0 x4.x4[0].VSS
flabel metal1 4446 2604 4480 2638 0 FreeSans 320 0 0 0 x4.x5[3].SW
flabel nwell 3890 3666 4560 3734 0 FreeSans 320 0 0 0 x4.x5[3].VDD
flabel pdiff 4478 2473 4536 2557 0 FreeSans 320 0 0 0 x4.x5[3].delay_signal
flabel metal4 3890 3665 3991 3734 0 FreeSans 320 0 0 0 x4.x5[3].VDD
flabel metal1 4925 2200 4959 2234 0 FreeSans 320 0 0 0 x4.x3[1].SW
flabel ndiff 4957 2272 5015 2356 0 FreeSans 320 0 0 0 x4.x3[1].delay_signal
flabel metal4 4364 1095 5036 1163 0 FreeSans 320 0 0 0 x4.x3[1].VSS
flabel metal1 4572 2604 4606 2638 0 FreeSans 320 0 0 0 x4.x5[2].SW
flabel nwell 4492 3666 5162 3734 0 FreeSans 320 0 0 0 x4.x5[2].VDD
flabel pdiff 4516 2473 4574 2557 0 FreeSans 320 0 0 0 x4.x5[2].delay_signal
flabel metal4 5061 3665 5162 3734 0 FreeSans 320 0 0 0 x4.x5[2].VDD
flabel metal1 5047 2200 5081 2234 0 FreeSans 320 0 0 0 x4.x3[0].SW
flabel ndiff 4991 2272 5049 2356 0 FreeSans 320 0 0 0 x4.x3[0].delay_signal
flabel metal4 4970 1095 5642 1163 0 FreeSans 320 0 0 0 x4.x3[0].VSS
flabel metal1 5658 2604 5692 2638 0 FreeSans 320 0 0 0 x4.x5[1].SW
flabel nwell 5102 3666 5772 3734 0 FreeSans 320 0 0 0 x4.x5[1].VDD
flabel pdiff 5690 2473 5748 2557 0 FreeSans 320 0 0 0 x4.x5[1].delay_signal
flabel metal4 5102 3665 5203 3734 0 FreeSans 320 0 0 0 x4.x5[1].VDD
flabel metal1 5781 2200 5815 2234 0 FreeSans 320 0 0 0 x4.x2.SW
flabel ndiff 5725 2272 5783 2356 0 FreeSans 320 0 0 0 x4.x2.delay_signal
flabel metal4 5704 1095 6376 1163 0 FreeSans 320 0 0 0 x4.x2.VSS
flabel metal1 5784 2604 5818 2638 0 FreeSans 320 0 0 0 x4.x5[0].SW
flabel nwell 5704 3666 6374 3734 0 FreeSans 320 0 0 0 x4.x5[0].VDD
flabel pdiff 5728 2473 5786 2557 0 FreeSans 320 0 0 0 x4.x5[0].delay_signal
flabel metal4 6273 3665 6374 3734 0 FreeSans 320 0 0 0 x4.x5[0].VDD
<< end >>
