magic
tech sky130A
magscale 1 2
timestamp 1697028858
<< error_s >>
rect 476 -710 6752 -674
rect 476 -852 512 -710
rect 1018 -778 2056 -776
rect 1018 -812 3090 -778
rect 1018 -852 1054 -812
rect 2020 -814 3090 -812
rect 3054 -852 3090 -814
rect 3220 -828 3642 -792
rect 4322 -828 4972 -792
rect 3220 -852 3344 -828
rect 3606 -852 4068 -828
rect 4322 -852 4358 -828
rect 4874 -844 4972 -828
rect 4936 -852 4972 -844
rect 5128 -852 5550 -844
rect 6716 -852 6752 -710
rect 476 -888 1018 -852
rect 3090 -888 3344 -852
rect 4068 -888 4322 -852
rect 4972 -888 5226 -852
rect 5550 -878 6752 -852
rect 6028 -888 6752 -878
rect 3220 -1398 3344 -888
rect 5128 -1398 5226 -888
rect 1200 -1442 1258 -1436
rect 1400 -1442 1458 -1436
rect 1816 -1442 1874 -1436
rect 1200 -1476 1212 -1442
rect 1400 -1476 1412 -1442
rect 1816 -1476 1828 -1442
rect 2228 -1444 2286 -1438
rect 2648 -1444 2706 -1438
rect 2850 -1444 2908 -1438
rect 1200 -1482 1258 -1476
rect 1400 -1482 1458 -1476
rect 1816 -1482 1874 -1476
rect 2228 -1478 2240 -1444
rect 2648 -1478 2660 -1444
rect 2850 -1478 2862 -1444
rect 2228 -1484 2286 -1478
rect 2648 -1484 2706 -1478
rect 2850 -1484 2908 -1478
rect 1808 -1722 1866 -1716
rect 1808 -1756 1820 -1722
rect 2274 -1734 2332 -1728
rect 2062 -1754 2120 -1748
rect 1808 -1762 1866 -1756
rect 2062 -1788 2074 -1754
rect 2274 -1768 2286 -1734
rect 2274 -1774 2332 -1768
rect 2062 -1794 2120 -1788
rect 4496 -1834 4554 -1828
rect 4716 -1834 4774 -1828
rect 4496 -1868 4508 -1834
rect 4716 -1868 4728 -1834
rect 4496 -1874 4554 -1868
rect 4716 -1874 4774 -1868
rect 2712 -1890 2770 -1884
rect 2904 -1890 2962 -1884
rect 2712 -1924 2724 -1890
rect 2904 -1924 2916 -1890
rect 1340 -1932 1398 -1926
rect 1532 -1932 1590 -1926
rect 2712 -1930 2770 -1924
rect 2904 -1930 2962 -1924
rect 1340 -1966 1352 -1932
rect 1532 -1966 1544 -1932
rect 1340 -1972 1398 -1966
rect 1532 -1972 1590 -1966
rect 4562 -2074 4620 -2068
rect 4762 -2074 4820 -2068
rect 4562 -2108 4574 -2074
rect 4762 -2108 4774 -2074
rect 4562 -2114 4620 -2108
rect 4762 -2114 4820 -2108
rect 2616 -2400 2674 -2394
rect 2808 -2400 2866 -2394
rect 2616 -2434 2628 -2400
rect 2808 -2434 2820 -2400
rect 1244 -2442 1302 -2436
rect 1436 -2442 1494 -2436
rect 2616 -2440 2674 -2434
rect 2808 -2440 2866 -2434
rect 1244 -2476 1256 -2442
rect 1436 -2476 1448 -2442
rect 1244 -2482 1302 -2476
rect 1436 -2482 1494 -2476
rect 5064 -2566 5204 -2474
rect 5318 -3080 5458 -2566
rect 7032 -2715 7062 -2686
<< nsubdiff >>
rect 512 -852 6716 -710
<< poly >>
rect 3416 -1568 3446 -1196
rect 4500 -1226 4566 -1210
rect 4500 -1260 4516 -1226
rect 4550 -1260 4566 -1226
rect 4500 -1278 4566 -1260
rect 4728 -1226 4794 -1210
rect 4728 -1260 4744 -1226
rect 4778 -1260 4794 -1226
rect 4728 -1280 4794 -1260
rect 5324 -1622 5354 -1231
rect 3414 -2683 3444 -2268
rect 4576 -2682 4606 -2344
rect 4776 -2682 4806 -2305
rect 4978 -2394 5008 -2296
rect 4942 -2410 5008 -2394
rect 4942 -2444 4958 -2410
rect 4992 -2444 5008 -2410
rect 4942 -2460 5008 -2444
rect 4978 -2682 5008 -2460
rect 5514 -2785 5544 -2337
rect 7032 -2716 7062 -2715
<< polycont >>
rect 4516 -1260 4550 -1226
rect 4744 -1260 4778 -1226
rect 4958 -2444 4992 -2410
<< locali >>
rect 508 -730 6712 -710
rect 508 -732 3130 -730
rect 508 -836 538 -732
rect 646 -836 754 -732
rect 862 -836 970 -732
rect 1078 -836 1186 -732
rect 1294 -836 1402 -732
rect 1510 -836 1618 -732
rect 1726 -836 1834 -732
rect 1942 -836 2050 -732
rect 2158 -836 2266 -732
rect 2374 -836 2482 -732
rect 2590 -836 2698 -732
rect 2806 -836 2914 -732
rect 3022 -834 3130 -732
rect 3238 -834 3346 -730
rect 3454 -834 3562 -730
rect 3670 -834 3778 -730
rect 3886 -834 3994 -730
rect 4102 -834 4210 -730
rect 4318 -834 4426 -730
rect 4534 -834 4642 -730
rect 4750 -834 4858 -730
rect 4966 -834 5074 -730
rect 5182 -834 5290 -730
rect 5398 -834 5506 -730
rect 5614 -834 5722 -730
rect 5830 -834 5938 -730
rect 6046 -834 6154 -730
rect 6262 -834 6370 -730
rect 6478 -834 6586 -730
rect 6694 -834 6712 -730
rect 3022 -836 6712 -834
rect 508 -852 6712 -836
rect 4500 -1260 4516 -1226
rect 4550 -1260 4566 -1226
rect 4728 -1260 4744 -1226
rect 4778 -1260 4794 -1226
rect 3328 -1942 4970 -1924
rect 3328 -1944 3474 -1942
rect 3328 -2002 3366 -1944
rect 3420 -2000 3474 -1944
rect 3528 -2000 3580 -1942
rect 3634 -2000 3688 -1942
rect 3742 -1944 4100 -1942
rect 3742 -2000 3798 -1944
rect 3420 -2002 3798 -2000
rect 3852 -2002 3900 -1944
rect 3954 -2002 4000 -1944
rect 4054 -2000 4100 -1944
rect 4154 -2000 4200 -1942
rect 4254 -1944 4500 -1942
rect 4254 -2000 4298 -1944
rect 4054 -2002 4298 -2000
rect 4352 -2002 4400 -1944
rect 4454 -2000 4500 -1944
rect 4554 -1944 4698 -1942
rect 4554 -2000 4600 -1944
rect 4454 -2002 4600 -2000
rect 4654 -2000 4698 -1944
rect 4752 -2000 4798 -1942
rect 4852 -2000 4898 -1942
rect 4952 -2000 4970 -1942
rect 4654 -2002 4970 -2000
rect 3328 -2022 4970 -2002
rect 4942 -2444 4958 -2410
rect 4992 -2444 5008 -2410
<< viali >>
rect 538 -836 646 -732
rect 754 -836 862 -732
rect 970 -836 1078 -732
rect 1186 -836 1294 -732
rect 1402 -836 1510 -732
rect 1618 -836 1726 -732
rect 1834 -836 1942 -732
rect 2050 -836 2158 -732
rect 2266 -836 2374 -732
rect 2482 -836 2590 -732
rect 2698 -836 2806 -732
rect 2914 -836 3022 -732
rect 3130 -834 3238 -730
rect 3346 -834 3454 -730
rect 3562 -834 3670 -730
rect 3778 -834 3886 -730
rect 3994 -834 4102 -730
rect 4210 -834 4318 -730
rect 4426 -834 4534 -730
rect 4642 -834 4750 -730
rect 4858 -834 4966 -730
rect 5074 -834 5182 -730
rect 5290 -834 5398 -730
rect 5506 -834 5614 -730
rect 5722 -834 5830 -730
rect 5938 -834 6046 -730
rect 6154 -834 6262 -730
rect 6370 -834 6478 -730
rect 6586 -834 6694 -730
rect 4516 -1260 4550 -1226
rect 4744 -1260 4778 -1226
rect 3366 -2002 3420 -1944
rect 3474 -2000 3528 -1942
rect 3580 -2000 3634 -1942
rect 3688 -2000 3742 -1942
rect 3798 -2002 3852 -1944
rect 3900 -2002 3954 -1944
rect 4000 -2002 4054 -1944
rect 4100 -2000 4154 -1942
rect 4200 -2000 4254 -1942
rect 4298 -2002 4352 -1944
rect 4400 -2002 4454 -1944
rect 4500 -2000 4554 -1942
rect 4600 -2002 4654 -1944
rect 4698 -2000 4752 -1942
rect 4798 -2000 4852 -1942
rect 4898 -2000 4952 -1942
rect 4958 -2444 4992 -2410
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 508 -710 708 -652
rect 508 -730 6716 -710
rect 508 -732 3130 -730
rect 508 -836 538 -732
rect 646 -836 754 -732
rect 862 -836 970 -732
rect 1078 -836 1186 -732
rect 1294 -836 1402 -732
rect 1510 -836 1618 -732
rect 1726 -836 1834 -732
rect 1942 -836 2050 -732
rect 2158 -836 2266 -732
rect 2374 -836 2482 -732
rect 2590 -836 2698 -732
rect 2806 -836 2914 -732
rect 3022 -834 3130 -732
rect 3238 -834 3346 -730
rect 3454 -834 3562 -730
rect 3670 -834 3778 -730
rect 3886 -834 3994 -730
rect 4102 -834 4210 -730
rect 4318 -834 4426 -730
rect 4534 -834 4642 -730
rect 4750 -834 4858 -730
rect 4966 -834 5074 -730
rect 5182 -834 5290 -730
rect 5398 -834 5506 -730
rect 5614 -834 5722 -730
rect 5830 -834 5938 -730
rect 6046 -834 6154 -730
rect 6262 -834 6370 -730
rect 6478 -834 6586 -730
rect 6694 -834 6716 -730
rect 3022 -836 6716 -834
rect 508 -852 6716 -836
rect 3452 -1222 3498 -1126
rect 4498 -1216 4566 -1210
rect 3452 -1268 3690 -1222
rect 0 -1600 200 -1400
rect 3452 -1654 3498 -1268
rect 3632 -1526 3690 -1268
rect 4498 -1268 4506 -1216
rect 4558 -1268 4566 -1216
rect 4498 -1278 4566 -1268
rect 4732 -1226 4790 -1220
rect 4732 -1260 4744 -1226
rect 4778 -1260 4790 -1226
rect 4732 -1410 4790 -1260
rect 4458 -1454 4790 -1410
rect 4458 -1670 4504 -1454
rect 4732 -1456 4790 -1454
rect 5364 -1272 5410 -1172
rect 5364 -1318 5650 -1272
rect 4760 -1494 4826 -1488
rect 4760 -1546 4768 -1494
rect 4820 -1546 4826 -1494
rect 4760 -1552 4826 -1546
rect 4766 -1656 4812 -1552
rect 5364 -1700 5410 -1318
rect 5592 -1576 5650 -1318
rect 0 -2000 200 -1800
rect 3326 -1942 4968 -1922
rect 3326 -1944 3474 -1942
rect 3326 -2002 3366 -1944
rect 3420 -2000 3474 -1944
rect 3528 -2000 3580 -1942
rect 3634 -2000 3688 -1942
rect 3742 -1944 4100 -1942
rect 3742 -2000 3798 -1944
rect 3420 -2002 3798 -2000
rect 3852 -2002 3900 -1944
rect 3954 -2002 4000 -1944
rect 4054 -2000 4100 -1944
rect 4154 -2000 4200 -1942
rect 4254 -1944 4500 -1942
rect 4254 -2000 4298 -1944
rect 4054 -2002 4298 -2000
rect 4352 -2002 4400 -1944
rect 4454 -2000 4500 -1944
rect 4554 -1944 4698 -1942
rect 4554 -2000 4600 -1944
rect 4454 -2002 4600 -2000
rect 4654 -2000 4698 -1944
rect 4752 -2000 4798 -1942
rect 4852 -2000 4898 -1942
rect 4952 -2000 4968 -1942
rect 4654 -2002 4968 -2000
rect 3326 -2020 4968 -2002
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 3450 -2611 3496 -2219
rect 4616 -2228 4764 -2156
rect 4612 -2302 4764 -2228
rect 3630 -2611 3688 -2353
rect 4612 -2410 4658 -2302
rect 4946 -2410 5004 -2404
rect 4612 -2444 4958 -2410
rect 4992 -2444 5006 -2410
rect 4612 -2446 5006 -2444
rect 3450 -2657 3688 -2611
rect 3450 -2747 3496 -2657
rect 4672 -2662 4712 -2446
rect 4946 -2450 5004 -2446
rect 4612 -2858 4770 -2662
rect 5550 -2700 5596 -2306
rect 5778 -2700 5836 -2442
rect 5550 -2746 5836 -2700
rect 5550 -2834 5596 -2746
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
<< via1 >>
rect 4506 -1226 4558 -1216
rect 4506 -1260 4516 -1226
rect 4516 -1260 4550 -1226
rect 4550 -1260 4558 -1226
rect 4506 -1268 4558 -1260
rect 4768 -1546 4820 -1494
<< rmetal2 >>
rect 4500 -1216 4564 -1210
rect 4500 -1268 4506 -1216
rect 4558 -1268 4564 -1216
rect 4500 -1502 4564 -1268
rect 4760 -1494 4826 -1488
rect 4760 -1502 4768 -1494
rect 4500 -1546 4768 -1502
rect 4820 -1546 4826 -1494
rect 4500 -1548 4826 -1546
rect 4760 -1552 4826 -1548
use sky130_fd_pr__nfet_01v8_PWNS5P  XM1
timestamp 1697007148
transform 1 0 2091 0 1 -2226
box -73 -430 73 488
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM2
timestamp 1697007148
transform 1 0 2789 0 1 -2162
box -221 -288 221 288
use sky130_fd_pr__nfet_01v8_lvt_F5PS5H  XM3
timestamp 1697007148
transform 1 0 1417 0 1 -2204
box -221 -288 221 288
use sky130_fd_pr__nfet_01v8_PWNS5P  XM4
timestamp 1697007148
transform 1 0 1837 0 1 -2194
box -73 -430 73 488
use sky130_fd_pr__nfet_01v8_PWNS5P  XM5
timestamp 1697007148
transform 1 0 2303 0 1 -2206
box -73 -430 73 488
use sky130_fd_pr__pfet_01v8_XGAKDL  XM6
timestamp 1697006309
transform 1 0 1845 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM7
timestamp 1697006309
transform 1 0 2257 0 1 -1197
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM8
timestamp 1697006309
transform 1 0 1429 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM9
timestamp 1697006309
transform 1 0 1229 0 1 -1195
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM10
timestamp 1697006309
transform 1 0 2677 0 1 -1197
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XGAKDL  XM11
timestamp 1697006309
transform 1 0 2879 0 1 -1197
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_MQX2PY  XM12
timestamp 1697008372
transform 1 0 3431 0 1 -1095
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1697008372
transform 1 0 3431 0 1 -1636
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM14
timestamp 1697012471
transform 1 0 3757 0 1 -1114
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM15
timestamp 1697012471
transform 1 0 3661 0 1 -1656
box -73 -138 73 188
use sky130_fd_pr__pfet_01v8_MQX2PY  XM16
timestamp 1697008372
transform 1 0 4533 0 1 -1095
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM17
timestamp 1697008372
transform 1 0 4761 0 1 -1095
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM18
timestamp 1697008372
transform 1 0 3429 0 -1 -2784
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM19
timestamp 1697022684
transform 1 0 4745 0 -1 -1712
box -73 -122 73 172
use sky130_fd_pr__nfet_01v8_L7T3GD  XM20
timestamp 1697008372
transform 1 0 3431 0 -1 -2207
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM21
timestamp 1697012471
transform 1 0 3755 0 -1 -2765
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM22
timestamp 1697012471
transform 1 0 3659 0 -1 -2221
box -73 -138 73 188
use sky130_fd_pr__nfet_01v8_9NW3WL  XM23
timestamp 1697022684
transform 1 0 4525 0 -1 -1712
box -73 -122 73 172
use sky130_fd_pr__pfet_01v8_MQX2PY  XM24
timestamp 1697008372
transform 1 0 4591 0 1 -2775
box -211 -303 211 303
use sky130_fd_pr__pfet_01v8_MQX2PY  XM25
timestamp 1697008372
transform 1 0 4791 0 1 -2775
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_9NW3WL  XM26
timestamp 1697022684
transform 1 0 4591 0 1 -2230
box -73 -122 73 172
use sky130_fd_pr__nfet_01v8_9NW3WL  XM27
timestamp 1697022684
transform 1 0 4791 0 1 -2230
box -73 -122 73 172
use sky130_fd_pr__pfet_01v8_MQX2PY  XM28
timestamp 1697008372
transform 1 0 4993 0 1 -2777
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM29
timestamp 1697008372
transform 1 0 4993 0 1 -2238
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_MQX2PY  XM30
timestamp 1697008372
transform 1 0 5339 0 1 -1147
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM31
timestamp 1697008372
transform 1 0 5339 0 1 -1698
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM32
timestamp 1697012471
transform 1 0 5717 0 1 -1164
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM33
timestamp 1697012471
transform 1 0 5623 0 1 -1708
box -73 -138 73 188
use sky130_fd_pr__pfet_01v8_MQX2PY  XM34
timestamp 1697008372
transform 1 0 5529 0 -1 -2869
box -211 -303 211 303
use sky130_fd_pr__nfet_01v8_L7T3GD  XM35
timestamp 1697008372
transform 1 0 5529 0 -1 -2276
box -73 -80 73 80
use sky130_fd_pr__pfet_01v8_HFBCFR  XM36
timestamp 1697012471
transform 1 0 5903 0 -1 -2854
box -311 -286 311 286
use sky130_fd_pr__nfet_01v8_648S5X  XM37
timestamp 1697012471
transform 1 0 5807 0 -1 -2312
box -73 -138 73 188
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 cdac_vn
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 cdac_vp
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 clk
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 X
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Y
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 P
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 Q
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 ready
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 X_drive
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 Y_drive
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 comp_outp
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 comp_outn
port 13 nsew
flabel metal1 508 -852 708 -652 0 FreeSans 256 0 0 0 VDD
port 3 nsew
<< end >>
