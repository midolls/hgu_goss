magic
tech sky130A
magscale 1 2
timestamp 1699322318
<< error_p >>
rect 39049 3126 39084 3160
rect 39050 3107 39084 3126
rect 38880 3058 38938 3064
rect 38880 3024 38892 3058
rect 38880 3018 38938 3024
rect 38880 2864 38938 2870
rect 38880 2830 38892 2864
rect 38880 2824 38938 2830
rect 39069 2728 39084 3107
rect 39103 3073 39138 3107
rect 39418 3073 39453 3107
rect 39103 2728 39137 3073
rect 39419 3054 39453 3073
rect 39249 3005 39307 3011
rect 39249 2971 39261 3005
rect 39249 2965 39307 2971
rect 39249 2811 39307 2817
rect 39249 2777 39261 2811
rect 39249 2771 39307 2777
rect 39103 2694 39118 2728
rect 39438 2675 39453 3054
rect 39472 3020 39507 3054
rect 39787 3020 39822 3054
rect 39472 2675 39506 3020
rect 39788 3001 39822 3020
rect 39618 2952 39676 2958
rect 39618 2918 39630 2952
rect 39618 2912 39676 2918
rect 39618 2758 39676 2764
rect 39618 2724 39630 2758
rect 39618 2718 39676 2724
rect 39472 2641 39487 2675
rect 39807 2622 39822 3001
rect 39841 2967 39876 3001
rect 40156 2967 40191 3001
rect 39841 2622 39875 2967
rect 40157 2948 40191 2967
rect 39987 2899 40045 2905
rect 39987 2865 39999 2899
rect 39987 2859 40045 2865
rect 39987 2705 40045 2711
rect 39987 2671 39999 2705
rect 39987 2665 40045 2671
rect 39841 2588 39856 2622
rect 40176 2569 40191 2948
rect 40210 2914 40245 2948
rect 40525 2914 40560 2948
rect 40210 2569 40244 2914
rect 40526 2895 40560 2914
rect 40356 2846 40414 2852
rect 40356 2812 40368 2846
rect 40356 2806 40414 2812
rect 40356 2652 40414 2658
rect 40356 2618 40368 2652
rect 40356 2612 40414 2618
rect 40210 2535 40225 2569
rect 40545 2516 40560 2895
rect 40579 2861 40614 2895
rect 40894 2861 40929 2895
rect 40579 2516 40613 2861
rect 40895 2842 40929 2861
rect 40725 2793 40783 2799
rect 40725 2759 40737 2793
rect 40725 2753 40783 2759
rect 40725 2599 40783 2605
rect 40725 2565 40737 2599
rect 40725 2559 40783 2565
rect 40579 2482 40594 2516
rect 40914 2463 40929 2842
rect 40948 2808 40983 2842
rect 41263 2808 41298 2842
rect 40948 2463 40982 2808
rect 41264 2789 41298 2808
rect 41094 2740 41152 2746
rect 41094 2706 41106 2740
rect 41094 2700 41152 2706
rect 41094 2546 41152 2552
rect 41094 2512 41106 2546
rect 41094 2506 41152 2512
rect 40948 2429 40963 2463
rect 41283 2410 41298 2789
rect 41317 2755 41352 2789
rect 41632 2755 41667 2789
rect 41317 2410 41351 2755
rect 41633 2736 41667 2755
rect 41463 2687 41521 2693
rect 41463 2653 41475 2687
rect 41463 2647 41521 2653
rect 41463 2493 41521 2499
rect 41463 2459 41475 2493
rect 41463 2453 41521 2459
rect 41317 2376 41332 2410
rect 41652 2357 41667 2736
rect 41686 2702 41721 2736
rect 42001 2702 42036 2736
rect 41686 2357 41720 2702
rect 42002 2683 42036 2702
rect 41832 2634 41890 2640
rect 41832 2600 41844 2634
rect 41832 2594 41890 2600
rect 41832 2440 41890 2446
rect 41832 2406 41844 2440
rect 41832 2400 41890 2406
rect 41686 2323 41701 2357
rect 42021 2304 42036 2683
rect 42055 2649 42090 2683
rect 42370 2649 42405 2683
rect 42055 2304 42089 2649
rect 42371 2630 42405 2649
rect 42201 2581 42259 2587
rect 42201 2547 42213 2581
rect 42201 2541 42259 2547
rect 42201 2387 42259 2393
rect 42201 2353 42213 2387
rect 42201 2347 42259 2353
rect 42055 2270 42070 2304
rect 42390 2251 42405 2630
rect 42424 2596 42459 2630
rect 42739 2596 42774 2630
rect 42424 2251 42458 2596
rect 42740 2577 42774 2596
rect 42570 2528 42628 2534
rect 42570 2494 42582 2528
rect 42570 2488 42628 2494
rect 42570 2334 42628 2340
rect 42570 2300 42582 2334
rect 42570 2294 42628 2300
rect 42424 2217 42439 2251
rect 42759 2198 42774 2577
rect 42793 2543 42828 2577
rect 43108 2543 43143 2577
rect 42793 2198 42827 2543
rect 43109 2524 43143 2543
rect 42939 2475 42997 2481
rect 42939 2441 42951 2475
rect 42939 2435 42997 2441
rect 42939 2281 42997 2287
rect 42939 2247 42951 2281
rect 42939 2241 42997 2247
rect 42793 2164 42808 2198
rect 43128 2145 43143 2524
rect 43162 2490 43197 2524
rect 43162 2145 43196 2490
rect 43308 2422 43366 2428
rect 43308 2388 43320 2422
rect 43308 2382 43366 2388
rect 43308 2228 43366 2234
rect 43308 2194 43320 2228
rect 43308 2188 43366 2194
rect 43162 2111 43177 2145
rect 6454 1040 6489 1074
rect 6454 1021 6488 1040
rect 6085 987 6120 1021
rect 6400 987 6435 1021
rect 6085 968 6119 987
rect 5716 934 5751 968
rect 6031 934 6066 968
rect 5716 915 5750 934
rect 5347 881 5382 915
rect 5662 881 5697 915
rect 5347 862 5381 881
rect 4978 828 5013 862
rect 5293 828 5328 862
rect 4978 809 5012 828
rect 4609 775 4644 809
rect 4924 775 4959 809
rect 4609 756 4643 775
rect 4555 722 4590 756
rect 4386 654 4444 660
rect 4432 620 4444 654
rect 4386 614 4444 620
rect 4386 460 4444 466
rect 4432 426 4444 460
rect 4386 420 4444 426
rect 4556 377 4590 722
rect 4609 377 4624 756
rect 4755 707 4813 713
rect 4801 673 4813 707
rect 4755 667 4813 673
rect 4755 513 4813 519
rect 4801 479 4813 513
rect 4755 473 4813 479
rect 4925 430 4959 775
rect 4978 430 4993 809
rect 5124 760 5182 766
rect 5170 726 5182 760
rect 5124 720 5182 726
rect 5124 566 5182 572
rect 5170 532 5182 566
rect 5124 526 5182 532
rect 5294 483 5328 828
rect 5347 483 5362 862
rect 5493 813 5551 819
rect 5539 779 5551 813
rect 5493 773 5551 779
rect 5493 619 5551 625
rect 5539 585 5551 619
rect 5493 579 5551 585
rect 5663 536 5697 881
rect 5716 536 5731 915
rect 5862 866 5920 872
rect 5908 832 5920 866
rect 5862 826 5920 832
rect 5862 672 5920 678
rect 5908 638 5920 672
rect 5862 632 5920 638
rect 6032 589 6066 934
rect 6085 589 6100 968
rect 6231 919 6289 925
rect 6277 885 6289 919
rect 6231 879 6289 885
rect 6231 725 6289 731
rect 6277 691 6289 725
rect 6231 685 6289 691
rect 6401 642 6435 987
rect 6454 642 6469 1021
rect 6420 608 6435 642
rect 6051 555 6066 589
rect 5682 502 5697 536
rect 5313 449 5328 483
rect 4944 396 4959 430
rect 4575 343 4590 377
<< error_s >>
rect 24526 4076 24584 4082
rect 25633 4076 25691 4082
rect 26740 4076 26798 4082
rect 27847 4076 27905 4082
rect 28954 4076 29012 4082
rect 30061 4076 30119 4082
rect 31168 4076 31226 4082
rect 32275 4076 32333 4082
rect 24526 4042 24538 4076
rect 25633 4042 25645 4076
rect 26740 4042 26752 4076
rect 27847 4042 27859 4076
rect 28954 4042 28966 4076
rect 30061 4042 30073 4076
rect 31168 4042 31180 4076
rect 32275 4042 32287 4076
rect 24526 4036 24584 4042
rect 25633 4036 25691 4042
rect 26740 4036 26798 4042
rect 27847 4036 27905 4042
rect 28954 4036 29012 4042
rect 30061 4036 30119 4042
rect 31168 4036 31226 4042
rect 32275 4036 32333 4042
rect 34790 4028 34848 4034
rect 34790 3994 34802 4028
rect 34790 3988 34848 3994
rect 23739 3331 23797 3337
rect 16081 3313 16139 3319
rect 17175 3313 17233 3319
rect 18269 3313 18327 3319
rect 19363 3313 19421 3319
rect 20457 3313 20515 3319
rect 21551 3313 21609 3319
rect 22645 3313 22703 3319
rect 16081 3279 16093 3313
rect 17175 3279 17187 3313
rect 18269 3279 18281 3313
rect 19363 3279 19375 3313
rect 20457 3279 20469 3313
rect 21551 3279 21563 3313
rect 22645 3279 22657 3313
rect 23739 3297 23751 3331
rect 23739 3291 23797 3297
rect 16081 3273 16139 3279
rect 17175 3273 17233 3279
rect 18269 3273 18327 3279
rect 19363 3273 19421 3279
rect 20457 3273 20515 3279
rect 21551 3273 21609 3279
rect 22645 3273 22703 3279
rect 16081 3119 16139 3125
rect 17175 3119 17233 3125
rect 18269 3119 18327 3125
rect 19363 3119 19421 3125
rect 20457 3119 20515 3125
rect 21551 3119 21609 3125
rect 22645 3119 22703 3125
rect 23739 3119 23797 3125
rect 16081 3085 16093 3119
rect 17175 3085 17187 3119
rect 18269 3085 18281 3119
rect 19363 3085 19375 3119
rect 20457 3085 20469 3119
rect 21551 3085 21563 3119
rect 22645 3085 22657 3119
rect 23739 3085 23751 3119
rect 16081 3079 16139 3085
rect 17175 3079 17233 3085
rect 18269 3079 18327 3085
rect 19363 3079 19421 3085
rect 20457 3079 20515 3085
rect 21551 3079 21609 3085
rect 22645 3079 22703 3085
rect 23739 3079 23797 3085
rect 15899 2947 15997 2986
rect 23980 2947 24233 3723
rect 24410 3469 24650 3723
rect 24664 3402 24904 3469
rect 24299 3363 24325 3395
rect 24664 2947 24906 3402
rect 25087 2947 25340 3723
rect 25517 3469 25757 3723
rect 25771 3402 26011 3469
rect 25406 3363 25432 3395
rect 25771 2947 26013 3402
rect 26194 2947 26447 3723
rect 26624 3469 26864 3723
rect 26878 3402 27118 3469
rect 26513 3363 26539 3395
rect 26878 2947 27120 3402
rect 27301 2947 27554 3723
rect 27731 3469 27971 3723
rect 27985 3402 28225 3469
rect 27620 3363 27646 3395
rect 27985 2947 28227 3402
rect 28408 2947 28661 3723
rect 28838 3469 29078 3723
rect 29092 3402 29332 3469
rect 28727 3363 28753 3395
rect 29092 2947 29334 3402
rect 29515 2947 29768 3723
rect 29945 3469 30185 3723
rect 30199 3402 30439 3469
rect 29834 3363 29860 3395
rect 30199 2947 30441 3402
rect 30622 2947 30875 3723
rect 31052 3469 31292 3723
rect 31306 3402 31546 3469
rect 30941 3363 30967 3395
rect 31306 2947 31548 3402
rect 31729 2947 31982 3723
rect 32048 3363 32074 3395
rect 34003 3283 34061 3289
rect 32909 3265 32967 3271
rect 32909 3231 32921 3265
rect 34003 3249 34015 3283
rect 34003 3243 34061 3249
rect 32909 3225 32967 3231
rect 32909 3071 32967 3077
rect 34003 3071 34061 3077
rect 32909 3037 32921 3071
rect 34003 3037 34015 3071
rect 32909 3031 32967 3037
rect 34003 3031 34061 3037
rect 10408 2902 10442 2916
rect 10488 2902 10522 2916
rect 11589 2902 11620 2919
rect 11666 2902 11700 2919
rect 11746 2902 11780 2919
rect 12112 2902 12146 2919
rect 12192 2902 12226 2919
rect 9808 2892 9933 2899
rect 9830 2865 9933 2892
rect 10408 2882 10569 2902
rect 10411 2868 10569 2882
rect 11623 2868 11781 2902
rect 12111 2868 12269 2902
rect 12272 2885 12303 2919
rect 12801 2902 12832 2919
rect 12878 2902 12912 2919
rect 12958 2902 12992 2919
rect 13324 2902 13358 2919
rect 13404 2902 13438 2919
rect 12835 2868 12993 2902
rect 13323 2868 13481 2902
rect 13484 2885 13515 2919
rect 14013 2902 14044 2919
rect 14090 2902 14124 2919
rect 14170 2902 14204 2919
rect 14536 2902 14570 2919
rect 14616 2902 14650 2919
rect 14047 2868 14205 2902
rect 14535 2868 14693 2902
rect 14696 2885 14727 2919
rect 15747 2868 15905 2902
rect 34244 2899 34497 3675
rect 34563 3315 34589 3347
rect 35638 3303 35673 3337
rect 35639 3284 35673 3303
rect 37942 3285 37977 3319
rect 35469 3235 35527 3241
rect 35469 3201 35481 3235
rect 35469 3195 35527 3201
rect 35437 3020 35465 3023
rect 35481 3016 35515 3023
rect 35531 3020 35559 3023
rect 35450 3004 35562 3016
rect 35443 2989 35562 3004
rect 35443 2975 35483 2989
rect 35425 2932 35483 2975
rect 35513 2975 35553 2989
rect 35513 2932 35571 2975
rect 35437 2928 35471 2932
rect 35525 2928 35559 2932
rect 35371 2907 35625 2921
rect 35287 2887 35625 2907
rect 35658 2887 35673 3284
rect 35692 3250 35727 3284
rect 36007 3250 36042 3284
rect 37943 3266 37977 3285
rect 35692 2887 35726 3250
rect 36008 3231 36042 3250
rect 35838 3182 35896 3188
rect 35838 3148 35850 3182
rect 35838 3142 35896 3148
rect 35838 2970 35896 2976
rect 35838 2936 35850 2970
rect 35838 2930 35896 2936
rect 9865 2816 9876 2865
rect 9899 2837 9933 2865
rect 15802 2838 15836 2868
rect 35287 2851 35388 2887
rect 35437 2878 35471 2882
rect 35525 2878 35559 2882
rect 35425 2862 35483 2878
rect 35513 2862 35571 2878
rect 35437 2853 35471 2862
rect 35525 2853 35559 2862
rect 35692 2853 35707 2887
rect 9899 2832 9964 2837
rect 15776 2834 15862 2838
rect 9899 2820 9933 2832
rect 9729 2797 9787 2803
rect 8198 2628 8233 2662
rect 8199 2609 8233 2628
rect 8029 2560 8087 2566
rect 8029 2526 8041 2560
rect 8029 2520 8087 2526
rect 8029 2348 8087 2354
rect 8029 2314 8041 2348
rect 8029 2308 8087 2314
rect 8218 2212 8233 2609
rect 8252 2575 8287 2609
rect 8567 2575 8602 2609
rect 8252 2212 8286 2575
rect 8568 2556 8602 2575
rect 8398 2507 8456 2513
rect 8398 2473 8410 2507
rect 8398 2467 8456 2473
rect 8398 2295 8456 2301
rect 8398 2261 8410 2295
rect 8398 2255 8456 2261
rect 8252 2178 8267 2212
rect 8587 2159 8602 2556
rect 8621 2522 8656 2556
rect 8936 2522 8971 2556
rect 8621 2159 8655 2522
rect 8937 2503 8971 2522
rect 8767 2454 8825 2460
rect 8767 2420 8779 2454
rect 8767 2414 8825 2420
rect 8767 2242 8825 2248
rect 8767 2208 8779 2242
rect 8767 2202 8825 2208
rect 8621 2125 8636 2159
rect 8956 2106 8971 2503
rect 8990 2469 9025 2503
rect 9305 2469 9340 2503
rect 9547 2486 9630 2793
rect 9729 2763 9741 2797
rect 9899 2794 9918 2820
rect 15772 2807 15862 2834
rect 10461 2800 10519 2806
rect 11673 2800 11731 2806
rect 12161 2800 12219 2806
rect 12885 2800 12943 2806
rect 13373 2800 13431 2806
rect 14097 2800 14155 2806
rect 14585 2800 14643 2806
rect 15797 2800 15855 2806
rect 9896 2780 9998 2794
rect 9729 2757 9787 2763
rect 9842 2744 9853 2754
rect 9836 2742 9853 2744
rect 9808 2716 9819 2720
rect 9808 2704 9825 2716
rect 9804 2682 9825 2704
rect 9836 2694 9857 2742
rect 9836 2682 9853 2694
rect 9776 2632 9831 2682
rect 9842 2678 9853 2682
rect 9865 2678 9876 2770
rect 9899 2766 9918 2780
rect 10461 2766 10473 2800
rect 11673 2766 11685 2800
rect 12161 2766 12173 2800
rect 12885 2766 12897 2800
rect 13373 2766 13385 2800
rect 14097 2766 14109 2800
rect 14585 2766 14597 2800
rect 15793 2766 15859 2800
rect 35656 2798 35862 2851
rect 36027 2834 36042 3231
rect 36061 3197 36096 3231
rect 36376 3197 36411 3231
rect 36061 2834 36095 3197
rect 36377 3178 36411 3197
rect 37773 3217 37831 3223
rect 37773 3183 37785 3217
rect 37962 3183 37977 3266
rect 36207 3129 36265 3135
rect 36207 3095 36219 3129
rect 36207 3089 36265 3095
rect 36207 2917 36265 2923
rect 36207 2883 36219 2917
rect 36207 2877 36265 2883
rect 36061 2800 36076 2834
rect 36396 2781 36411 3178
rect 36430 3144 36465 3178
rect 36745 3144 36780 3178
rect 37773 3177 37831 3183
rect 36430 2781 36464 3144
rect 36746 3125 36780 3144
rect 36576 3076 36634 3082
rect 36576 3042 36588 3076
rect 36576 3036 36634 3042
rect 36576 2864 36634 2870
rect 36576 2830 36588 2864
rect 36576 2824 36634 2830
rect 9899 2752 9970 2766
rect 10461 2760 10519 2766
rect 11673 2760 11731 2766
rect 12161 2760 12219 2766
rect 12885 2760 12943 2766
rect 13373 2760 13431 2766
rect 14097 2760 14155 2766
rect 14585 2760 14643 2766
rect 15797 2760 15855 2766
rect 9899 2682 9933 2752
rect 15781 2747 15867 2750
rect 36430 2747 36445 2781
rect 15777 2732 15867 2747
rect 15781 2719 15841 2732
rect 36765 2728 36780 3125
rect 36799 3091 36834 3125
rect 37114 3091 37149 3125
rect 36799 2728 36833 3091
rect 37115 3072 37149 3091
rect 37859 3073 37863 3144
rect 37867 3073 37869 3145
rect 36945 3023 37003 3029
rect 36945 2989 36957 3023
rect 36945 2983 37003 2989
rect 36945 2811 37003 2817
rect 36945 2777 36957 2811
rect 36945 2771 37003 2777
rect 15781 2707 15867 2719
rect 9808 2628 9819 2632
rect 9842 2628 9853 2632
rect 9836 2616 9853 2628
rect 9836 2606 9857 2616
rect 9836 2604 9853 2606
rect 9842 2594 9853 2604
rect 9729 2585 9787 2591
rect 9729 2551 9741 2585
rect 9729 2545 9787 2551
rect 9865 2540 9876 2632
rect 9899 2628 9918 2682
rect 15769 2664 15879 2707
rect 36799 2694 36814 2728
rect 37134 2675 37149 3072
rect 37168 3038 37203 3072
rect 37168 2675 37202 3038
rect 37859 3023 37877 3073
rect 37895 3033 37897 3145
rect 37909 3057 37935 3149
rect 37737 3007 37813 3023
rect 37817 3007 37877 3023
rect 37754 2995 37857 3007
rect 37747 2989 37857 2995
rect 37314 2970 37372 2976
rect 37747 2975 37787 2989
rect 37314 2936 37326 2970
rect 37314 2930 37372 2936
rect 37729 2923 37787 2975
rect 37817 2975 37835 2989
rect 37909 2975 37935 3011
rect 37943 2975 37977 3183
rect 37817 2923 37859 2975
rect 37889 2923 37977 2975
rect 37909 2921 37935 2923
rect 37943 2921 37977 2923
rect 37675 2887 37977 2921
rect 37996 3232 38031 3266
rect 38311 3232 38346 3266
rect 37996 2887 38030 3232
rect 38312 3213 38346 3232
rect 38142 3164 38200 3170
rect 38142 3130 38154 3164
rect 38142 3124 38200 3130
rect 38142 2970 38200 2976
rect 38142 2936 38154 2970
rect 38142 2930 38200 2936
rect 37741 2869 37775 2873
rect 37901 2869 37935 2873
rect 37729 2862 37787 2869
rect 37817 2862 37859 2869
rect 37889 2862 37947 2869
rect 37741 2853 37775 2862
rect 37901 2853 37935 2862
rect 37996 2853 38011 2887
rect 37996 2834 38001 2853
rect 38331 2834 38346 3213
rect 38365 3179 38400 3213
rect 38680 3179 38715 3213
rect 38365 2834 38399 3179
rect 38681 3160 38715 3179
rect 38511 3111 38569 3117
rect 38511 3077 38523 3111
rect 38511 3071 38569 3077
rect 38511 2917 38569 2923
rect 38511 2883 38523 2917
rect 38511 2877 38569 2883
rect 38365 2800 38380 2834
rect 38700 2781 38715 3160
rect 38734 3126 38769 3160
rect 38734 2781 38768 3126
rect 37314 2758 37372 2764
rect 37314 2724 37326 2758
rect 38734 2747 38749 2781
rect 37314 2718 37372 2724
rect 15769 2652 15799 2664
rect 15853 2652 15879 2664
rect 15753 2635 15793 2652
rect 15859 2635 15899 2652
rect 37168 2641 37183 2675
rect 15765 2631 15799 2632
rect 15853 2631 15887 2632
rect 9899 2544 9933 2628
rect 15809 2598 15876 2606
rect 10461 2588 10519 2594
rect 11673 2588 11731 2594
rect 12161 2588 12219 2594
rect 12885 2588 12943 2594
rect 13373 2588 13431 2594
rect 14097 2588 14155 2594
rect 14585 2588 14643 2594
rect 10461 2554 10473 2588
rect 11673 2554 11685 2588
rect 12161 2554 12173 2588
rect 12885 2554 12897 2588
rect 13373 2554 13385 2588
rect 14097 2554 14109 2588
rect 14585 2554 14597 2588
rect 15782 2587 15876 2598
rect 15793 2554 15876 2587
rect 10461 2548 10519 2554
rect 11673 2548 11731 2554
rect 12161 2548 12219 2554
rect 12885 2548 12943 2554
rect 13373 2548 13431 2554
rect 14097 2548 14155 2554
rect 14585 2548 14643 2554
rect 9865 2483 9876 2494
rect 9899 2490 9918 2544
rect 15793 2540 15859 2554
rect 9899 2483 9933 2490
rect 10289 2487 10315 2519
rect 11021 2490 11047 2522
rect 11633 2490 11659 2522
rect 12233 2490 12259 2522
rect 12845 2490 12871 2522
rect 13445 2490 13471 2522
rect 14057 2490 14083 2522
rect 14657 2490 14683 2522
rect 15269 2490 15295 2522
rect 15782 2512 15868 2540
rect 35431 2518 35477 2532
rect 37735 2509 37781 2532
rect 35403 2490 35505 2504
rect 9808 2478 9933 2483
rect 15748 2482 15902 2486
rect 8990 2106 9024 2469
rect 9306 2450 9340 2469
rect 9830 2451 9933 2478
rect 15728 2452 15922 2482
rect 37707 2481 37809 2504
rect 9136 2401 9194 2407
rect 9325 2406 9340 2450
rect 9136 2367 9148 2401
rect 9136 2361 9194 2367
rect 9306 2352 9340 2406
rect 9359 2416 9394 2450
rect 9679 2449 9976 2451
rect 9674 2416 9709 2449
rect 9359 2352 9393 2416
rect 9675 2397 9709 2416
rect 9830 2406 9888 2449
rect 9918 2406 9976 2449
rect 15782 2418 15868 2428
rect 9842 2402 9876 2406
rect 9930 2402 9964 2406
rect 9483 2352 9538 2382
rect 9694 2354 9709 2397
rect 9324 2321 9340 2352
rect 9344 2350 9394 2352
rect 9344 2321 9408 2350
rect 9479 2321 9589 2352
rect 9675 2350 9709 2354
rect 9650 2321 9709 2350
rect 9728 2363 9763 2397
rect 9776 2363 10030 2397
rect 9728 2352 9762 2363
rect 9842 2352 9876 2356
rect 9930 2352 9964 2356
rect 9728 2321 9743 2352
rect 9830 2338 9888 2352
rect 9918 2338 9976 2352
rect 9842 2329 9876 2338
rect 9344 2316 9709 2321
rect 9344 2312 9394 2316
rect 9407 2312 9661 2316
rect 9136 2189 9194 2195
rect 9136 2155 9148 2189
rect 9136 2149 9194 2155
rect 8990 2072 9005 2106
rect 9325 2053 9340 2287
rect 9359 2257 9393 2312
rect 9439 2293 9629 2305
rect 9435 2287 9633 2293
rect 9461 2257 9465 2267
rect 9359 2088 9394 2257
rect 9473 2245 9507 2271
rect 9460 2211 9507 2245
rect 9473 2195 9507 2211
rect 9561 2267 9595 2271
rect 9561 2257 9607 2267
rect 9561 2245 9595 2257
rect 9561 2211 9600 2245
rect 9561 2195 9595 2211
rect 9470 2178 9502 2183
rect 9457 2170 9502 2178
rect 9558 2170 9598 2183
rect 9457 2157 9598 2170
rect 9470 2137 9503 2157
rect 9558 2142 9598 2157
rect 9470 2136 9502 2137
rect 9501 2088 9502 2136
rect 9505 2129 9598 2142
rect 9505 2109 9551 2129
rect 9517 2106 9551 2109
rect 9528 2102 9551 2106
rect 9558 2102 9598 2129
rect 9359 2057 9420 2088
rect 9450 2068 9502 2088
rect 9444 2057 9502 2068
rect 9558 2089 9589 2102
rect 9558 2088 9567 2089
rect 9675 2088 9709 2316
rect 9558 2068 9610 2088
rect 9558 2057 9616 2068
rect 9640 2057 9709 2088
rect 9359 2053 9393 2057
rect 9359 2047 9374 2053
rect 9694 2047 9709 2057
rect 9359 2034 9393 2047
rect 9675 2034 9709 2047
rect 9359 2032 9502 2034
rect 9558 2032 9709 2034
rect 9359 2023 9464 2032
rect 9596 2023 9709 2032
rect 9359 2011 9452 2023
rect 9608 2011 9709 2023
rect 9359 2005 9461 2011
rect 9599 2005 9709 2011
rect 9728 2005 9762 2312
rect 9848 2311 9876 2329
rect 9920 2311 9967 2338
rect 9848 2298 9888 2311
rect 9918 2298 9967 2311
rect 9848 2280 9967 2298
rect 9855 2268 9967 2280
rect 9886 2261 9920 2268
rect 9323 1981 9762 2005
rect 9780 1981 9796 2025
rect 9323 1964 9760 1981
rect 9692 1911 9760 1964
rect 9784 1954 9901 1966
rect 9784 1947 10062 1954
rect 9818 1920 9867 1932
rect 9818 1913 10028 1920
rect 15513 1772 15547 1990
rect 15655 1950 15721 1982
rect 15561 1914 15815 1948
rect 15627 1903 15661 1907
rect 15715 1903 15749 1907
rect 15615 1889 15673 1903
rect 15703 1889 15761 1903
rect 15627 1880 15661 1889
rect 15633 1862 15661 1880
rect 15705 1862 15752 1889
rect 15633 1849 15673 1862
rect 15703 1849 15752 1862
rect 15633 1831 15752 1849
rect 15640 1819 15752 1831
rect 15655 1812 15721 1819
rect 15655 1796 15673 1812
rect 15703 1796 15721 1812
rect 15829 1787 15863 1990
rect 15829 1772 15879 1787
rect 9775 1517 9810 1551
rect 9406 1464 9441 1498
rect 9037 1411 9072 1445
rect 8668 1358 8703 1392
rect 8299 1305 8334 1339
rect 7930 1252 7965 1286
rect 7561 1199 7596 1233
rect 7192 1146 7227 1180
rect 6823 1093 6858 1127
rect 6600 972 6658 978
rect 6600 938 6612 972
rect 6600 932 6658 938
rect 6600 778 6658 784
rect 6600 744 6612 778
rect 6600 738 6658 744
rect 6789 661 6804 1074
rect 6823 729 6857 1093
rect 6969 1025 7027 1031
rect 6969 991 6981 1025
rect 6969 985 7027 991
rect 6969 831 7027 837
rect 6969 797 6981 831
rect 6969 791 7027 797
rect 6823 695 6858 729
rect 7158 714 7173 1127
rect 7192 782 7226 1146
rect 7338 1078 7396 1084
rect 7338 1044 7350 1078
rect 7338 1038 7396 1044
rect 7338 884 7396 890
rect 7338 850 7350 884
rect 7338 844 7396 850
rect 7192 748 7227 782
rect 7527 767 7542 1180
rect 7561 835 7595 1199
rect 7707 1131 7765 1137
rect 7707 1097 7719 1131
rect 7707 1091 7765 1097
rect 7707 937 7765 943
rect 7707 903 7719 937
rect 7707 897 7765 903
rect 7561 801 7596 835
rect 7896 820 7911 1233
rect 7930 888 7964 1252
rect 8076 1184 8134 1190
rect 8076 1150 8088 1184
rect 8076 1144 8134 1150
rect 8076 990 8134 996
rect 8076 956 8088 990
rect 8076 950 8134 956
rect 7930 854 7965 888
rect 8265 873 8280 1286
rect 8299 941 8333 1305
rect 8445 1237 8503 1243
rect 8445 1203 8457 1237
rect 8445 1197 8503 1203
rect 8445 1043 8503 1049
rect 8445 1009 8457 1043
rect 8445 1003 8503 1009
rect 8299 907 8334 941
rect 8634 926 8649 1339
rect 8668 994 8702 1358
rect 8814 1290 8872 1296
rect 8814 1256 8826 1290
rect 8814 1250 8872 1256
rect 8814 1096 8872 1102
rect 8814 1062 8826 1096
rect 8814 1056 8872 1062
rect 8668 960 8703 994
rect 9003 979 9018 1392
rect 9037 1047 9071 1411
rect 9183 1343 9241 1349
rect 9183 1309 9195 1343
rect 9183 1303 9241 1309
rect 9183 1149 9241 1155
rect 9183 1115 9195 1149
rect 9183 1109 9241 1115
rect 9037 1013 9072 1047
rect 9372 1032 9387 1445
rect 9406 1100 9440 1464
rect 9552 1202 9610 1208
rect 9552 1168 9564 1202
rect 9552 1162 9610 1168
rect 9406 1066 9441 1100
rect 9741 1085 9756 1498
rect 9775 1377 9809 1517
rect 9953 1449 9979 1455
rect 9897 1415 9931 1449
rect 9933 1415 9979 1449
rect 9953 1409 9979 1415
rect 9981 1381 10007 1483
rect 15477 1462 15899 1772
rect 15924 1681 15947 1822
rect 15952 1653 15975 1800
rect 15924 1594 15933 1640
rect 15952 1600 15961 1653
rect 9775 1293 9810 1377
rect 9775 1239 9809 1293
rect 9817 1289 9843 1381
rect 9855 1265 9857 1377
rect 9883 1376 9885 1377
rect 9878 1365 9893 1376
rect 9883 1305 9885 1365
rect 9889 1305 9893 1365
rect 9875 1271 9893 1305
rect 9917 1255 9935 1271
rect 15513 1262 15547 1462
rect 15659 1456 15709 1462
rect 15659 1440 15709 1446
rect 15623 1424 15753 1440
rect 15640 1412 15743 1424
rect 15633 1406 15743 1412
rect 15633 1392 15673 1406
rect 15615 1340 15673 1392
rect 15703 1392 15743 1406
rect 15703 1340 15761 1392
rect 15615 1315 15761 1338
rect 15621 1304 15755 1315
rect 15655 1270 15721 1302
rect 15829 1262 15863 1462
rect 9775 1207 9810 1239
rect 9817 1207 9843 1243
rect 9893 1239 9935 1255
rect 9939 1239 10015 1255
rect 9902 1224 10005 1239
rect 9917 1221 10005 1224
rect 9917 1207 9935 1221
rect 9775 1155 9863 1207
rect 9893 1155 9935 1207
rect 9965 1207 10005 1221
rect 9965 1155 10023 1207
rect 9775 1153 9809 1155
rect 9817 1153 9843 1155
rect 9775 1119 10077 1153
rect 9817 1101 9851 1105
rect 9977 1101 10011 1105
rect 9805 1094 9863 1101
rect 9893 1094 9935 1101
rect 9965 1094 10023 1101
rect 9805 1066 9810 1094
rect 9817 1085 9851 1094
rect 9977 1085 10011 1094
rect 9971 741 10017 764
rect 9943 713 10045 736
<< nwell >>
rect 9791 2389 15997 2986
rect 9742 2388 15997 2389
rect 9262 2322 15997 2388
rect 9262 2300 9760 2322
rect 9264 2298 9760 2300
rect 9453 2146 9501 2202
rect 9791 1692 15997 2322
<< ndiff >>
rect 11664 1549 11722 1561
rect 11664 1489 11676 1549
rect 11710 1489 11722 1549
rect 11664 1477 11722 1489
rect 12875 1549 12933 1561
rect 12875 1489 12887 1549
rect 12921 1489 12933 1549
rect 12875 1477 12933 1489
rect 14215 1549 14273 1561
rect 14215 1489 14227 1549
rect 14261 1489 14273 1549
rect 14215 1477 14273 1489
rect 14962 1549 15020 1561
rect 14962 1489 14974 1549
rect 15008 1489 15020 1549
rect 14962 1477 15020 1489
<< pdiff >>
rect 9453 2146 9501 2202
rect 11309 1750 11367 1762
rect 11309 1690 11321 1750
rect 11355 1690 11367 1750
rect 11309 1678 11367 1690
rect 12520 1750 12578 1762
rect 12520 1690 12532 1750
rect 12566 1690 12578 1750
rect 12520 1678 12578 1690
rect 13733 1750 13791 1762
rect 13733 1690 13745 1750
rect 13779 1690 13791 1750
rect 13733 1678 13791 1690
rect 14947 1750 15005 1762
rect 14947 1690 14959 1750
rect 14993 1690 15005 1750
rect 14947 1678 15005 1690
<< ndiffc >>
rect 10927 1489 10961 1549
rect 11676 1489 11710 1549
rect 12887 1489 12921 1549
rect 14227 1489 14261 1549
rect 14974 1489 15008 1549
<< pdiffc >>
rect 10572 1690 10606 1750
rect 11321 1690 11355 1750
rect 12532 1690 12566 1750
rect 13745 1690 13779 1750
rect 14959 1690 14993 1750
<< psubdiff >>
rect 9370 1714 9394 1748
rect 9428 1714 9512 1748
rect 9546 1714 9656 1748
rect 9690 1714 9732 1748
rect 9370 1712 9732 1714
<< nsubdiff >>
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9344 2350 9760 2352
rect 9344 2316 9374 2350
rect 9408 2316 9504 2350
rect 9538 2316 9650 2350
rect 9684 2316 9760 2350
rect 15782 2342 15868 2368
rect 9344 2312 9760 2316
rect 15781 2245 15867 2271
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 15781 2185 15867 2211
<< psubdiffcont >>
rect 9394 1714 9428 1748
rect 9512 1714 9546 1748
rect 9656 1714 9690 1748
<< nsubdiffcont >>
rect 15802 2834 15836 2868
rect 15807 2690 15841 2724
rect 15808 2538 15842 2572
rect 15808 2368 15842 2402
rect 9374 2316 9408 2350
rect 9504 2316 9538 2350
rect 9650 2316 9684 2350
rect 15807 2211 15841 2245
<< poly >>
rect 15544 1636 15703 1656
rect 15544 1602 15556 1636
rect 15590 1602 15703 1636
rect 15544 1583 15703 1602
rect 15765 1577 15891 1656
rect 9881 1449 9947 1465
rect 9881 1422 9897 1449
rect 9863 1415 9897 1422
rect 9931 1422 9947 1449
rect 9931 1415 9965 1422
rect 9863 1392 9965 1415
<< polycont >>
rect 15556 1602 15590 1636
rect 9897 1415 9931 1449
<< locali >>
rect 9938 2868 10053 2908
rect 15776 2868 15862 2894
rect 15776 2834 15802 2868
rect 15836 2834 15862 2868
rect 15776 2808 15862 2834
rect 15781 2724 15867 2750
rect 15781 2690 15807 2724
rect 15841 2690 15867 2724
rect 15781 2664 15867 2690
rect 15782 2572 15868 2598
rect 15782 2538 15808 2572
rect 15842 2538 15868 2572
rect 15782 2512 15868 2538
rect 15782 2402 15868 2428
rect 15782 2368 15808 2402
rect 15842 2368 15868 2402
rect 9358 2316 9374 2350
rect 9408 2316 9424 2350
rect 9488 2316 9504 2350
rect 9538 2316 9558 2350
rect 9634 2318 9650 2350
rect 9684 2318 9704 2350
rect 15782 2342 15868 2368
rect 15781 2245 15867 2271
rect 15781 2211 15807 2245
rect 15841 2211 15867 2245
rect 9453 2178 9501 2202
rect 15781 2185 15867 2211
rect 9453 2146 9457 2178
rect 9491 2146 9501 2178
rect 9647 2012 9681 2021
rect 9780 2013 9829 2025
rect 9647 1987 9650 2012
rect 9780 1979 9789 2013
rect 9823 2008 9829 2013
rect 9823 1979 10112 2008
rect 9780 1973 10112 1979
rect 9780 1966 9829 1973
rect 10077 1950 10112 1973
rect 10077 1938 10126 1950
rect 9818 1920 9867 1932
rect 9818 1886 9827 1920
rect 9861 1886 10028 1920
rect 10077 1904 10086 1938
rect 10120 1904 10126 1938
rect 10077 1891 10126 1904
rect 9818 1873 9867 1886
rect 9987 1844 10028 1886
rect 10078 1845 10127 1857
rect 10078 1844 10087 1845
rect 9987 1811 10087 1844
rect 10121 1811 10127 1845
rect 9987 1810 10127 1811
rect 10078 1798 10127 1810
rect 9378 1748 9454 1756
rect 9378 1714 9394 1748
rect 9428 1714 9454 1748
rect 9496 1748 9572 1756
rect 10572 1750 10606 1766
rect 9496 1714 9512 1748
rect 9546 1714 9572 1748
rect 9638 1714 9656 1744
rect 9690 1714 9706 1744
rect 10572 1674 10606 1690
rect 11321 1750 11355 1766
rect 11321 1674 11355 1690
rect 12532 1750 12566 1766
rect 12532 1674 12566 1690
rect 13745 1750 13779 1766
rect 13745 1674 13779 1690
rect 14959 1750 14993 1766
rect 14959 1674 14993 1690
rect 15540 1602 15556 1636
rect 15590 1602 15606 1636
rect 10927 1549 10961 1565
rect 10927 1473 10961 1489
rect 11676 1549 11710 1565
rect 11676 1473 11710 1489
rect 12887 1549 12921 1565
rect 12887 1473 12921 1489
rect 14227 1549 14261 1565
rect 14227 1473 14261 1489
rect 14974 1549 15008 1565
rect 14974 1473 15008 1489
rect 9881 1415 9897 1449
rect 9931 1415 9947 1449
<< viali >>
rect 15802 2834 15836 2868
rect 15807 2690 15841 2724
rect 15808 2538 15842 2572
rect 15808 2368 15842 2402
rect 15807 2211 15841 2245
rect 9457 2144 9491 2178
rect 9566 2089 9600 2123
rect 9376 1979 9410 2013
rect 9650 1978 9684 2012
rect 9789 1979 9823 2013
rect 9827 1886 9861 1920
rect 10086 1904 10120 1938
rect 10087 1811 10121 1845
rect 10572 1690 10606 1750
rect 11321 1690 11355 1750
rect 12532 1690 12566 1750
rect 13745 1690 13779 1750
rect 14959 1690 14993 1750
rect 15556 1602 15590 1636
rect 10927 1489 10961 1549
rect 11676 1489 11710 1549
rect 12887 1489 12921 1549
rect 14227 1489 14261 1549
rect 14974 1489 15008 1549
rect 9897 1415 9931 1449
<< metal1 >>
rect 9963 2937 10053 2953
rect 9963 2926 9982 2937
rect 9945 2885 9982 2926
rect 10034 2885 10053 2937
rect 9945 2870 10053 2885
rect 15772 2875 15862 2891
rect 9945 2838 9998 2870
rect 15772 2823 15791 2875
rect 15843 2823 15862 2875
rect 15772 2807 15862 2823
rect 15777 2731 15867 2747
rect 15777 2679 15796 2731
rect 15848 2679 15867 2731
rect 15777 2663 15867 2679
rect 15778 2579 15868 2595
rect 15778 2527 15797 2579
rect 15849 2527 15868 2579
rect 15778 2511 15868 2527
rect 15778 2409 15868 2425
rect 15778 2357 15797 2409
rect 15849 2357 15868 2409
rect 9358 2332 9424 2350
rect 9358 2316 9365 2332
rect 9363 2280 9365 2316
rect 9417 2316 9424 2332
rect 9494 2331 9550 2342
rect 9417 2280 9419 2316
rect 9363 2269 9419 2280
rect 9494 2279 9496 2331
rect 9548 2279 9550 2331
rect 9634 2332 9704 2350
rect 15778 2341 15868 2357
rect 9634 2318 9640 2332
rect 9494 2268 9550 2279
rect 9638 2280 9640 2318
rect 9692 2318 9704 2332
rect 9692 2280 9694 2318
rect 9638 2269 9694 2280
rect 15777 2252 15867 2268
rect 9445 2178 9808 2185
rect 9445 2144 9457 2178
rect 9491 2157 9808 2178
rect 9491 2144 9503 2157
rect 9445 2137 9503 2144
rect 9550 2123 9617 2129
rect 9550 2089 9566 2123
rect 9600 2110 9617 2123
rect 9600 2089 9752 2110
rect 9550 2082 9752 2089
rect 9630 2021 9696 2023
rect 9368 2016 9422 2020
rect 9367 2013 9422 2016
rect 9238 1979 9376 2013
rect 9410 1979 9422 2013
rect 9367 1976 9422 1979
rect 9367 1972 9421 1976
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 9724 1938 9752 2082
rect 9780 2025 9808 2157
rect 9956 2130 10027 2214
rect 15777 2200 15796 2252
rect 15848 2200 15867 2252
rect 15777 2184 15867 2200
rect 9780 2013 9829 2025
rect 9780 1979 9789 2013
rect 9823 1979 9829 2013
rect 9780 1966 9829 1979
rect 9724 1920 9867 1938
rect 9724 1910 9827 1920
rect 9818 1886 9827 1910
rect 9861 1886 9867 1920
rect 9818 1873 9867 1886
rect 9381 1786 9437 1797
rect 9381 1756 9383 1786
rect 9378 1734 9383 1756
rect 9435 1756 9437 1786
rect 9501 1786 9557 1797
rect 9501 1756 9503 1786
rect 9435 1734 9454 1756
rect 9378 1714 9454 1734
rect 9496 1734 9503 1756
rect 9555 1756 9557 1786
rect 9644 1786 9700 1797
rect 9555 1734 9572 1756
rect 9644 1744 9646 1786
rect 9496 1714 9572 1734
rect 9638 1734 9646 1744
rect 9698 1744 9700 1786
rect 9698 1734 9706 1744
rect 9638 1714 9706 1734
rect 9895 1643 9943 2089
rect 9275 1596 9943 1643
rect 9895 1455 9943 1596
rect 9885 1449 9943 1455
rect 9644 1443 9709 1444
rect 9644 1442 9650 1443
rect 9548 1440 9650 1442
rect 9546 1394 9650 1440
rect 9644 1391 9650 1394
rect 9702 1391 9709 1443
rect 9885 1415 9897 1449
rect 9931 1415 9943 1449
rect 9885 1409 9943 1415
rect 9981 1640 10027 2130
rect 15695 2010 15785 2026
rect 15695 1999 15714 2010
rect 15620 1958 15714 1999
rect 15766 1958 15785 2010
rect 10077 1943 10126 1950
rect 10077 1938 10696 1943
rect 10077 1904 10086 1938
rect 10120 1904 10696 1938
rect 10077 1896 10696 1904
rect 10077 1891 10126 1896
rect 10078 1849 10127 1857
rect 10647 1849 10696 1896
rect 15620 1940 15785 1958
rect 15620 1894 15667 1940
rect 10078 1845 10579 1849
rect 10078 1811 10087 1845
rect 10121 1811 10579 1845
rect 10078 1803 10579 1811
rect 10647 1803 15068 1849
rect 10078 1802 10567 1803
rect 10647 1802 11093 1803
rect 10078 1798 10127 1802
rect 15709 1793 15947 1822
rect 10566 1750 10612 1762
rect 10566 1690 10572 1750
rect 10606 1690 10612 1750
rect 10566 1640 10612 1690
rect 11315 1750 11361 1762
rect 11315 1690 11321 1750
rect 11355 1690 11361 1750
rect 11315 1640 11361 1690
rect 12526 1750 12572 1762
rect 12526 1690 12532 1750
rect 12566 1690 12572 1750
rect 12526 1640 12572 1690
rect 13739 1750 13785 1762
rect 13739 1690 13745 1750
rect 13779 1690 13785 1750
rect 13739 1640 13785 1690
rect 14953 1750 14999 1762
rect 15709 1756 15755 1793
rect 14953 1690 14959 1750
rect 14993 1690 14999 1750
rect 14953 1640 14999 1690
rect 15783 1749 15873 1765
rect 15901 1764 15947 1793
rect 15783 1697 15802 1749
rect 15854 1697 15873 1749
rect 15540 1640 15606 1642
rect 9981 1636 15606 1640
rect 9981 1602 15556 1636
rect 15590 1602 15606 1636
rect 9981 1598 15606 1602
rect 9981 1368 10027 1598
rect 10921 1549 10967 1598
rect 10921 1489 10927 1549
rect 10961 1489 10967 1549
rect 10921 1477 10967 1489
rect 11670 1549 11716 1598
rect 11670 1489 11676 1549
rect 11710 1489 11716 1549
rect 11670 1477 11716 1489
rect 12881 1549 12927 1598
rect 12881 1489 12887 1549
rect 12921 1489 12927 1549
rect 12881 1477 12927 1489
rect 14221 1549 14267 1598
rect 14221 1489 14227 1549
rect 14261 1489 14267 1549
rect 14221 1477 14267 1489
rect 14968 1549 15014 1598
rect 15544 1596 15606 1598
rect 15639 1633 15667 1683
rect 15783 1681 15873 1697
rect 15751 1633 15933 1640
rect 15639 1604 15933 1633
rect 15639 1556 15667 1604
rect 15751 1594 15933 1604
rect 14968 1489 14974 1549
rect 15008 1489 15014 1549
rect 14968 1477 15014 1489
rect 15783 1546 15873 1562
rect 15783 1494 15802 1546
rect 15854 1494 15873 1546
rect 15709 1450 15755 1480
rect 15783 1478 15873 1494
rect 15901 1450 15947 1481
rect 10131 1391 10138 1443
rect 10190 1441 10196 1443
rect 10190 1424 10913 1441
rect 10190 1394 10929 1424
rect 11603 1399 12997 1445
rect 14153 1399 14335 1445
rect 10190 1391 10196 1394
rect 10131 1390 10196 1391
rect 10871 1389 10929 1394
rect 10013 1293 10027 1368
rect 9932 359 10039 375
rect 9932 307 9968 359
rect 10020 307 10039 359
rect 9932 291 10039 307
rect 11727 268 11785 1399
rect 14153 268 14211 1399
rect 15009 267 15068 1448
rect 15709 1421 15947 1450
rect 15621 1300 15667 1344
rect 15621 1284 15782 1300
rect 15621 1232 15711 1284
rect 15763 1232 15782 1284
rect 15621 1216 15782 1232
<< via1 >>
rect 9982 2885 10034 2937
rect 15791 2868 15843 2875
rect 15791 2834 15802 2868
rect 15802 2834 15836 2868
rect 15836 2834 15843 2868
rect 15791 2823 15843 2834
rect 15796 2724 15848 2731
rect 15796 2690 15807 2724
rect 15807 2690 15841 2724
rect 15841 2690 15848 2724
rect 15796 2679 15848 2690
rect 15797 2572 15849 2579
rect 15797 2538 15808 2572
rect 15808 2538 15842 2572
rect 15842 2538 15849 2572
rect 15797 2527 15849 2538
rect 15797 2402 15849 2409
rect 15797 2368 15808 2402
rect 15808 2368 15842 2402
rect 15842 2368 15849 2402
rect 15797 2357 15849 2368
rect 9365 2280 9417 2332
rect 9496 2279 9548 2331
rect 9640 2280 9692 2332
rect 9638 2012 9690 2021
rect 9638 1978 9650 2012
rect 9650 1978 9684 2012
rect 9684 1978 9690 2012
rect 9638 1969 9690 1978
rect 15796 2245 15848 2252
rect 15796 2211 15807 2245
rect 15807 2211 15841 2245
rect 15841 2211 15848 2245
rect 15796 2200 15848 2211
rect 9383 1734 9435 1786
rect 9503 1734 9555 1786
rect 9646 1734 9698 1786
rect 9650 1391 9702 1443
rect 15714 1958 15766 2010
rect 15802 1697 15854 1749
rect 15802 1494 15854 1546
rect 10138 1391 10190 1443
rect 9968 307 10020 359
rect 15711 1232 15763 1284
<< metal2 >>
rect 9971 2939 10045 2943
rect 9971 2883 9980 2939
rect 10036 2883 10045 2939
rect 9971 2879 10045 2883
rect 15780 2877 15854 2881
rect 15780 2821 15789 2877
rect 15845 2821 15854 2877
rect 15780 2817 15854 2821
rect 15785 2733 15859 2737
rect 15785 2677 15794 2733
rect 15850 2677 15859 2733
rect 15785 2673 15859 2677
rect 15786 2581 15860 2585
rect 15786 2525 15795 2581
rect 15851 2525 15860 2581
rect 15786 2521 15860 2525
rect 15786 2411 15860 2415
rect 15786 2355 15795 2411
rect 15851 2355 15860 2411
rect 15786 2351 15860 2355
rect 9363 2334 9419 2343
rect 9363 2269 9419 2278
rect 9494 2333 9550 2342
rect 9494 2268 9550 2277
rect 9638 2334 9694 2343
rect 9638 2269 9694 2278
rect 15785 2254 15859 2258
rect 15785 2198 15794 2254
rect 15850 2198 15859 2254
rect 15785 2194 15859 2198
rect 9630 1969 9638 2021
rect 9690 1969 9696 2021
rect 9630 1968 9696 1969
rect 15703 2012 15777 2016
rect 9648 1892 9694 1968
rect 15703 1956 15712 2012
rect 15768 1956 15777 2012
rect 15703 1952 15777 1956
rect 9648 1846 9887 1892
rect 9381 1788 9437 1797
rect 9381 1723 9437 1732
rect 9501 1788 9557 1797
rect 9501 1723 9557 1732
rect 9644 1788 9700 1797
rect 9644 1723 9700 1732
rect 9644 1443 9709 1444
rect 9644 1391 9650 1443
rect 9702 1440 9709 1443
rect 9841 1440 9887 1846
rect 15791 1751 15865 1755
rect 15791 1695 15800 1751
rect 15856 1695 15865 1751
rect 15791 1691 15865 1695
rect 15791 1548 15865 1552
rect 15791 1492 15800 1548
rect 15856 1492 15865 1548
rect 15791 1488 15865 1492
rect 10131 1440 10138 1443
rect 9702 1394 10138 1440
rect 9702 1391 9709 1394
rect 10131 1391 10138 1394
rect 10190 1391 10196 1443
rect 10131 1390 10196 1391
rect 15700 1286 15774 1290
rect 15700 1230 15709 1286
rect 15765 1230 15774 1286
rect 15700 1226 15774 1230
rect 9957 361 10031 365
rect 9957 305 9966 361
rect 10022 305 10031 361
rect 9957 301 10031 305
<< via2 >>
rect 9980 2937 10036 2939
rect 9980 2885 9982 2937
rect 9982 2885 10034 2937
rect 10034 2885 10036 2937
rect 9980 2883 10036 2885
rect 15789 2875 15845 2877
rect 15789 2823 15791 2875
rect 15791 2823 15843 2875
rect 15843 2823 15845 2875
rect 15789 2821 15845 2823
rect 15794 2731 15850 2733
rect 15794 2679 15796 2731
rect 15796 2679 15848 2731
rect 15848 2679 15850 2731
rect 15794 2677 15850 2679
rect 15795 2579 15851 2581
rect 15795 2527 15797 2579
rect 15797 2527 15849 2579
rect 15849 2527 15851 2579
rect 15795 2525 15851 2527
rect 15795 2409 15851 2411
rect 15795 2357 15797 2409
rect 15797 2357 15849 2409
rect 15849 2357 15851 2409
rect 15795 2355 15851 2357
rect 9363 2332 9419 2334
rect 9363 2280 9365 2332
rect 9365 2280 9417 2332
rect 9417 2280 9419 2332
rect 9363 2278 9419 2280
rect 9494 2331 9550 2333
rect 9494 2279 9496 2331
rect 9496 2279 9548 2331
rect 9548 2279 9550 2331
rect 9494 2277 9550 2279
rect 9638 2332 9694 2334
rect 9638 2280 9640 2332
rect 9640 2280 9692 2332
rect 9692 2280 9694 2332
rect 9638 2278 9694 2280
rect 15794 2252 15850 2254
rect 15794 2200 15796 2252
rect 15796 2200 15848 2252
rect 15848 2200 15850 2252
rect 15794 2198 15850 2200
rect 15712 2010 15768 2012
rect 15712 1958 15714 2010
rect 15714 1958 15766 2010
rect 15766 1958 15768 2010
rect 15712 1956 15768 1958
rect 9381 1786 9437 1788
rect 9381 1734 9383 1786
rect 9383 1734 9435 1786
rect 9435 1734 9437 1786
rect 9381 1732 9437 1734
rect 9501 1786 9557 1788
rect 9501 1734 9503 1786
rect 9503 1734 9555 1786
rect 9555 1734 9557 1786
rect 9501 1732 9557 1734
rect 9644 1786 9700 1788
rect 9644 1734 9646 1786
rect 9646 1734 9698 1786
rect 9698 1734 9700 1786
rect 9644 1732 9700 1734
rect 15800 1749 15856 1751
rect 15800 1697 15802 1749
rect 15802 1697 15854 1749
rect 15854 1697 15856 1749
rect 15800 1695 15856 1697
rect 15800 1546 15856 1548
rect 15800 1494 15802 1546
rect 15802 1494 15854 1546
rect 15854 1494 15856 1546
rect 15800 1492 15856 1494
rect 15709 1284 15765 1286
rect 15709 1232 15711 1284
rect 15711 1232 15763 1284
rect 15763 1232 15765 1284
rect 15709 1230 15765 1232
rect 9966 359 10022 361
rect 9966 307 9968 359
rect 9968 307 10020 359
rect 10020 307 10022 359
rect 9966 305 10022 307
<< metal3 >>
rect 9945 2943 10071 2953
rect 9945 2879 9976 2943
rect 10040 2879 10071 2943
rect 9945 2870 10071 2879
rect 15754 2881 15880 2891
rect 15754 2817 15785 2881
rect 15849 2817 15880 2881
rect 15754 2807 15880 2817
rect 15759 2737 15885 2747
rect 15759 2673 15790 2737
rect 15854 2673 15885 2737
rect 15759 2663 15885 2673
rect 15760 2585 15886 2595
rect 15760 2521 15791 2585
rect 15855 2521 15886 2585
rect 15760 2511 15886 2521
rect 15760 2415 15886 2425
rect 9344 2352 9462 2353
rect 9593 2352 9737 2353
rect 9344 2338 9737 2352
rect 15760 2351 15791 2415
rect 15855 2351 15886 2415
rect 15760 2341 15886 2351
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2274 9737 2338
rect 9554 2273 9737 2274
rect 9344 2257 9737 2273
rect 15759 2258 15885 2268
rect 9449 2256 9593 2257
rect 15759 2194 15790 2258
rect 15854 2194 15885 2258
rect 15759 2184 15885 2194
rect 15677 2016 15803 2026
rect 15677 1952 15708 2016
rect 15772 1952 15803 2016
rect 15677 1942 15803 1952
rect 9484 1807 9576 1808
rect 9370 1792 9743 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9743 1792
rect 9370 1711 9743 1728
rect 15765 1755 15891 1765
rect 15765 1691 15796 1755
rect 15860 1691 15891 1755
rect 15765 1681 15891 1691
rect 15765 1552 15891 1562
rect 15765 1488 15796 1552
rect 15860 1488 15891 1552
rect 15765 1478 15891 1488
rect 15791 1477 15865 1478
rect 15675 1290 15800 1300
rect 15675 1226 15705 1290
rect 15769 1226 15800 1290
rect 15675 1216 15800 1226
rect 9932 365 10057 375
rect 9932 301 9962 365
rect 10026 301 10057 365
rect 9932 291 10057 301
<< via3 >>
rect 9976 2939 10040 2943
rect 9976 2883 9980 2939
rect 9980 2883 10036 2939
rect 10036 2883 10040 2939
rect 9976 2879 10040 2883
rect 15785 2877 15849 2881
rect 15785 2821 15789 2877
rect 15789 2821 15845 2877
rect 15845 2821 15849 2877
rect 15785 2817 15849 2821
rect 15790 2733 15854 2737
rect 15790 2677 15794 2733
rect 15794 2677 15850 2733
rect 15850 2677 15854 2733
rect 15790 2673 15854 2677
rect 15791 2581 15855 2585
rect 15791 2525 15795 2581
rect 15795 2525 15851 2581
rect 15851 2525 15855 2581
rect 15791 2521 15855 2525
rect 15791 2411 15855 2415
rect 15791 2355 15795 2411
rect 15795 2355 15851 2411
rect 15851 2355 15855 2411
rect 15791 2351 15855 2355
rect 9359 2334 9423 2338
rect 9359 2278 9363 2334
rect 9363 2278 9419 2334
rect 9419 2278 9423 2334
rect 9359 2274 9423 2278
rect 9490 2333 9554 2337
rect 9490 2277 9494 2333
rect 9494 2277 9550 2333
rect 9550 2277 9554 2333
rect 9490 2273 9554 2277
rect 9634 2334 9698 2338
rect 9634 2278 9638 2334
rect 9638 2278 9694 2334
rect 9694 2278 9698 2334
rect 9634 2274 9698 2278
rect 15790 2254 15854 2258
rect 15790 2198 15794 2254
rect 15794 2198 15850 2254
rect 15850 2198 15854 2254
rect 15790 2194 15854 2198
rect 15708 2012 15772 2016
rect 15708 1956 15712 2012
rect 15712 1956 15768 2012
rect 15768 1956 15772 2012
rect 15708 1952 15772 1956
rect 9377 1788 9441 1792
rect 9377 1732 9381 1788
rect 9381 1732 9437 1788
rect 9437 1732 9441 1788
rect 9377 1728 9441 1732
rect 9497 1788 9561 1792
rect 9497 1732 9501 1788
rect 9501 1732 9557 1788
rect 9557 1732 9561 1788
rect 9497 1728 9561 1732
rect 9640 1788 9704 1792
rect 9640 1732 9644 1788
rect 9644 1732 9700 1788
rect 9700 1732 9704 1788
rect 9640 1728 9704 1732
rect 15796 1751 15860 1755
rect 15796 1695 15800 1751
rect 15800 1695 15856 1751
rect 15856 1695 15860 1751
rect 15796 1691 15860 1695
rect 15796 1548 15860 1552
rect 15796 1492 15800 1548
rect 15800 1492 15856 1548
rect 15856 1492 15860 1548
rect 15796 1488 15860 1492
rect 15705 1286 15769 1290
rect 15705 1230 15709 1286
rect 15709 1230 15765 1286
rect 15765 1230 15769 1286
rect 15705 1226 15769 1230
rect 9962 361 10026 365
rect 9962 305 9966 361
rect 9966 305 10022 361
rect 10022 305 10026 361
rect 9962 301 10026 305
<< metal4 >>
rect 9945 2948 10071 2953
rect 9344 2943 15993 2948
rect 9344 2879 9976 2943
rect 10040 2881 15993 2943
rect 10040 2879 15785 2881
rect 9344 2870 15785 2879
rect 9344 2338 9762 2870
rect 9344 2274 9359 2338
rect 9423 2337 9634 2338
rect 9423 2274 9490 2337
rect 9344 2273 9490 2274
rect 9554 2274 9634 2337
rect 9698 2332 9762 2338
rect 15675 2817 15785 2870
rect 15849 2817 15993 2881
rect 15675 2737 15993 2817
rect 15675 2673 15790 2737
rect 15854 2673 15993 2737
rect 15675 2585 15993 2673
rect 15675 2521 15791 2585
rect 15855 2521 15993 2585
rect 15675 2415 15993 2521
rect 15675 2351 15791 2415
rect 15855 2351 15993 2415
rect 9698 2274 9761 2332
rect 9554 2273 9761 2274
rect 9344 2255 9761 2273
rect 15675 2258 15993 2351
rect 15675 2194 15790 2258
rect 15854 2194 15993 2258
rect 15675 2016 15993 2194
rect 15675 1952 15708 2016
rect 15772 1952 15993 2016
rect 15675 1940 15993 1952
rect 9370 1792 9747 1807
rect 9370 1728 9377 1792
rect 9441 1728 9497 1792
rect 9561 1728 9640 1792
rect 9704 1728 9747 1792
rect 15675 1755 15873 1765
rect 9372 369 9748 1728
rect 15675 1691 15796 1755
rect 15860 1691 15873 1755
rect 15675 1681 15873 1691
rect 15675 1300 15735 1681
rect 15933 1562 15993 1940
rect 15795 1552 15993 1562
rect 15795 1488 15796 1552
rect 15860 1488 15993 1552
rect 15795 1478 15993 1488
rect 15675 1290 15993 1300
rect 15675 1226 15705 1290
rect 15769 1226 15993 1290
rect 9932 369 10057 375
rect 15675 369 15993 1226
rect 9372 365 15993 369
rect 9372 301 9962 365
rect 10026 301 15993 365
rect 9372 291 15993 301
use hgu_nfet_hvt_stack_in_delay  hgu_nfet_hvt_stack_in_delay_0
timestamp 1699322317
transform 1 0 37644 0 1 2304
box -90 -800 5904 1051
use hgu_pfet_hvt_stack_in_delay  hgu_pfet_hvt_stack_in_delay_0
timestamp 1699322316
transform 1 0 35340 0 1 2304
box -98 -800 2214 1069
use hgu_sw_cap  hgu_sw_cap_0
timestamp 1699322316
transform 1 0 15952 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap  hgu_sw_cap_1
timestamp 1699322316
transform 1 0 32780 0 1 2352
box -53 -800 1041 1775
use hgu_sw_cap_pmos  hgu_sw_cap_pmos_0
timestamp 1699322316
transform 1 0 33874 0 1 2352
box -53 -800 1054 1856
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 32413 0 1 1600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1697965495
transform 1 0 34928 0 1 1552
box -38 -48 314 592
use hgu_sw_cap_nmos  x2
timestamp 1699184270
transform -1 0 15982 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap_nmos  x3[0]
timestamp 1699184270
transform -1 0 15248 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x3[0]
timestamp 1699322316
transform 1 0 18140 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_nmos  x3[1]
timestamp 1699184270
transform 1 0 13234 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x3[1]
timestamp 1699322316
transform 1 0 17046 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_nmos  x4[0]
timestamp 1699184270
transform -1 0 13910 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x4[0]
timestamp 1699322316
transform 1 0 22516 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_nmos  x4[1]
timestamp 1699184270
transform 1 0 11896 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x4[1]
timestamp 1699322316
transform 1 0 21422 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_nmos  x4[2]
timestamp 1699184270
transform -1 0 12698 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x4[2]
timestamp 1699322316
transform 1 0 20328 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_nmos  x4[3]
timestamp 1699184270
transform 1 0 10684 0 1 -246
box 368 546 1040 1833
use hgu_sw_cap  x4[3]
timestamp 1699322316
transform 1 0 19234 0 1 2400
box -53 -800 1041 1775
use hgu_sw_cap_pmos  x5[0]
timestamp 1699322316
transform -1 0 15984 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[0]
timestamp 1699322316
transform 1 0 31359 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[1]
timestamp 1699322316
transform 1 0 13968 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[1]
timestamp 1699322316
transform 1 0 30252 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[2]
timestamp 1699322316
transform -1 0 14772 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[2]
timestamp 1699322316
transform 1 0 29145 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[3]
timestamp 1699322316
transform 1 0 12756 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[3]
timestamp 1699322316
transform 1 0 28038 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[4]
timestamp 1699322316
transform -1 0 13560 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[4]
timestamp 1699322316
transform 1 0 26931 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[5]
timestamp 1699322316
transform 1 0 11544 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[5]
timestamp 1699322316
transform 1 0 25824 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[6]
timestamp 1699322316
transform -1 0 12348 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[6]
timestamp 1699322316
transform 1 0 24717 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[7]
timestamp 1699322316
transform 1 0 10332 0 -1 3485
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x5[7]
timestamp 1699322316
transform 1 0 23610 0 1 2400
box -53 -800 1054 1856
use hgu_sw_cap_pmos  x6
timestamp 1699322316
transform 1 0 9600 0 -1 3482
box -53 -800 1054 1856
use hgu_sw_cap_nmos  x7
timestamp 1699184270
transform 1 0 9952 0 1 -246
box 368 546 1040 1833
use hgu_pfet_hvt_stack_in_delay  x8
timestamp 1699322316
transform -1 0 10061 0 -1 2980
box -98 -800 2214 1069
use hgu_nfet_hvt_stack_in_delay  x9
timestamp 1699322317
transform -1 0 10108 0 1 536
box -90 -800 5904 1051
use sky130_fd_sc_hd__inv_1  x10
timestamp 1697965495
transform 1 0 9300 0 1 1760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x11
timestamp 1697965495
transform -1 0 9760 0 1 1760
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_MVW3GX  XM1
timestamp 1698807554
transform 1 0 15828 0 -1 1520
box -125 -130 125 68
use sky130_fd_pr__nfet_01v8_L7T3GD  XM13
timestamp 1698825334
transform 1 0 15688 0 1 1520
box -211 -252 211 252
use sky130_fd_pr__nfet_01v8_L7T3GD  XM15
timestamp 1698825334
transform 1 0 15688 0 1 1382
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM46
timestamp 1698807554
transform 1 0 15688 0 1 1723
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_hvt_M479BZ  XM47
timestamp 1698807554
transform 1 0 15688 0 1 1861
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_hvt_M433PY  XM48
timestamp 1698807554
transform 1 0 15828 0 1 1723
box -161 -139 161 90
<< labels >>
flabel metal1 9275 1596 9943 1643 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 15751 1594 15933 1640 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 9238 1979 9376 2013 0 FreeSans 320 0 0 0 code[3]
port 5 nsew
flabel metal1 14153 268 14211 1445 0 FreeSans 320 0 0 0 code[1]
port 8 nsew
flabel metal1 11727 268 11785 1445 0 FreeSans 320 0 0 0 code[2]
port 10 nsew
flabel metal4 9344 2338 9762 2948 0 FreeSans 320 0 0 0 VDD
port 17 nsew
flabel metal4 9372 291 9748 1728 0 FreeSans 320 0 0 0 VSS
port 19 nsew
flabel metal2 9702 1394 10138 1440 0 FreeSans 320 0 0 0 code_offset
port 21 nsew
flabel metal1 15009 267 15068 1448 0 FreeSans 320 0 0 0 code[0]
port 22 nsew
<< end >>
