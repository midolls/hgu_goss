magic
tech sky130A
magscale 1 2
timestamp 1698472922
<< checkpaint >>
rect -1260 -1660 1460 1460
<< pwell >>
rect 1006 1014 1032 1046
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
<< metal3 >>
rect 686 1686 1358 1688
rect 686 1622 790 1686
rect 854 1622 870 1686
rect 934 1622 950 1686
rect 1014 1622 1030 1686
rect 1094 1622 1110 1686
rect 1174 1622 1190 1686
rect 1254 1622 1358 1686
rect 686 1620 1358 1622
rect 686 1574 752 1620
rect 686 1510 687 1574
rect 751 1510 752 1574
rect 686 1494 752 1510
rect 686 1430 687 1494
rect 751 1430 752 1494
rect 686 1414 752 1430
rect 686 1350 687 1414
rect 751 1350 752 1414
rect 686 1334 752 1350
rect 686 1270 687 1334
rect 751 1270 752 1334
rect 686 1254 752 1270
rect 686 1190 687 1254
rect 751 1190 752 1254
rect 686 1174 752 1190
rect 686 1110 687 1174
rect 751 1110 752 1174
rect 686 1094 752 1110
rect 686 1030 687 1094
rect 751 1030 752 1094
rect 686 1014 752 1030
rect 686 950 687 1014
rect 751 950 752 1014
rect 686 934 752 950
rect 686 870 687 934
rect 751 870 752 934
rect 686 854 752 870
rect 686 790 687 854
rect 751 790 752 854
rect 686 726 752 790
rect 812 726 872 1620
rect 932 666 992 1560
rect 1052 726 1112 1620
rect 1292 1574 1358 1620
rect 1172 666 1232 1560
rect 1292 1510 1293 1574
rect 1357 1510 1358 1574
rect 1292 1494 1358 1510
rect 1292 1430 1293 1494
rect 1357 1430 1358 1494
rect 1292 1414 1358 1430
rect 1292 1350 1293 1414
rect 1357 1350 1358 1414
rect 1292 1334 1358 1350
rect 1292 1270 1293 1334
rect 1357 1270 1358 1334
rect 1292 1254 1358 1270
rect 1292 1190 1293 1254
rect 1357 1190 1358 1254
rect 1292 1174 1358 1190
rect 1292 1110 1293 1174
rect 1357 1110 1358 1174
rect 1292 1094 1358 1110
rect 1292 1030 1293 1094
rect 1357 1030 1358 1094
rect 1292 1014 1358 1030
rect 1292 950 1293 1014
rect 1357 950 1358 1014
rect 1292 934 1358 950
rect 1292 870 1293 934
rect 1357 870 1358 934
rect 1292 854 1358 870
rect 1292 790 1293 854
rect 1357 790 1358 854
rect 1292 726 1358 790
rect 812 664 1232 666
rect 812 600 870 664
rect 934 600 950 664
rect 1014 600 1030 664
rect 1094 600 1110 664
rect 1174 600 1232 664
rect 812 598 1232 600
<< via3 >>
rect 790 1622 854 1686
rect 870 1622 934 1686
rect 950 1622 1014 1686
rect 1030 1622 1094 1686
rect 1110 1622 1174 1686
rect 1190 1622 1254 1686
rect 687 1510 751 1574
rect 687 1430 751 1494
rect 687 1350 751 1414
rect 687 1270 751 1334
rect 687 1190 751 1254
rect 687 1110 751 1174
rect 687 1030 751 1094
rect 687 950 751 1014
rect 687 870 751 934
rect 687 790 751 854
rect 1293 1510 1357 1574
rect 1293 1430 1357 1494
rect 1293 1350 1357 1414
rect 1293 1270 1357 1334
rect 1293 1190 1357 1254
rect 1293 1110 1357 1174
rect 1293 1030 1357 1094
rect 1293 950 1357 1014
rect 1293 870 1357 934
rect 1293 790 1357 854
rect 870 600 934 664
rect 950 600 1014 664
rect 1030 600 1094 664
rect 1110 600 1174 664
<< metal4 >>
rect 686 1686 1358 1688
rect 686 1622 790 1686
rect 854 1622 870 1686
rect 934 1622 950 1686
rect 1014 1622 1030 1686
rect 1094 1622 1110 1686
rect 1174 1622 1190 1686
rect 1254 1622 1358 1686
rect 686 1620 1358 1622
rect 686 1574 752 1620
rect 686 1510 687 1574
rect 751 1510 752 1574
rect 686 1494 752 1510
rect 686 1430 687 1494
rect 751 1430 752 1494
rect 686 1414 752 1430
rect 686 1350 687 1414
rect 751 1350 752 1414
rect 686 1334 752 1350
rect 686 1270 687 1334
rect 751 1270 752 1334
rect 686 1254 752 1270
rect 686 1190 687 1254
rect 751 1190 752 1254
rect 686 1174 752 1190
rect 686 1110 687 1174
rect 751 1110 752 1174
rect 686 1094 752 1110
rect 686 1030 687 1094
rect 751 1030 752 1094
rect 686 1014 752 1030
rect 686 950 687 1014
rect 751 950 752 1014
rect 686 934 752 950
rect 686 870 687 934
rect 751 870 752 934
rect 686 854 752 870
rect 686 790 687 854
rect 751 790 752 854
rect 686 726 752 790
rect 812 666 872 1560
rect 932 726 992 1620
rect 1052 666 1112 1560
rect 1172 726 1232 1620
rect 1292 1574 1358 1620
rect 1292 1510 1293 1574
rect 1357 1510 1358 1574
rect 1292 1494 1358 1510
rect 1292 1430 1293 1494
rect 1357 1430 1358 1494
rect 1292 1414 1358 1430
rect 1292 1350 1293 1414
rect 1357 1350 1358 1414
rect 1292 1334 1358 1350
rect 1292 1270 1293 1334
rect 1357 1270 1358 1334
rect 1292 1254 1358 1270
rect 1292 1190 1293 1254
rect 1357 1190 1358 1254
rect 1292 1174 1358 1190
rect 1292 1110 1293 1174
rect 1357 1110 1358 1174
rect 1292 1094 1358 1110
rect 1292 1030 1293 1094
rect 1357 1030 1358 1094
rect 1292 1014 1358 1030
rect 1292 950 1293 1014
rect 1357 950 1358 1014
rect 1292 934 1358 950
rect 1292 870 1293 934
rect 1357 870 1358 934
rect 1292 854 1358 870
rect 1292 790 1293 854
rect 1357 790 1358 854
rect 1292 726 1358 790
rect 812 664 1232 666
rect 812 600 870 664
rect 934 600 950 664
rect 1014 600 1030 664
rect 1094 600 1110 664
rect 1174 600 1232 664
rect 812 598 1232 600
<< labels >>
flabel space 1006 1016 1032 1048 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 948 1348 974 1380 0 FreeSans 320 0 0 0 C1
port 4 nsew
flabel metal4 1066 758 1092 790 0 FreeSans 320 0 0 0 C0
port 6 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 C1
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 C0
<< end >>
