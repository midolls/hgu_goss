magic
tech sky130A
magscale 1 2
timestamp 1699450567
<< pwell >>
rect -1151 -358 1151 358
<< mvnnmos >>
rect -923 -100 -743 100
rect -685 -100 -505 100
rect -447 -100 -267 100
rect -209 -100 -29 100
rect 29 -100 209 100
rect 267 -100 447 100
rect 505 -100 685 100
rect 743 -100 923 100
<< mvndiff >>
rect -981 88 -923 100
rect -981 -88 -969 88
rect -935 -88 -923 88
rect -981 -100 -923 -88
rect -743 88 -685 100
rect -743 -88 -731 88
rect -697 -88 -685 88
rect -743 -100 -685 -88
rect -505 88 -447 100
rect -505 -88 -493 88
rect -459 -88 -447 88
rect -505 -100 -447 -88
rect -267 88 -209 100
rect -267 -88 -255 88
rect -221 -88 -209 88
rect -267 -100 -209 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 209 88 267 100
rect 209 -88 221 88
rect 255 -88 267 88
rect 209 -100 267 -88
rect 447 88 505 100
rect 447 -88 459 88
rect 493 -88 505 88
rect 447 -100 505 -88
rect 685 88 743 100
rect 685 -88 697 88
rect 731 -88 743 88
rect 685 -100 743 -88
rect 923 88 981 100
rect 923 -88 935 88
rect 969 -88 981 88
rect 923 -100 981 -88
<< mvndiffc >>
rect -969 -88 -935 88
rect -731 -88 -697 88
rect -493 -88 -459 88
rect -255 -88 -221 88
rect -17 -88 17 88
rect 221 -88 255 88
rect 459 -88 493 88
rect 697 -88 731 88
rect 935 -88 969 88
<< mvpsubdiff >>
rect -1115 310 1115 322
rect -1115 276 -1007 310
rect 1007 276 1115 310
rect -1115 264 1115 276
rect -1115 214 -1057 264
rect -1115 -214 -1103 214
rect -1069 -214 -1057 214
rect 1057 214 1115 264
rect -1115 -264 -1057 -214
rect 1057 -214 1069 214
rect 1103 -214 1115 214
rect 1057 -264 1115 -214
rect -1115 -276 1115 -264
rect -1115 -310 -1007 -276
rect 1007 -310 1115 -276
rect -1115 -322 1115 -310
<< mvpsubdiffcont >>
rect -1007 276 1007 310
rect -1103 -214 -1069 214
rect 1069 -214 1103 214
rect -1007 -310 1007 -276
<< poly >>
rect -923 172 -743 188
rect -923 138 -907 172
rect -759 138 -743 172
rect -923 100 -743 138
rect -685 172 -505 188
rect -685 138 -669 172
rect -521 138 -505 172
rect -685 100 -505 138
rect -447 172 -267 188
rect -447 138 -431 172
rect -283 138 -267 172
rect -447 100 -267 138
rect -209 172 -29 188
rect -209 138 -193 172
rect -45 138 -29 172
rect -209 100 -29 138
rect 29 172 209 188
rect 29 138 45 172
rect 193 138 209 172
rect 29 100 209 138
rect 267 172 447 188
rect 267 138 283 172
rect 431 138 447 172
rect 267 100 447 138
rect 505 172 685 188
rect 505 138 521 172
rect 669 138 685 172
rect 505 100 685 138
rect 743 172 923 188
rect 743 138 759 172
rect 907 138 923 172
rect 743 100 923 138
rect -923 -138 -743 -100
rect -923 -172 -907 -138
rect -759 -172 -743 -138
rect -923 -188 -743 -172
rect -685 -138 -505 -100
rect -685 -172 -669 -138
rect -521 -172 -505 -138
rect -685 -188 -505 -172
rect -447 -138 -267 -100
rect -447 -172 -431 -138
rect -283 -172 -267 -138
rect -447 -188 -267 -172
rect -209 -138 -29 -100
rect -209 -172 -193 -138
rect -45 -172 -29 -138
rect -209 -188 -29 -172
rect 29 -138 209 -100
rect 29 -172 45 -138
rect 193 -172 209 -138
rect 29 -188 209 -172
rect 267 -138 447 -100
rect 267 -172 283 -138
rect 431 -172 447 -138
rect 267 -188 447 -172
rect 505 -138 685 -100
rect 505 -172 521 -138
rect 669 -172 685 -138
rect 505 -188 685 -172
rect 743 -138 923 -100
rect 743 -172 759 -138
rect 907 -172 923 -138
rect 743 -188 923 -172
<< polycont >>
rect -907 138 -759 172
rect -669 138 -521 172
rect -431 138 -283 172
rect -193 138 -45 172
rect 45 138 193 172
rect 283 138 431 172
rect 521 138 669 172
rect 759 138 907 172
rect -907 -172 -759 -138
rect -669 -172 -521 -138
rect -431 -172 -283 -138
rect -193 -172 -45 -138
rect 45 -172 193 -138
rect 283 -172 431 -138
rect 521 -172 669 -138
rect 759 -172 907 -138
<< locali >>
rect -1103 276 -1007 310
rect 1007 276 1103 310
rect -1103 214 -1069 276
rect 1069 214 1103 276
rect -923 138 -907 172
rect -759 138 -743 172
rect -685 138 -669 172
rect -521 138 -505 172
rect -447 138 -431 172
rect -283 138 -267 172
rect -209 138 -193 172
rect -45 138 -29 172
rect 29 138 45 172
rect 193 138 209 172
rect 267 138 283 172
rect 431 138 447 172
rect 505 138 521 172
rect 669 138 685 172
rect 743 138 759 172
rect 907 138 923 172
rect -969 88 -935 104
rect -969 -104 -935 -88
rect -731 88 -697 104
rect -731 -104 -697 -88
rect -493 88 -459 104
rect -493 -104 -459 -88
rect -255 88 -221 104
rect -255 -104 -221 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 221 88 255 104
rect 221 -104 255 -88
rect 459 88 493 104
rect 459 -104 493 -88
rect 697 88 731 104
rect 697 -104 731 -88
rect 935 88 969 104
rect 935 -104 969 -88
rect -923 -172 -907 -138
rect -759 -172 -743 -138
rect -685 -172 -669 -138
rect -521 -172 -505 -138
rect -447 -172 -431 -138
rect -283 -172 -267 -138
rect -209 -172 -193 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 193 -172 209 -138
rect 267 -172 283 -138
rect 431 -172 447 -138
rect 505 -172 521 -138
rect 669 -172 685 -138
rect 743 -172 759 -138
rect 907 -172 923 -138
rect -1103 -276 -1069 -214
rect 1069 -276 1103 -214
rect -1103 -310 -1007 -276
rect 1007 -310 1103 -276
<< viali >>
rect -907 138 -759 172
rect -669 138 -521 172
rect -431 138 -283 172
rect -193 138 -45 172
rect 45 138 193 172
rect 283 138 431 172
rect 521 138 669 172
rect 759 138 907 172
rect -969 -88 -935 88
rect -731 -88 -697 88
rect -493 -88 -459 88
rect -255 -88 -221 88
rect -17 -88 17 88
rect 221 -88 255 88
rect 459 -88 493 88
rect 697 -88 731 88
rect 935 -88 969 88
rect -907 -172 -759 -138
rect -669 -172 -521 -138
rect -431 -172 -283 -138
rect -193 -172 -45 -138
rect 45 -172 193 -138
rect 283 -172 431 -138
rect 521 -172 669 -138
rect 759 -172 907 -138
<< metal1 >>
rect -919 172 -747 178
rect -919 138 -907 172
rect -759 138 -747 172
rect -919 132 -747 138
rect -681 172 -509 178
rect -681 138 -669 172
rect -521 138 -509 172
rect -681 132 -509 138
rect -443 172 -271 178
rect -443 138 -431 172
rect -283 138 -271 172
rect -443 132 -271 138
rect -205 172 -33 178
rect -205 138 -193 172
rect -45 138 -33 172
rect -205 132 -33 138
rect 33 172 205 178
rect 33 138 45 172
rect 193 138 205 172
rect 33 132 205 138
rect 271 172 443 178
rect 271 138 283 172
rect 431 138 443 172
rect 271 132 443 138
rect 509 172 681 178
rect 509 138 521 172
rect 669 138 681 172
rect 509 132 681 138
rect 747 172 919 178
rect 747 138 759 172
rect 907 138 919 172
rect 747 132 919 138
rect -975 88 -929 100
rect -975 -88 -969 88
rect -935 -88 -929 88
rect -975 -100 -929 -88
rect -737 88 -691 100
rect -737 -88 -731 88
rect -697 -88 -691 88
rect -737 -100 -691 -88
rect -499 88 -453 100
rect -499 -88 -493 88
rect -459 -88 -453 88
rect -499 -100 -453 -88
rect -261 88 -215 100
rect -261 -88 -255 88
rect -221 -88 -215 88
rect -261 -100 -215 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 215 88 261 100
rect 215 -88 221 88
rect 255 -88 261 88
rect 215 -100 261 -88
rect 453 88 499 100
rect 453 -88 459 88
rect 493 -88 499 88
rect 453 -100 499 -88
rect 691 88 737 100
rect 691 -88 697 88
rect 731 -88 737 88
rect 691 -100 737 -88
rect 929 88 975 100
rect 929 -88 935 88
rect 969 -88 975 88
rect 929 -100 975 -88
rect -919 -138 -747 -132
rect -919 -172 -907 -138
rect -759 -172 -747 -138
rect -919 -178 -747 -172
rect -681 -138 -509 -132
rect -681 -172 -669 -138
rect -521 -172 -509 -138
rect -681 -178 -509 -172
rect -443 -138 -271 -132
rect -443 -172 -431 -138
rect -283 -172 -271 -138
rect -443 -178 -271 -172
rect -205 -138 -33 -132
rect -205 -172 -193 -138
rect -45 -172 -33 -138
rect -205 -178 -33 -172
rect 33 -138 205 -132
rect 33 -172 45 -138
rect 193 -172 205 -138
rect 33 -178 205 -172
rect 271 -138 443 -132
rect 271 -172 283 -138
rect 431 -172 443 -138
rect 271 -178 443 -172
rect 509 -138 681 -132
rect 509 -172 521 -138
rect 669 -172 681 -138
rect 509 -178 681 -172
rect 747 -138 919 -132
rect 747 -172 759 -138
rect 907 -172 919 -138
rect 747 -178 919 -172
<< properties >>
string FIXED_BBOX -1086 -293 1086 293
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 1.0 l 0.9 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
