magic
tech sky130A
timestamp 1698913202
<< nwell >>
rect -19 618 295 625
rect -19 536 296 618
rect 295 529 296 536
<< psubdiff >>
rect 1 293 277 295
rect 1 276 78 293
rect 95 276 277 293
<< nsubdiff >>
rect 0 594 276 595
rect 0 577 61 594
rect 78 577 276 594
rect 0 576 276 577
<< psubdiffcont >>
rect 78 276 95 293
<< nsubdiffcont >>
rect 61 577 78 594
<< locali >>
rect 53 594 86 595
rect 53 578 61 594
rect 78 578 86 594
rect 85 410 193 427
rect 69 293 103 294
rect 69 276 78 293
rect 95 276 103 293
<< viali >>
rect 37 409 54 426
rect 225 412 242 429
<< metal1 >>
rect 0 554 275 603
rect 219 429 304 433
rect -27 426 62 429
rect -27 409 37 426
rect 54 409 62 426
rect -27 405 62 409
rect 219 412 225 429
rect 242 412 304 429
rect 219 408 304 412
rect -27 404 53 405
rect 0 265 275 314
use sky130_fd_sc_hd__inv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697965495
transform 1 0 0 0 1 300
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x2
timestamp 1697965495
transform 1 0 138 0 1 300
box -19 -24 157 296
<< labels >>
flabel metal1 0 554 275 603 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 0 265 275 314 0 FreeSans 160 0 0 0 VSS
port 1 nsew
flabel metal1 -27 404 53 429 0 FreeSans 160 0 0 0 in
port 2 nsew
flabel metal1 224 408 304 433 0 FreeSans 160 0 0 0 out
port 4 nsew
<< end >>
