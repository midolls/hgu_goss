magic
tech sky130A
timestamp 1699890160
<< psubdiff >>
rect 1046 2019 1068 2069
<< metal4 >>
rect 772 2096 795 2142
rect 1136 2107 1159 2153
rect 836 1681 856 1723
use hgu_cdac_unit  x1[0]
timestamp 1699890160
transform 1 0 0 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[1]
timestamp 1699890160
transform -1 0 1022 0 -1 2892
box 343 299 679 913
use hgu_cdac_unit  x1[2]
timestamp 1699890160
transform 1 0 303 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[3]
timestamp 1699890160
transform -1 0 1325 0 -1 2892
box 343 299 679 913
use hgu_cdac_unit  x1[4]
timestamp 1699890160
transform 1 0 606 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[5]
timestamp 1699890160
transform -1 0 1628 0 -1 2892
box 343 299 679 913
use hgu_cdac_unit  x1[6]
timestamp 1699890160
transform 1 0 909 0 1 1100
box 343 299 679 913
use hgu_cdac_unit  x1[7]
timestamp 1699890160
transform -1 0 1931 0 -1 2892
box 343 299 679 913
<< labels >>
flabel psubdiff 1046 2019 1068 2069 0 FreeSans 160 0 0 0 SUB
port 1 nsew
flabel metal4 1136 2107 1159 2153 0 FreeSans 160 0 0 0 CBOT
port 3 nsew
flabel metal4 772 2096 795 2142 0 FreeSans 160 0 0 0 CTOP
port 5 nsew
flabel metal4 836 1681 856 1723 0 FreeSans 160 0 0 0 CTOP
port 8 nsew
<< end >>
