* NGSPICE file created from edit_distance_state.ext - technology: sky130A

.subckt edit_distance_state in out VSS VDD
X0 x2.A in.t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1 out.t0 x2.A VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2 x2.A in.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3 out.t1 x2.A VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 in.n0 in.t0 230.502
R1 in.n0 in.t1 157.821
R2 in.n1 in.n0 8.66327
R3 in in.n1 3.61504
R4 in.n1 in 2.02684
R5 VDD.n7 VDD 551.928
R6 VDD VDD.t2 258.87
R7 VDD.t0 VDD 258.87
R8 VDD.n0 VDD.t3 164.91
R9 VDD.n15 VDD.t1 152.88
R10 VDD.n6 VDD.n5 50.5268
R11 VDD.n8 VDD.n7 39.0751
R12 VDD.n16 VDD.n15 20.8387
R13 VDD.n14 VDD.n13 9.3005
R14 VDD.n11 VDD.n10 9.3005
R15 VDD.n10 VDD.n9 9.3005
R16 VDD.n9 VDD.t0 7.32698
R17 VDD.n4 VDD.n3 6.02403
R18 VDD.n10 VDD.n6 3.15839
R19 VDD.n12 VDD.n11 3.1005
R20 VDD.n9 VDD.n8 2.44266
R21 VDD.n0 VDD 0.563874
R22 VDD.n11 VDD.n4 0.376971
R23 VDD.n1 VDD 0.352541
R24 VDD.n12 VDD.n2 0.105045
R25 VDD.n1 VDD 0.0974388
R26 VDD.n16 VDD.n14 0.0857273
R27 VDD VDD.n0 0.0745681
R28 VDD.n2 VDD.n1 0.0527727
R29 VDD.n14 VDD.n12 0.0198182
R30 VDD VDD.n16 0.0198182
R31 out.n0 out.t0 137.917
R32 out out.t1 106.635
R33 out.n1 out 13.357
R34 out out.n1 5.56572
R35 out.n1 out 4.66888
R36 out out.n0 2.22659
R37 out.n0 out 1.55202
R38 VSS.n3 VSS 2764.95
R39 VSS VSS.t2 1409.06
R40 VSS.t0 VSS 1409.06
R41 VSS.n4 VSS.n3 585
R42 VSS.n3 VSS.t0 505.137
R43 VSS.n0 VSS.t3 118.326
R44 VSS.n7 VSS.t1 111.924
R45 VSS.n8 VSS.n7 11.427
R46 VSS.n5 VSS.n4 6.89281
R47 VSS.n6 VSS.n5 4.6505
R48 VSS.n0 VSS 0.553346
R49 VSS.n1 VSS 0.352541
R50 VSS.n6 VSS.n2 0.0979576
R51 VSS.n8 VSS.n6 0.0979576
R52 VSS.n1 VSS 0.0974388
R53 VSS VSS.n0 0.0662933
R54 VSS.n2 VSS.n1 0.0492288
R55 VSS VSS.n8 0.0185085
C0 VDD VSS 1.19f
.ends

