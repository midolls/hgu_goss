** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_clk_async.sch
**.subckt hgu_clk_async VDD ASYNC_CLK_SAR VSS sample_clk EOC READY
*.ipin VDD
*.opin ASYNC_CLK_SAR
*.ipin VSS
*.ipin sample_clk
*.ipin EOC
*.ipin READY
x3 net2 VSS sample_clk VGND VNB VPB VPWR net4 sky130_fd_sc_hd__mux2_1
x8 net4 VSS EOC VGND VNB VPB VPWR ASYNC_CLK_SAR sky130_fd_sc_hd__mux2_1
x27 sample_clk VDD net5 net6 VGND VNB VPB VPWR net2 net7 sky130_fd_sc_hd__dfbbp_1
x9 net1 VGND VNB VPB VPWR net6 sky130_fd_sc_hd__inv_1
x10 net3 VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
C1 net1 VSS 5f m=1
C2 net3 VSS 5f m=1
C3 net2 VSS 5f m=1
C4 net4 VSS 5f m=1
x2 VDD READY net1 VSS hgu_delay_no_code
x4 VDD ASYNC_CLK_SAR net3 VSS hgu_delay_no_code
**.ends

* expanding   symbol:  hgu_delay_no_code.sym # of pins=4
** sym_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sym
** sch_path: /foss/designs/hgu_goss/hgu/xschem/hgu_delay_no_code.sch
.subckt hgu_delay_no_code VDD IN OUT VSS
*.ipin IN
*.ipin VDD
*.ipin VSS
*.opin OUT
XM1 net1 IN VSS VSS sky130_fd_pr__nfet_01v8 L=3.69 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 IN VDD VDD sky130_fd_pr__pfet_01v8 L=1.5 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 VSS net1 VSS VSS sky130_fd_pr__nfet_01v8 L=2.045 W=1.375 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 OUT net1 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 OUT net1 net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 VDD OUT net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS OUT net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
