magic
tech sky130A
magscale 1 2
timestamp 1699484509
<< error_s >>
rect 1098 5136 1148 5141
rect 1178 5136 1244 5141
rect 1274 5136 1340 5141
rect 1370 5136 1436 5141
rect 1562 5136 1628 5143
rect 1692 5139 1708 5140
rect 1146 5091 1148 5122
rect 1178 5091 1244 5122
rect 1274 5091 1340 5122
rect 1370 5091 1436 5122
rect 1562 5093 1628 5124
rect 1708 5108 1724 5124
rect 1518 3988 1576 3994
rect 1518 3954 1530 3988
rect 1518 3948 1576 3954
rect 1579 2627 1595 2643
rect 1597 2627 1613 2643
rect 1675 2627 1691 2643
rect 1693 2627 1709 2643
rect 1563 2611 1579 2627
rect 1613 2611 1629 2627
rect 1659 2611 1675 2627
rect 1709 2611 1725 2627
rect 985 1384 1820 1409
rect 959 1373 1849 1381
rect 949 1348 1856 1373
<< nwell >>
rect 1482 5138 1509 5140
rect 1589 5138 1708 5139
rect 1098 5082 1132 5131
rect 1290 5124 1324 5137
rect 1148 5093 1466 5124
rect 1481 5105 1708 5138
rect 1481 5104 1666 5105
rect 1482 5103 1509 5104
rect 1290 5088 1324 5093
rect 1578 5089 1612 5104
rect 1487 4022 1601 4036
rect 1487 4018 1507 4022
rect 1593 4018 1601 4022
rect 1487 4015 1601 4018
rect 1487 4011 1593 4015
rect 1487 3933 1502 4011
rect 1507 3940 1593 4011
rect 1594 3933 1601 4015
rect 1487 3916 1601 3933
rect 1487 3883 1614 3916
rect 949 3845 1858 3883
<< nsubdiff >>
rect 1498 3881 1614 3916
<< poly >>
rect 1146 5091 1465 5122
rect 1532 5093 1658 5124
rect 1532 4004 1562 4010
rect 1514 3988 1580 4004
rect 1514 3954 1530 3988
rect 1564 3954 1580 3988
rect 1514 3940 1580 3954
rect 1147 3635 1466 3666
rect 1532 3635 1658 3666
<< polycont >>
rect 1530 3954 1564 3988
<< locali >>
rect 1098 5105 1708 5139
rect 1098 5055 1132 5105
rect 1290 5055 1324 5105
rect 1482 5075 1483 5104
rect 1482 5055 1516 5075
rect 1578 5055 1612 5105
rect 1674 5055 1708 5105
rect 1514 3954 1530 3988
rect 1564 3954 1580 3988
rect 1498 3881 1614 3916
<< viali >>
rect 1530 3954 1564 3988
<< metal1 >>
rect 1518 3988 1576 3994
rect 1290 3671 1324 3979
rect 1518 3954 1530 3988
rect 1564 3954 1576 3988
rect 1518 3948 1576 3954
rect 1674 3759 1708 4036
rect 1292 1239 1326 1492
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_0
timestamp 1699479866
transform 1 0 1595 0 1 3334
box -204 -473 227 1797
use sky130_fd_pr__nfet_01v8_5AY3TR  sky130_fd_pr__nfet_01v8_5AY3TR_3
timestamp 1699479866
transform 1 0 1596 0 1 906
box -204 -473 227 1797
use sky130_fd_pr__nfet_01v8_YCY3T5  sky130_fd_pr__nfet_01v8_YCY3T5_2
timestamp 1699479866
transform 1 0 1308 0 1 906
box -323 -449 289 449
use sky130_fd_pr__pfet_01v8_UJB66J  sky130_fd_pr__pfet_01v8_UJB66J_2
timestamp 1699484509
transform 1 0 1596 0 1 2089
box -399 -741 263 769
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_0
timestamp 1699484509
transform 1 0 1307 0 1 4586
box -359 -741 551 905
use sky130_fd_pr__pfet_01v8_UJKTUG  sky130_fd_pr__pfet_01v8_UJKTUG_3
timestamp 1699484509
transform 1 0 1308 0 1 2089
box -359 -741 551 905
use sky130_fd_pr__pfet_01v8_UJB66J  XM1
timestamp 1699484509
transform 1 0 1595 0 1 4586
box -399 -741 263 769
use sky130_fd_pr__nfet_01v8_YCY3T5  XM4
timestamp 1699479866
transform 1 0 1307 0 1 3334
box -323 -449 289 449
<< labels >>
flabel space 1675 1169 1709 1551 0 FreeSans 320 0 0 0 tah_vn
port 5 nsew
flabel metal1 1300 1355 1320 1384 0 FreeSans 320 0 0 0 vin
port 8 nsew
flabel metal1 1294 3797 1317 3826 0 FreeSans 320 0 0 0 vip
port 3 nsew
<< end >>
