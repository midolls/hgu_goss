* NGSPICE file created from hgu_delay_no_code_flat.ext - technology: sky130A

.subckt hgu_delay_no_code_flat IN OUT code[3] code[1] code[2] code[0] code_offset
+ VSS VDD
X0 x9.output_stack x10.Y.t2 x5[7].floating.t7 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X1 x9.output_stack code[2].t0 x4[3].floating VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X2 x5[7].floating.t6 x10.Y.t3 x9.output_stack VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X3 x9.output_stack code_offset.t0 x7.floating VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X4 a_15703_1340# OUT.t2 VDD.t15 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 x3[1].floating code[1].t0 x9.output_stack VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X6 a_9893_879# IN.t0 a_9805_879# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X7 a_9965_465# IN.t1 a_9893_465# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_9918_2268# IN.t2 a_9830_2130# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X9 a_9965_1017# IN.t3 a_9893_1017# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_9918_2544# IN.t4 a_9830_2682# VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_15703_1340# x9.output_stack VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X12 a_15703_1681# x9.output_stack OUT.t1 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X13 x4[3].floating code[2].t1 x9.output_stack VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X14 VDD.t3 OUT.t3 a_15703_1340# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_9893_465# IN.t5 a_9805_327# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X16 VDD.t10 code_offset.t1 x6.SW VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X17 VSS.t10 IN.t6 a_9893_327# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 x9.output_stack x10.Y.t4 x5[7].floating.t5 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X19 x5[7].floating.t4 x10.Y.t5 x9.output_stack VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X20 a_9918_2544# IN.t7 a_9830_2406# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X21 x9.output_stack code[1].t1 x3[1].floating VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X22 a_9965_741# IN.t8 a_9893_741# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 a_9893_327# IN.t9 a_9805_327# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X24 x10.Y.t1 code[3].t0 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X25 a_15703_1681# x9.output_stack VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X26 x9.output_stack x6.SW x6.floating VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X27 VSS.t12 code_offset.t2 x6.SW VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X28 a_9893_1293# IN.t10 a_9805_1155# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X29 x5[7].floating.t3 x10.Y.t6 x9.output_stack VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X30 a_15703_1681# OUT.t4 VSS.t6 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X31 a_9893_741# IN.t11 a_9805_603# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X32 x9.output_stack IN.t12 a_9830_2130# VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X33 x5[7].floating.t2 x10.Y.t7 x9.output_stack VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.101 ps=0.9 w=0.42 l=0.15
X34 x9.output_stack x10.Y.t8 x5[7].floating.t1 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X35 x9.output_stack code[2].t2 x4[3].floating VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.122 ps=1.42 w=0.42 l=0.15
X36 a_9965_465# IN.t13 a_9893_603# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X37 a_9918_2268# IN.t14 a_9830_2406# VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X38 x4[3].floating code[2].t3 x9.output_stack VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0966 ps=0.88 w=0.42 l=0.15
X39 a_15703_1340# x9.output_stack OUT.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0651 pd=0.73 as=0.122 ps=1.42 w=0.42 l=0.15
X40 x9.output_stack IN.t15 a_9893_1293# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X41 x10.Y.t0 code[3].t1 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X42 a_9893_1155# IN.t16 a_9805_1155# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X43 VDD.t6 IN.t17 a_9830_2682# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X44 x9.output_stack x10.Y.t9 x5[7].floating.t0 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.101 pd=0.9 as=0.122 ps=1.42 w=0.42 l=0.15
X45 VSS.t5 OUT.t5 a_15703_1681# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0651 ps=0.73 w=0.42 l=0.15
X46 x2.floating code[0].t0 x9.output_stack VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.124 ps=1.43 w=0.42 l=0.15
X47 a_9893_603# IN.t18 a_9805_603# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
X48 a_9965_1017# IN.t19 a_9893_1155# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X49 a_9965_741# IN.t20 a_9893_879# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0441 ps=0.63 w=0.42 l=0.15
X50 a_9893_1017# IN.t21 a_9805_879# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.122 ps=1.42 w=0.42 l=0.15
R0 x10.Y x10.Y.t6 154.847
R1 x10.Y x10.Y.t8 154.8
R2 x10.Y x10.Y.t7 154.8
R3 x10.Y x10.Y.t2 154.8
R4 x10.Y x10.Y.t3 154.8
R5 x10.Y x10.Y.t4 154.8
R6 x10.Y x10.Y.t5 154.8
R7 x10.Y x10.Y.t9 154.8
R8 x10.Y.n0 x10.Y 134.239
R9 x10.Y x10.Y.t0 106.635
R10 x10.Y.n2 x10.Y.t1 24.6567
R11 x10.Y.n5 x10.Y.n4 12.4089
R12 x10.Y.n3 x10.Y.n2 9.12522
R13 x10.Y.n4 x10.Y.n3 7.34048
R14 x10.Y.n5 x10.Y 2.22659
R15 x10.Y.n2 x10.Y.n1 1.93377
R16 x10.Y x10.Y.n5 1.55202
R17 x10.Y.n3 x10.Y.n0 0.69928
R18 x5[7].floating.n95 x5[7].floating.t7 68.0345
R19 x5[7].floating.n24 x5[7].floating.t2 68.0345
R20 x5[7].floating.n42 x5[7].floating.t1 68.0345
R21 x5[7].floating.n54 x5[7].floating.t3 68.0345
R22 x5[7].floating.n154 x5[7].floating.t0 68.0345
R23 x5[7].floating.n142 x5[7].floating.t4 68.0345
R24 x5[7].floating.n12 x5[7].floating.t5 68.0345
R25 x5[7].floating.n109 x5[7].floating.t6 68.0345
R26 x5[7].floating.n73 x5[7].floating.n35 0.660401
R27 x5[7].floating.n91 x5[7].floating.n90 0.660401
R28 x5[7].floating.n130 x5[7].floating.n20 0.660401
R29 x5[7].floating.n139 x5[7].floating.n5 0.660401
R30 x5[7].floating.n121 x5[7].floating.n120 0.660401
R31 x5[7].floating.n60 x5[7].floating.n59 0.320345
R32 x5[7].floating.n160 x5[7].floating.n159 0.308269
R33 x5[7].floating.n161 x5[7].floating.n160 0.173084
R34 x5[7].floating.n61 x5[7].floating.n60 0.162103
R35 x5[7].floating.n160 x5[7].floating 0.100688
R36 x5[7].floating.n60 x5[7].floating 0.0755007
R37 x5[7].floating.n36 x5[7].floating.n35 0.0716912
R38 x5[7].floating.n35 x5[7].floating.n34 0.0716912
R39 x5[7].floating.n6 x5[7].floating.n5 0.0716912
R40 x5[7].floating.n5 x5[7].floating.n4 0.0716912
R41 x5[7].floating.n74 x5[7].floating.n73 0.0716912
R42 x5[7].floating.n122 x5[7].floating.n121 0.0716912
R43 x5[7].floating.n140 x5[7].floating.n139 0.0716912
R44 x5[7].floating.n120 x5[7].floating.n105 0.0716912
R45 x5[7].floating.n120 x5[7].floating.n119 0.0716912
R46 x5[7].floating.n40 x5[7].floating.n39 0.0557941
R47 x5[7].floating.n39 x5[7].floating.n38 0.0557941
R48 x5[7].floating.n38 x5[7].floating.n37 0.0557941
R49 x5[7].floating.n37 x5[7].floating.n36 0.0557941
R50 x5[7].floating.n34 x5[7].floating.n33 0.0557941
R51 x5[7].floating.n33 x5[7].floating.n32 0.0557941
R52 x5[7].floating.n32 x5[7].floating.n31 0.0557941
R53 x5[7].floating.n31 x5[7].floating.n30 0.0557941
R54 x5[7].floating.n10 x5[7].floating.n9 0.0557941
R55 x5[7].floating.n9 x5[7].floating.n8 0.0557941
R56 x5[7].floating.n8 x5[7].floating.n7 0.0557941
R57 x5[7].floating.n7 x5[7].floating.n6 0.0557941
R58 x5[7].floating.n4 x5[7].floating.n3 0.0557941
R59 x5[7].floating.n3 x5[7].floating.n2 0.0557941
R60 x5[7].floating.n2 x5[7].floating.n1 0.0557941
R61 x5[7].floating.n1 x5[7].floating.n0 0.0557941
R62 x5[7].floating.n69 x5[7].floating.n68 0.0557941
R63 x5[7].floating.n70 x5[7].floating.n69 0.0557941
R64 x5[7].floating.n71 x5[7].floating.n70 0.0557941
R65 x5[7].floating.n72 x5[7].floating.n71 0.0557941
R66 x5[7].floating.n76 x5[7].floating.n75 0.0557941
R67 x5[7].floating.n77 x5[7].floating.n76 0.0557941
R68 x5[7].floating.n78 x5[7].floating.n77 0.0557941
R69 x5[7].floating.n86 x5[7].floating.n85 0.0557941
R70 x5[7].floating.n85 x5[7].floating.n84 0.0557941
R71 x5[7].floating.n84 x5[7].floating.n83 0.0557941
R72 x5[7].floating.n83 x5[7].floating.n82 0.0557941
R73 x5[7].floating.n124 x5[7].floating.n123 0.0557941
R74 x5[7].floating.n125 x5[7].floating.n124 0.0557941
R75 x5[7].floating.n126 x5[7].floating.n125 0.0557941
R76 x5[7].floating.n135 x5[7].floating.n134 0.0557941
R77 x5[7].floating.n136 x5[7].floating.n135 0.0557941
R78 x5[7].floating.n137 x5[7].floating.n136 0.0557941
R79 x5[7].floating.n138 x5[7].floating.n137 0.0557941
R80 x5[7].floating.n171 x5[7].floating.n170 0.0557941
R81 x5[7].floating.n170 x5[7].floating.n169 0.0557941
R82 x5[7].floating.n169 x5[7].floating.n168 0.0557941
R83 x5[7].floating.n102 x5[7].floating.n101 0.0557941
R84 x5[7].floating.n103 x5[7].floating.n102 0.0557941
R85 x5[7].floating.n104 x5[7].floating.n103 0.0557941
R86 x5[7].floating.n105 x5[7].floating.n104 0.0557941
R87 x5[7].floating.n119 x5[7].floating.n118 0.0557941
R88 x5[7].floating.n118 x5[7].floating.n117 0.0557941
R89 x5[7].floating.n117 x5[7].floating.n116 0.0557941
R90 x5[7].floating.n116 x5[7].floating.n115 0.0557941
R91 x5[7].floating.n65 x5[7].floating.n64 0.0537206
R92 x5[7].floating.n90 x5[7].floating.n89 0.0537206
R93 x5[7].floating.n131 x5[7].floating.n130 0.0537206
R94 x5[7].floating.n164 x5[7].floating.n163 0.0537206
R95 x5[7].floating.n64 x5[7].floating.n63 0.0530294
R96 x5[7].floating.n90 x5[7].floating.n81 0.0530294
R97 x5[7].floating.n130 x5[7].floating.n129 0.0530294
R98 x5[7].floating.n165 x5[7].floating.n164 0.0530294
R99 x5[7].floating.n92 x5[7].floating.n91 0.0529559
R100 x5[7].floating.n50 x5[7].floating.n49 0.0529559
R101 x5[7].floating.n20 x5[7].floating.n19 0.0529559
R102 x5[7].floating.n151 x5[7].floating.n150 0.0529559
R103 x5[7].floating.n51 x5[7].floating.n50 0.0524559
R104 x5[7].floating.n91 x5[7].floating.n21 0.0524559
R105 x5[7].floating.n106 x5[7].floating.n20 0.0524559
R106 x5[7].floating.n150 x5[7].floating.n149 0.0524559
R107 x5[7].floating.n79 x5[7].floating.n78 0.0523382
R108 x5[7].floating.n127 x5[7].floating.n126 0.0523382
R109 x5[7].floating.n168 x5[7].floating.n167 0.0523382
R110 x5[7].floating.n68 x5[7].floating.n67 0.0516471
R111 x5[7].floating.n87 x5[7].floating.n86 0.0516471
R112 x5[7].floating.n134 x5[7].floating.n133 0.0516471
R113 x5[7].floating.n73 x5[7].floating 0.0495735
R114 x5[7].floating.n121 x5[7].floating 0.0495735
R115 x5[7].floating.n139 x5[7].floating 0.0495735
R116 x5[7].floating.n98 x5[7].floating.n97 0.0408846
R117 x5[7].floating.n45 x5[7].floating.n44 0.0408846
R118 x5[7].floating.n157 x5[7].floating.n156 0.0408846
R119 x5[7].floating.n15 x5[7].floating.n14 0.0408846
R120 x5[7].floating.n75 x5[7].floating 0.0336765
R121 x5[7].floating.n123 x5[7].floating 0.0336765
R122 x5[7].floating x5[7].floating.n171 0.0336765
R123 x5[7].floating.n30 x5[7].floating.n29 0.0271618
R124 x5[7].floating.n115 x5[7].floating.n114 0.0271618
R125 x5[7].floating.n101 x5[7].floating.n100 0.0266618
R126 x5[7].floating.n41 x5[7].floating.n40 0.0266618
R127 x5[7].floating.n11 x5[7].floating.n10 0.0266618
R128 x5[7].floating x5[7].floating.n72 0.0226176
R129 x5[7].floating x5[7].floating.n74 0.0226176
R130 x5[7].floating.n82 x5[7].floating 0.0226176
R131 x5[7].floating x5[7].floating.n122 0.0226176
R132 x5[7].floating x5[7].floating.n138 0.0226176
R133 x5[7].floating x5[7].floating.n140 0.0226176
R134 x5[7].floating.n63 x5[7].floating.n62 0.0191618
R135 x5[7].floating.n81 x5[7].floating.n80 0.0191618
R136 x5[7].floating.n129 x5[7].floating.n128 0.0191618
R137 x5[7].floating.n166 x5[7].floating.n165 0.0191618
R138 x5[7].floating.n66 x5[7].floating.n65 0.0184706
R139 x5[7].floating.n89 x5[7].floating.n88 0.0184706
R140 x5[7].floating.n132 x5[7].floating.n131 0.0184706
R141 x5[7].floating.n163 x5[7].floating.n162 0.0184706
R142 x5[7].floating.n100 x5[7].floating.n99 0.014
R143 x5[7].floating.n52 x5[7].floating.n51 0.014
R144 x5[7].floating.n46 x5[7].floating.n41 0.014
R145 x5[7].floating.n22 x5[7].floating.n21 0.014
R146 x5[7].floating.n16 x5[7].floating.n11 0.014
R147 x5[7].floating.n149 x5[7].floating.n148 0.014
R148 x5[7].floating.n159 x5[7].floating.n158 0.014
R149 x5[7].floating.n107 x5[7].floating.n106 0.014
R150 x5[7].floating.n93 x5[7].floating.n92 0.0135
R151 x5[7].floating.n59 x5[7].floating.n58 0.0135
R152 x5[7].floating.n49 x5[7].floating.n48 0.0135
R153 x5[7].floating.n29 x5[7].floating.n28 0.0135
R154 x5[7].floating.n19 x5[7].floating.n18 0.0135
R155 x5[7].floating.n146 x5[7].floating.n141 0.0135
R156 x5[7].floating.n152 x5[7].floating.n151 0.0135
R157 x5[7].floating.n114 x5[7].floating.n113 0.0135
R158 x5[7].floating.n27 x5[7].floating.n26 0.0120385
R159 x5[7].floating.n57 x5[7].floating.n56 0.0120385
R160 x5[7].floating.n145 x5[7].floating.n144 0.0120385
R161 x5[7].floating.n112 x5[7].floating.n111 0.0120385
R162 x5[7].floating.n67 x5[7].floating.n66 0.00464706
R163 x5[7].floating.n88 x5[7].floating.n87 0.00464706
R164 x5[7].floating.n133 x5[7].floating.n132 0.00464706
R165 x5[7].floating.n162 x5[7].floating.n161 0.00464706
R166 x5[7].floating.n62 x5[7].floating.n61 0.00395588
R167 x5[7].floating.n80 x5[7].floating.n79 0.00395588
R168 x5[7].floating.n128 x5[7].floating.n127 0.00395588
R169 x5[7].floating.n167 x5[7].floating.n166 0.00395588
R170 x5[7].floating.n110 x5[7].floating.n109 0.00359614
R171 x5[7].floating.n25 x5[7].floating.n24 0.00359614
R172 x5[7].floating.n55 x5[7].floating.n54 0.00359614
R173 x5[7].floating.n143 x5[7].floating.n142 0.00359614
R174 x5[7].floating.n94 x5[7].floating.n93 0.0035
R175 x5[7].floating.n58 x5[7].floating.n53 0.0035
R176 x5[7].floating.n48 x5[7].floating.n47 0.0035
R177 x5[7].floating.n28 x5[7].floating.n23 0.0035
R178 x5[7].floating.n18 x5[7].floating.n17 0.0035
R179 x5[7].floating.n147 x5[7].floating.n146 0.0035
R180 x5[7].floating.n153 x5[7].floating.n152 0.0035
R181 x5[7].floating.n113 x5[7].floating.n108 0.0035
R182 x5[7].floating.n99 x5[7].floating.n94 0.003
R183 x5[7].floating.n53 x5[7].floating.n52 0.003
R184 x5[7].floating.n47 x5[7].floating.n46 0.003
R185 x5[7].floating.n23 x5[7].floating.n22 0.003
R186 x5[7].floating.n17 x5[7].floating.n16 0.003
R187 x5[7].floating.n148 x5[7].floating.n147 0.003
R188 x5[7].floating.n158 x5[7].floating.n153 0.003
R189 x5[7].floating.n108 x5[7].floating.n107 0.003
R190 x5[7].floating.n155 x5[7].floating.n154 0.00277942
R191 x5[7].floating.n96 x5[7].floating.n95 0.0023396
R192 x5[7].floating.n43 x5[7].floating.n42 0.0023396
R193 x5[7].floating.n13 x5[7].floating.n12 0.0023396
R194 x5[7].floating.n157 x5[7].floating.n155 0.00233747
R195 x5[7].floating.n98 x5[7].floating.n96 0.00200689
R196 x5[7].floating.n45 x5[7].floating.n43 0.00200689
R197 x5[7].floating.n15 x5[7].floating.n13 0.00200689
R198 x5[7].floating.n27 x5[7].floating.n25 0.0010233
R199 x5[7].floating.n57 x5[7].floating.n55 0.0010233
R200 x5[7].floating.n145 x5[7].floating.n143 0.0010233
R201 x5[7].floating.n112 x5[7].floating.n110 0.0010233
R202 x5[7].floating.n99 x5[7].floating.n98 0.00053972
R203 x5[7].floating.n58 x5[7].floating.n57 0.00053972
R204 x5[7].floating.n46 x5[7].floating.n45 0.00053972
R205 x5[7].floating.n28 x5[7].floating.n27 0.00053972
R206 x5[7].floating.n16 x5[7].floating.n15 0.00053972
R207 x5[7].floating.n146 x5[7].floating.n145 0.00053972
R208 x5[7].floating.n158 x5[7].floating.n157 0.00053972
R209 x5[7].floating.n113 x5[7].floating.n112 0.00053972
R210 VDD.n1717 VDD.n4 426
R211 VDD.n1741 VDD.n2 351
R212 VDD.t9 VDD.n3 258.856
R213 VDD VDD.n1715 242.981
R214 VDD.n707 VDD.n119 198.118
R215 VDD.n530 VDD.n130 198.118
R216 VDD.n353 VDD.n141 198.118
R217 VDD.n997 VDD.n996 198.118
R218 VDD.n352 VDD.n142 198.118
R219 VDD.n529 VDD.n131 198.118
R220 VDD.n706 VDD.n120 198.118
R221 VDD.t12 VDD.n1739 188.965
R222 VDD.n892 VDD.n891 185
R223 VDD.n1053 VDD.n879 185
R224 VDD.n922 VDD.n920 185
R225 VDD.n1032 VDD.n918 185
R226 VDD.n1002 VDD.n1000 185
R227 VDD.n1052 VDD.n1051 185
R228 VDD.n1052 VDD.n108 185
R229 VDD.n931 VDD.n930 185
R230 VDD.n931 VDD.n108 185
R231 VDD.n1031 VDD.n1030 185
R232 VDD.n1031 VDD.n108 185
R233 VDD.n1011 VDD.n1010 185
R234 VDD.n998 VDD.n957 185
R235 VDD.n884 VDD.n883 185
R236 VDD.n179 VDD.n72 185
R237 VDD.n151 VDD.n149 185
R238 VDD.n227 VDD.n226 185
R239 VDD.n1664 VDD.n236 185
R240 VDD.n254 VDD.n237 185
R241 VDD.n1639 VDD.n1638 185
R242 VDD.n1641 VDD.n1640 185
R243 VDD.n1611 VDD.n1610 185
R244 VDD.n1620 VDD.n1619 185
R245 VDD.n1605 VDD.n1604 185
R246 VDD.n1607 VDD.n1606 185
R247 VDD.n1577 VDD.n1576 185
R248 VDD.n1586 VDD.n1585 185
R249 VDD.n1571 VDD.n1570 185
R250 VDD.n1573 VDD.n1572 185
R251 VDD.n351 VDD.n350 185
R252 VDD.n370 VDD.n369 185
R253 VDD.n386 VDD.n385 185
R254 VDD.n402 VDD.n401 185
R255 VDD.n1501 VDD.n417 185
R256 VDD.n431 VDD.n418 185
R257 VDD.n1476 VDD.n1475 185
R258 VDD.n1478 VDD.n1477 185
R259 VDD.n1448 VDD.n1447 185
R260 VDD.n1457 VDD.n1456 185
R261 VDD.n1442 VDD.n1441 185
R262 VDD.n1444 VDD.n1443 185
R263 VDD.n1414 VDD.n1413 185
R264 VDD.n1423 VDD.n1422 185
R265 VDD.n1408 VDD.n1407 185
R266 VDD.n1410 VDD.n1409 185
R267 VDD.n528 VDD.n527 185
R268 VDD.n547 VDD.n546 185
R269 VDD.n563 VDD.n562 185
R270 VDD.n579 VDD.n578 185
R271 VDD.n1338 VDD.n594 185
R272 VDD.n608 VDD.n595 185
R273 VDD.n1313 VDD.n1312 185
R274 VDD.n1315 VDD.n1314 185
R275 VDD.n1285 VDD.n1284 185
R276 VDD.n1294 VDD.n1293 185
R277 VDD.n1279 VDD.n1278 185
R278 VDD.n1281 VDD.n1280 185
R279 VDD.n1251 VDD.n1250 185
R280 VDD.n1260 VDD.n1259 185
R281 VDD.n1245 VDD.n1244 185
R282 VDD.n1247 VDD.n1246 185
R283 VDD.n705 VDD.n704 185
R284 VDD.n724 VDD.n723 185
R285 VDD.n740 VDD.n739 185
R286 VDD.n756 VDD.n755 185
R287 VDD.n1175 VDD.n771 185
R288 VDD.n785 VDD.n772 185
R289 VDD.n1150 VDD.n1149 185
R290 VDD.n1152 VDD.n1151 185
R291 VDD.n1122 VDD.n1121 185
R292 VDD.n1131 VDD.n1130 185
R293 VDD.n1116 VDD.n1115 185
R294 VDD.n1118 VDD.n1117 185
R295 VDD.n1088 VDD.n1087 185
R296 VDD.n1097 VDD.n1096 185
R297 VDD.n1082 VDD.n1081 185
R298 VDD.n1084 VDD.n1083 185
R299 VDD.n758 VDD.n757 185
R300 VDD.n742 VDD.n741 185
R301 VDD.n726 VDD.n725 185
R302 VDD.n711 VDD.n710 185
R303 VDD.n787 VDD.n786 185
R304 VDD.n709 VDD.n708 185
R305 VDD.n581 VDD.n580 185
R306 VDD.n565 VDD.n564 185
R307 VDD.n549 VDD.n548 185
R308 VDD.n534 VDD.n533 185
R309 VDD.n610 VDD.n609 185
R310 VDD.n532 VDD.n531 185
R311 VDD.n404 VDD.n403 185
R312 VDD.n388 VDD.n387 185
R313 VDD.n372 VDD.n371 185
R314 VDD.n357 VDD.n356 185
R315 VDD.n433 VDD.n432 185
R316 VDD.n355 VDD.n354 185
R317 VDD.n235 VDD.n234 185
R318 VDD.n225 VDD.n150 185
R319 VDD.n198 VDD.n197 185
R320 VDD.n256 VDD.n255 185
R321 VDD.n169 VDD.n168 185
R322 VDD.n1735 VDD.n2 185
R323 VDD.n1739 VDD.n2 185
R324 VDD.n1740 VDD 160.49
R325 VDD.n1743 VDD.t13 152.88
R326 VDD.n28 VDD.t10 152.879
R327 VDD.n1740 VDD.t12 113.897
R328 VDD.n1132 VDD.n1131 111.177
R329 VDD.n1098 VDD.n1097 111.177
R330 VDD.n710 VDD.n118 111.177
R331 VDD.n725 VDD.n100 111.177
R332 VDD.n741 VDD.n116 111.177
R333 VDD.n757 VDD.n102 111.177
R334 VDD.n1295 VDD.n1294 111.177
R335 VDD.n1261 VDD.n1260 111.177
R336 VDD.n533 VDD.n129 111.177
R337 VDD.n548 VDD.n91 111.177
R338 VDD.n564 VDD.n127 111.177
R339 VDD.n580 VDD.n93 111.177
R340 VDD.n1458 VDD.n1457 111.177
R341 VDD.n1424 VDD.n1423 111.177
R342 VDD.n356 VDD.n140 111.177
R343 VDD.n371 VDD.n82 111.177
R344 VDD.n387 VDD.n138 111.177
R345 VDD.n403 VDD.n84 111.177
R346 VDD.n1621 VDD.n1620 111.177
R347 VDD.n1587 VDD.n1586 111.177
R348 VDD.n197 VDD.n196 111.177
R349 VDD.n1687 VDD.n150 111.177
R350 VDD.n234 VDD.n75 111.177
R351 VDD.n1055 VDD.n892 111.177
R352 VDD.n1052 VDD.n893 111.177
R353 VDD.n1034 VDD.n931 111.177
R354 VDD.n1031 VDD.n932 111.177
R355 VDD.n1716 VDD.t9 108.719
R356 VDD.n1742 VDD.n1741 92.5005
R357 VDD.n1741 VDD.n1740 92.5005
R358 VDD.n1718 VDD.n1717 92.5005
R359 VDD.n1717 VDD.n1716 92.5005
R360 VDD.n1737 VDD.n1736 92.5005
R361 VDD.n1738 VDD.n1737 92.5005
R362 VDD.n880 VDD.n108 85.9427
R363 VDD.n997 VDD.n108 85.9427
R364 VDD.n1688 VDD.n74 85.9427
R365 VDD.n1688 VDD.n148 85.9427
R366 VDD.n1688 VDD.n76 85.9427
R367 VDD.n1688 VDD.n146 85.9427
R368 VDD.n1688 VDD.n144 85.9427
R369 VDD.n1688 VDD.n142 85.9427
R370 VDD.n1688 VDD.n141 85.9427
R371 VDD.n1688 VDD.n139 85.9427
R372 VDD.n1688 VDD.n83 85.9427
R373 VDD.n1688 VDD.n137 85.9427
R374 VDD.n1688 VDD.n85 85.9427
R375 VDD.n1688 VDD.n135 85.9427
R376 VDD.n1688 VDD.n133 85.9427
R377 VDD.n1688 VDD.n131 85.9427
R378 VDD.n1688 VDD.n130 85.9427
R379 VDD.n1688 VDD.n128 85.9427
R380 VDD.n1688 VDD.n92 85.9427
R381 VDD.n1688 VDD.n126 85.9427
R382 VDD.n1688 VDD.n94 85.9427
R383 VDD.n1688 VDD.n124 85.9427
R384 VDD.n1688 VDD.n122 85.9427
R385 VDD.n1688 VDD.n120 85.9427
R386 VDD.n1688 VDD.n119 85.9427
R387 VDD.n1688 VDD.n117 85.9427
R388 VDD.n1688 VDD.n101 85.9427
R389 VDD.n1688 VDD.n115 85.9427
R390 VDD.n1688 VDD.n103 85.9427
R391 VDD.n1688 VDD.n113 85.9427
R392 VDD.n1688 VDD.n111 85.9427
R393 VDD.n1716 VDD 77.6572
R394 VDD.n45 VDD.t1 70.3649
R395 VDD.n977 VDD.t6 68.0287
R396 VDD.n1689 VDD.n72 67.5405
R397 VDD.n1082 VDD.n109 67.5405
R398 VDD.n785 VDD.n104 67.3307
R399 VDD.n608 VDD.n95 67.3307
R400 VDD.n431 VDD.n86 67.3307
R401 VDD.n254 VDD.n77 67.3307
R402 VDD.n1012 VDD.n1011 67.3307
R403 VDD.n1639 VDD.n79 67.3307
R404 VDD.n1605 VDD.n80 67.3307
R405 VDD.n1571 VDD.n81 67.3307
R406 VDD.n1476 VDD.n88 67.3307
R407 VDD.n1442 VDD.n89 67.3307
R408 VDD.n1408 VDD.n90 67.3307
R409 VDD.n1313 VDD.n97 67.3307
R410 VDD.n1279 VDD.n98 67.3307
R411 VDD.n1245 VDD.n99 67.3307
R412 VDD.n1150 VDD.n106 67.3307
R413 VDD.n1116 VDD.n107 67.3307
R414 VDD.t14 VDD.t0 47.6077
R415 VDD.n38 VDD.t15 47.1434
R416 VDD.n38 VDD.t3 47.1434
R417 VDD.n1737 VDD.n2 39.0005
R418 VDD.n353 VDD.n352 33.746
R419 VDD.n530 VDD.n529 33.746
R420 VDD.n707 VDD.n706 33.746
R421 VDD.n1739 VDD.n1738 33.6517
R422 VDD.n1650 VDD.n257 32.9702
R423 VDD.n1487 VDD.n434 32.9702
R424 VDD.n1324 VDD.n611 32.9702
R425 VDD.n1161 VDD.n788 32.9702
R426 VDD.n995 VDD.n994 29.4128
R427 VDD.n1151 VDD.n1150 28.2358
R428 VDD.n1117 VDD.n1116 28.2358
R429 VDD.n1083 VDD.n1082 28.2358
R430 VDD.n786 VDD.n785 28.2358
R431 VDD.n1314 VDD.n1313 28.2358
R432 VDD.n1280 VDD.n1279 28.2358
R433 VDD.n1246 VDD.n1245 28.2358
R434 VDD.n609 VDD.n608 28.2358
R435 VDD.n1477 VDD.n1476 28.2358
R436 VDD.n1443 VDD.n1442 28.2358
R437 VDD.n1409 VDD.n1408 28.2358
R438 VDD.n432 VDD.n431 28.2358
R439 VDD.n1640 VDD.n1639 28.2358
R440 VDD.n1606 VDD.n1605 28.2358
R441 VDD.n1572 VDD.n1571 28.2358
R442 VDD.n168 VDD.n72 28.2358
R443 VDD.n255 VDD.n254 28.2358
R444 VDD.n1053 VDD.n1052 28.2358
R445 VDD.n931 VDD.n920 28.2358
R446 VDD.n1032 VDD.n1031 28.2358
R447 VDD.n1011 VDD.n1000 28.2358
R448 VDD.n1721 VDD.n1720 27.3454
R449 VDD.n1735 VDD.n1 22.8875
R450 VDD.t0 VDD.t2 21.1252
R451 VDD.n981 VDD.n980 20.7428
R452 VDD.n993 VDD.n984 20.7428
R453 VDD.n992 VDD.n987 20.7428
R454 VDD.n991 VDD.n990 20.7428
R455 VDD.n1713 VDD.n1712 20.7428
R456 VDD.n993 VDD.t4 18.5229
R457 VDD.t8 VDD 16.5329
R458 VDD.n992 VDD.t7 16.3798
R459 VDD.n1744 VDD.n1743 15.4666
R460 VDD.n28 VDD 15.1421
R461 VDD.n995 VDD.n977 13.3673
R462 VDD.n1121 VDD.n113 13.1177
R463 VDD.n1087 VDD.n111 13.1177
R464 VDD.n723 VDD.n117 13.1177
R465 VDD.n739 VDD.n101 13.1177
R466 VDD.n755 VDD.n115 13.1177
R467 VDD.n1175 VDD.n103 13.1177
R468 VDD.n1284 VDD.n124 13.1177
R469 VDD.n1250 VDD.n122 13.1177
R470 VDD.n704 VDD.n120 13.1177
R471 VDD.n546 VDD.n128 13.1177
R472 VDD.n562 VDD.n92 13.1177
R473 VDD.n578 VDD.n126 13.1177
R474 VDD.n1338 VDD.n94 13.1177
R475 VDD.n1447 VDD.n135 13.1177
R476 VDD.n1413 VDD.n133 13.1177
R477 VDD.n527 VDD.n131 13.1177
R478 VDD.n369 VDD.n139 13.1177
R479 VDD.n385 VDD.n83 13.1177
R480 VDD.n401 VDD.n137 13.1177
R481 VDD.n1501 VDD.n85 13.1177
R482 VDD.n1610 VDD.n146 13.1177
R483 VDD.n1576 VDD.n144 13.1177
R484 VDD.n350 VDD.n142 13.1177
R485 VDD.n149 VDD.n74 13.1177
R486 VDD.n226 VDD.n148 13.1177
R487 VDD.n1664 VDD.n76 13.1177
R488 VDD.n892 VDD.n880 13.1177
R489 VDD.n998 VDD.n997 13.1177
R490 VDD.n883 VDD.n880 13.1177
R491 VDD.n1620 VDD.n146 13.1177
R492 VDD.n1586 VDD.n144 13.1177
R493 VDD.n1457 VDD.n135 13.1177
R494 VDD.n1423 VDD.n133 13.1177
R495 VDD.n1294 VDD.n124 13.1177
R496 VDD.n1260 VDD.n122 13.1177
R497 VDD.n1131 VDD.n113 13.1177
R498 VDD.n1097 VDD.n111 13.1177
R499 VDD.n757 VDD.n103 13.1177
R500 VDD.n741 VDD.n115 13.1177
R501 VDD.n725 VDD.n101 13.1177
R502 VDD.n710 VDD.n117 13.1177
R503 VDD.n708 VDD.n119 13.1177
R504 VDD.n580 VDD.n94 13.1177
R505 VDD.n564 VDD.n126 13.1177
R506 VDD.n548 VDD.n92 13.1177
R507 VDD.n533 VDD.n128 13.1177
R508 VDD.n531 VDD.n130 13.1177
R509 VDD.n403 VDD.n85 13.1177
R510 VDD.n387 VDD.n137 13.1177
R511 VDD.n371 VDD.n83 13.1177
R512 VDD.n356 VDD.n139 13.1177
R513 VDD.n354 VDD.n141 13.1177
R514 VDD.n234 VDD.n76 13.1177
R515 VDD.n150 VDD.n148 13.1177
R516 VDD.n197 VDD.n74 13.1177
R517 VDD.n1713 VDD.t16 12.5529
R518 VDD.n1737 VDD.n4 12.0005
R519 VDD.n1742 VDD.n1 11.9758
R520 VDD.n852 VDD.n109 11.5452
R521 VDD.n1690 VDD.n1689 11.5452
R522 VDD.n991 VDD.t16 11.4813
R523 VDD.n1721 VDD.n1718 11.2229
R524 VDD.n1738 VDD.n3 10.3547
R525 VDD.t7 VDD.n991 9.64439
R526 VDD.n1153 VDD.n114 9.38471
R527 VDD.n1163 VDD.n105 9.38471
R528 VDD.n1316 VDD.n125 9.38471
R529 VDD.n1326 VDD.n96 9.38471
R530 VDD.n1479 VDD.n136 9.38471
R531 VDD.n1489 VDD.n87 9.38471
R532 VDD.n1642 VDD.n147 9.38471
R533 VDD.n1652 VDD.n78 9.38471
R534 VDD.n1650 VDD.n1649 9.3005
R535 VDD.n1569 VDD.n1568 9.3005
R536 VDD.n1603 VDD.n1602 9.3005
R537 VDD.n1637 VDD.n1636 9.3005
R538 VDD.n260 VDD.n257 9.3005
R539 VDD.n1618 VDD.n1617 9.3005
R540 VDD.n1584 VDD.n1583 9.3005
R541 VDD.n1487 VDD.n1486 9.3005
R542 VDD.n1406 VDD.n1405 9.3005
R543 VDD.n1440 VDD.n1439 9.3005
R544 VDD.n1474 VDD.n1473 9.3005
R545 VDD.n437 VDD.n434 9.3005
R546 VDD.n1455 VDD.n1454 9.3005
R547 VDD.n1421 VDD.n1420 9.3005
R548 VDD.n1324 VDD.n1323 9.3005
R549 VDD.n1243 VDD.n1242 9.3005
R550 VDD.n1277 VDD.n1276 9.3005
R551 VDD.n1311 VDD.n1310 9.3005
R552 VDD.n614 VDD.n611 9.3005
R553 VDD.n1292 VDD.n1291 9.3005
R554 VDD.n1258 VDD.n1257 9.3005
R555 VDD.n1161 VDD.n1160 9.3005
R556 VDD.n1080 VDD.n1079 9.3005
R557 VDD.n1114 VDD.n1113 9.3005
R558 VDD.n1148 VDD.n1147 9.3005
R559 VDD.n791 VDD.n788 9.3005
R560 VDD.n1129 VDD.n1128 9.3005
R561 VDD.n1095 VDD.n1094 9.3005
R562 VDD.n1173 VDD.n1172 9.3005
R563 VDD.n1187 VDD.n1186 9.3005
R564 VDD.n1199 VDD.n1198 9.3005
R565 VDD.n1211 VDD.n1210 9.3005
R566 VDD.n1223 VDD.n1222 9.3005
R567 VDD.n1336 VDD.n1335 9.3005
R568 VDD.n1350 VDD.n1349 9.3005
R569 VDD.n1362 VDD.n1361 9.3005
R570 VDD.n1374 VDD.n1373 9.3005
R571 VDD.n1386 VDD.n1385 9.3005
R572 VDD.n1499 VDD.n1498 9.3005
R573 VDD.n1513 VDD.n1512 9.3005
R574 VDD.n1525 VDD.n1524 9.3005
R575 VDD.n1537 VDD.n1536 9.3005
R576 VDD.n1549 VDD.n1548 9.3005
R577 VDD.n1662 VDD.n1661 9.3005
R578 VDD.n233 VDD.n232 9.3005
R579 VDD.n224 VDD.n155 9.3005
R580 VDD.n181 VDD.n180 9.3005
R581 VDD.n200 VDD.n199 9.3005
R582 VDD.n890 VDD.n889 9.3005
R583 VDD.n1050 VDD.n1049 9.3005
R584 VDD.n929 VDD.n928 9.3005
R585 VDD.n1029 VDD.n1028 9.3005
R586 VDD.n1009 VDD.n1008 9.3005
R587 VDD.n1057 VDD.n1056 9.3005
R588 VDD.n1056 VDD.n1055 9.3005
R589 VDD.n921 VDD.n896 9.3005
R590 VDD.n921 VDD.n893 9.3005
R591 VDD.n1036 VDD.n1035 9.3005
R592 VDD.n1035 VDD.n1034 9.3005
R593 VDD.n1001 VDD.n935 9.3005
R594 VDD.n1001 VDD.n932 9.3005
R595 VDD.n1015 VDD.n1014 9.3005
R596 VDD.n1014 VDD.n1013 9.3005
R597 VDD.n882 VDD.n881 9.3005
R598 VDD.n882 VDD.n108 9.3005
R599 VDD.n348 VDD.n321 9.3005
R600 VDD.n349 VDD.n348 9.3005
R601 VDD.n1574 VDD.n297 9.3005
R602 VDD.n1575 VDD.n1574 9.3005
R603 VDD.n1608 VDD.n264 9.3005
R604 VDD.n1609 VDD.n1608 9.3005
R605 VDD.n1642 VDD.n261 9.3005
R606 VDD.n1623 VDD.n1622 9.3005
R607 VDD.n1622 VDD.n1621 9.3005
R608 VDD.n1589 VDD.n1588 9.3005
R609 VDD.n1588 VDD.n1587 9.3005
R610 VDD.n525 VDD.n498 9.3005
R611 VDD.n526 VDD.n525 9.3005
R612 VDD.n1411 VDD.n474 9.3005
R613 VDD.n1412 VDD.n1411 9.3005
R614 VDD.n1445 VDD.n441 9.3005
R615 VDD.n1446 VDD.n1445 9.3005
R616 VDD.n1479 VDD.n438 9.3005
R617 VDD.n1460 VDD.n1459 9.3005
R618 VDD.n1459 VDD.n1458 9.3005
R619 VDD.n1426 VDD.n1425 9.3005
R620 VDD.n1425 VDD.n1424 9.3005
R621 VDD.n702 VDD.n675 9.3005
R622 VDD.n703 VDD.n702 9.3005
R623 VDD.n1248 VDD.n651 9.3005
R624 VDD.n1249 VDD.n1248 9.3005
R625 VDD.n1282 VDD.n618 9.3005
R626 VDD.n1283 VDD.n1282 9.3005
R627 VDD.n1316 VDD.n615 9.3005
R628 VDD.n1297 VDD.n1296 9.3005
R629 VDD.n1296 VDD.n1295 9.3005
R630 VDD.n1263 VDD.n1262 9.3005
R631 VDD.n1262 VDD.n1261 9.3005
R632 VDD.n1085 VDD.n828 9.3005
R633 VDD.n1086 VDD.n1085 9.3005
R634 VDD.n1119 VDD.n795 9.3005
R635 VDD.n1120 VDD.n1119 9.3005
R636 VDD.n1153 VDD.n792 9.3005
R637 VDD.n1134 VDD.n1133 9.3005
R638 VDD.n1133 VDD.n1132 9.3005
R639 VDD.n1100 VDD.n1099 9.3005
R640 VDD.n1099 VDD.n1098 9.3005
R641 VDD.n853 VDD.n852 9.3005
R642 VDD.n1178 VDD.n1177 9.3005
R643 VDD.n1177 VDD.n1176 9.3005
R644 VDD.n1190 VDD.n1189 9.3005
R645 VDD.n1189 VDD.n102 9.3005
R646 VDD.n1688 VDD.n102 9.3005
R647 VDD.n1202 VDD.n1201 9.3005
R648 VDD.n1201 VDD.n116 9.3005
R649 VDD.n1688 VDD.n116 9.3005
R650 VDD.n1214 VDD.n1213 9.3005
R651 VDD.n1213 VDD.n100 9.3005
R652 VDD.n1688 VDD.n100 9.3005
R653 VDD.n1164 VDD.n1163 9.3005
R654 VDD.n1226 VDD.n1225 9.3005
R655 VDD.n1225 VDD.n118 9.3005
R656 VDD.n1688 VDD.n118 9.3005
R657 VDD.n1341 VDD.n1340 9.3005
R658 VDD.n1340 VDD.n1339 9.3005
R659 VDD.n1353 VDD.n1352 9.3005
R660 VDD.n1352 VDD.n93 9.3005
R661 VDD.n1688 VDD.n93 9.3005
R662 VDD.n1365 VDD.n1364 9.3005
R663 VDD.n1364 VDD.n127 9.3005
R664 VDD.n1688 VDD.n127 9.3005
R665 VDD.n1377 VDD.n1376 9.3005
R666 VDD.n1376 VDD.n91 9.3005
R667 VDD.n1688 VDD.n91 9.3005
R668 VDD.n1327 VDD.n1326 9.3005
R669 VDD.n1389 VDD.n1388 9.3005
R670 VDD.n1388 VDD.n129 9.3005
R671 VDD.n1688 VDD.n129 9.3005
R672 VDD.n1504 VDD.n1503 9.3005
R673 VDD.n1503 VDD.n1502 9.3005
R674 VDD.n1516 VDD.n1515 9.3005
R675 VDD.n1515 VDD.n84 9.3005
R676 VDD.n1688 VDD.n84 9.3005
R677 VDD.n1528 VDD.n1527 9.3005
R678 VDD.n1527 VDD.n138 9.3005
R679 VDD.n1688 VDD.n138 9.3005
R680 VDD.n1540 VDD.n1539 9.3005
R681 VDD.n1539 VDD.n82 9.3005
R682 VDD.n1688 VDD.n82 9.3005
R683 VDD.n1490 VDD.n1489 9.3005
R684 VDD.n1552 VDD.n1551 9.3005
R685 VDD.n1551 VDD.n140 9.3005
R686 VDD.n1688 VDD.n140 9.3005
R687 VDD.n1667 VDD.n1666 9.3005
R688 VDD.n1666 VDD.n1665 9.3005
R689 VDD.n228 VDD.n157 9.3005
R690 VDD.n228 VDD.n75 9.3005
R691 VDD.n1688 VDD.n75 9.3005
R692 VDD.n1686 VDD.n1685 9.3005
R693 VDD.n1687 VDD.n1686 9.3005
R694 VDD.n1688 VDD.n1687 9.3005
R695 VDD.n1653 VDD.n1652 9.3005
R696 VDD.n1691 VDD.n1690 9.3005
R697 VDD.n195 VDD.n194 9.3005
R698 VDD.n196 VDD.n195 9.3005
R699 VDD.n1720 VDD.n1719 9.3005
R700 VDD.n1734 VDD.n1733 9.3005
R701 VDD.n1734 VDD.n4 9.3005
R702 VDD.n4 VDD.n3 9.3005
R703 VDD.n180 VDD.n179 8.92171
R704 VDD.n199 VDD.n198 8.92171
R705 VDD.n225 VDD.n224 8.92171
R706 VDD.n235 VDD.n233 8.92171
R707 VDD.n1662 VDD.n237 8.92171
R708 VDD.n1638 VDD.n1637 8.92171
R709 VDD.n1619 VDD.n1618 8.92171
R710 VDD.n1604 VDD.n1603 8.92171
R711 VDD.n1585 VDD.n1584 8.92171
R712 VDD.n1570 VDD.n1569 8.92171
R713 VDD.n1549 VDD.n357 8.92171
R714 VDD.n1537 VDD.n372 8.92171
R715 VDD.n1525 VDD.n388 8.92171
R716 VDD.n1513 VDD.n404 8.92171
R717 VDD.n1499 VDD.n418 8.92171
R718 VDD.n1475 VDD.n1474 8.92171
R719 VDD.n1456 VDD.n1455 8.92171
R720 VDD.n1441 VDD.n1440 8.92171
R721 VDD.n1422 VDD.n1421 8.92171
R722 VDD.n1407 VDD.n1406 8.92171
R723 VDD.n1386 VDD.n534 8.92171
R724 VDD.n1374 VDD.n549 8.92171
R725 VDD.n1362 VDD.n565 8.92171
R726 VDD.n1350 VDD.n581 8.92171
R727 VDD.n1336 VDD.n595 8.92171
R728 VDD.n1312 VDD.n1311 8.92171
R729 VDD.n1293 VDD.n1292 8.92171
R730 VDD.n1278 VDD.n1277 8.92171
R731 VDD.n1259 VDD.n1258 8.92171
R732 VDD.n1244 VDD.n1243 8.92171
R733 VDD.n1223 VDD.n711 8.92171
R734 VDD.n1211 VDD.n726 8.92171
R735 VDD.n1199 VDD.n742 8.92171
R736 VDD.n1187 VDD.n758 8.92171
R737 VDD.n1173 VDD.n772 8.92171
R738 VDD.n1149 VDD.n1148 8.92171
R739 VDD.n1130 VDD.n1129 8.92171
R740 VDD.n1115 VDD.n1114 8.92171
R741 VDD.n1096 VDD.n1095 8.92171
R742 VDD.n1081 VDD.n1080 8.92171
R743 VDD.n891 VDD.n890 8.92171
R744 VDD.n1051 VDD.n1050 8.92171
R745 VDD.n930 VDD.n929 8.92171
R746 VDD.n1030 VDD.n1029 8.92171
R747 VDD.n1010 VDD.n1009 8.92171
R748 VDD.n1054 VDD.n108 8.77616
R749 VDD.n919 VDD.n108 8.77616
R750 VDD.n1033 VDD.n108 8.77616
R751 VDD.n999 VDD.n108 8.77616
R752 VDD.n1688 VDD.n147 8.77616
R753 VDD.n1688 VDD.n145 8.77616
R754 VDD.n1688 VDD.n143 8.77616
R755 VDD.n1688 VDD.n136 8.77616
R756 VDD.n1688 VDD.n134 8.77616
R757 VDD.n1688 VDD.n132 8.77616
R758 VDD.n1688 VDD.n125 8.77616
R759 VDD.n1688 VDD.n123 8.77616
R760 VDD.n1688 VDD.n121 8.77616
R761 VDD.n1688 VDD.n114 8.77616
R762 VDD.n1688 VDD.n112 8.77616
R763 VDD.n1688 VDD.n110 8.77616
R764 VDD.n1688 VDD.n105 8.77616
R765 VDD.n1688 VDD.n96 8.77616
R766 VDD.n1688 VDD.n87 8.77616
R767 VDD.n1688 VDD.n78 8.77616
R768 VDD.n1688 VDD.n73 8.77616
R769 VDD.n1012 VDD.n108 5.63319
R770 VDD.n1688 VDD.n77 5.63319
R771 VDD.n1688 VDD.n81 5.63319
R772 VDD.n1688 VDD.n80 5.63319
R773 VDD.n1688 VDD.n79 5.63319
R774 VDD.n1688 VDD.n86 5.63319
R775 VDD.n1688 VDD.n90 5.63319
R776 VDD.n1688 VDD.n89 5.63319
R777 VDD.n1688 VDD.n88 5.63319
R778 VDD.n1688 VDD.n95 5.63319
R779 VDD.n1688 VDD.n99 5.63319
R780 VDD.n1688 VDD.n98 5.63319
R781 VDD.n1688 VDD.n97 5.63319
R782 VDD.n1688 VDD.n104 5.63319
R783 VDD.n1688 VDD.n107 5.63319
R784 VDD.n1688 VDD.n106 5.63319
R785 VDD.n1689 VDD.n1688 5.1329
R786 VDD.n1688 VDD.n109 5.1329
R787 VDD.n1715 VDD.t14 5.05206
R788 VDD.t4 VDD.n992 4.74591
R789 VDD.n7 VDD.n1 4.6505
R790 VDD.n1722 VDD.n1721 4.6505
R791 VDD.n1692 VDD.n1691 4.54027
R792 VDD.n1069 VDD.n853 4.54027
R793 VDD.n40 VDD.n39 4.52882
R794 VDD.n178 VDD.n70 4.5005
R795 VDD.n71 VDD.n70 4.5005
R796 VDD.n183 VDD.n182 4.5005
R797 VDD.n202 VDD.n201 4.5005
R798 VDD.n1648 VDD.n1647 4.5005
R799 VDD.n240 VDD.n238 4.5005
R800 VDD.n346 VDD.n339 4.5005
R801 VDD.n345 VDD.n344 4.5005
R802 VDD.n322 VDD.n320 4.5005
R803 VDD.n1567 VDD.n1566 4.5005
R804 VDD.n1567 VDD.n319 4.5005
R805 VDD.n1579 VDD.n1578 4.5005
R806 VDD.n298 VDD.n296 4.5005
R807 VDD.n1601 VDD.n1600 4.5005
R808 VDD.n1601 VDD.n295 4.5005
R809 VDD.n1613 VDD.n1612 4.5005
R810 VDD.n265 VDD.n263 4.5005
R811 VDD.n1635 VDD.n1634 4.5005
R812 VDD.n1635 VDD.n262 4.5005
R813 VDD.n281 VDD.n280 4.5005
R814 VDD.n1646 VDD.n258 4.5005
R815 VDD.n1645 VDD.n1644 4.5005
R816 VDD.n1644 VDD.n1643 4.5005
R817 VDD.n305 VDD.n293 4.5005
R818 VDD.n1616 VDD.n1615 4.5005
R819 VDD.n292 VDD.n290 4.5005
R820 VDD.n294 VDD.n292 4.5005
R821 VDD.n329 VDD.n317 4.5005
R822 VDD.n1582 VDD.n1581 4.5005
R823 VDD.n316 VDD.n314 4.5005
R824 VDD.n318 VDD.n316 4.5005
R825 VDD.n1485 VDD.n1484 4.5005
R826 VDD.n420 VDD.n419 4.5005
R827 VDD.n523 VDD.n516 4.5005
R828 VDD.n522 VDD.n521 4.5005
R829 VDD.n499 VDD.n497 4.5005
R830 VDD.n1404 VDD.n1403 4.5005
R831 VDD.n1404 VDD.n496 4.5005
R832 VDD.n1416 VDD.n1415 4.5005
R833 VDD.n475 VDD.n473 4.5005
R834 VDD.n1438 VDD.n1437 4.5005
R835 VDD.n1438 VDD.n472 4.5005
R836 VDD.n1450 VDD.n1449 4.5005
R837 VDD.n442 VDD.n440 4.5005
R838 VDD.n1472 VDD.n1471 4.5005
R839 VDD.n1472 VDD.n439 4.5005
R840 VDD.n458 VDD.n457 4.5005
R841 VDD.n1483 VDD.n435 4.5005
R842 VDD.n1482 VDD.n1481 4.5005
R843 VDD.n1481 VDD.n1480 4.5005
R844 VDD.n482 VDD.n470 4.5005
R845 VDD.n1453 VDD.n1452 4.5005
R846 VDD.n469 VDD.n467 4.5005
R847 VDD.n471 VDD.n469 4.5005
R848 VDD.n506 VDD.n494 4.5005
R849 VDD.n1419 VDD.n1418 4.5005
R850 VDD.n493 VDD.n491 4.5005
R851 VDD.n495 VDD.n493 4.5005
R852 VDD.n1322 VDD.n1321 4.5005
R853 VDD.n597 VDD.n596 4.5005
R854 VDD.n700 VDD.n693 4.5005
R855 VDD.n699 VDD.n698 4.5005
R856 VDD.n676 VDD.n674 4.5005
R857 VDD.n1241 VDD.n1240 4.5005
R858 VDD.n1241 VDD.n673 4.5005
R859 VDD.n1253 VDD.n1252 4.5005
R860 VDD.n652 VDD.n650 4.5005
R861 VDD.n1275 VDD.n1274 4.5005
R862 VDD.n1275 VDD.n649 4.5005
R863 VDD.n1287 VDD.n1286 4.5005
R864 VDD.n619 VDD.n617 4.5005
R865 VDD.n1309 VDD.n1308 4.5005
R866 VDD.n1309 VDD.n616 4.5005
R867 VDD.n635 VDD.n634 4.5005
R868 VDD.n1320 VDD.n612 4.5005
R869 VDD.n1319 VDD.n1318 4.5005
R870 VDD.n1318 VDD.n1317 4.5005
R871 VDD.n659 VDD.n647 4.5005
R872 VDD.n1290 VDD.n1289 4.5005
R873 VDD.n646 VDD.n644 4.5005
R874 VDD.n648 VDD.n646 4.5005
R875 VDD.n683 VDD.n671 4.5005
R876 VDD.n1256 VDD.n1255 4.5005
R877 VDD.n670 VDD.n668 4.5005
R878 VDD.n672 VDD.n670 4.5005
R879 VDD.n1159 VDD.n1158 4.5005
R880 VDD.n774 VDD.n773 4.5005
R881 VDD.n854 VDD.n851 4.5005
R882 VDD.n1090 VDD.n1089 4.5005
R883 VDD.n829 VDD.n827 4.5005
R884 VDD.n1112 VDD.n1111 4.5005
R885 VDD.n1112 VDD.n826 4.5005
R886 VDD.n1124 VDD.n1123 4.5005
R887 VDD.n796 VDD.n794 4.5005
R888 VDD.n1146 VDD.n1145 4.5005
R889 VDD.n1146 VDD.n793 4.5005
R890 VDD.n812 VDD.n811 4.5005
R891 VDD.n1157 VDD.n789 4.5005
R892 VDD.n1156 VDD.n1155 4.5005
R893 VDD.n1155 VDD.n1154 4.5005
R894 VDD.n836 VDD.n824 4.5005
R895 VDD.n1127 VDD.n1126 4.5005
R896 VDD.n823 VDD.n821 4.5005
R897 VDD.n825 VDD.n823 4.5005
R898 VDD.n861 VDD.n848 4.5005
R899 VDD.n1093 VDD.n1092 4.5005
R900 VDD.n847 VDD.n845 4.5005
R901 VDD.n849 VDD.n847 4.5005
R902 VDD.n1078 VDD.n1077 4.5005
R903 VDD.n1078 VDD.n850 4.5005
R904 VDD.n713 VDD.n712 4.5005
R905 VDD.n1171 VDD.n1170 4.5005
R906 VDD.n760 VDD.n759 4.5005
R907 VDD.n770 VDD.n768 4.5005
R908 VDD.n1174 VDD.n770 4.5005
R909 VDD.n1185 VDD.n1184 4.5005
R910 VDD.n744 VDD.n743 4.5005
R911 VDD.n754 VDD.n752 4.5005
R912 VDD.n1188 VDD.n754 4.5005
R913 VDD.n1197 VDD.n1196 4.5005
R914 VDD.n728 VDD.n727 4.5005
R915 VDD.n738 VDD.n736 4.5005
R916 VDD.n1200 VDD.n738 4.5005
R917 VDD.n722 VDD.n720 4.5005
R918 VDD.n1212 VDD.n722 4.5005
R919 VDD.n1209 VDD.n1208 4.5005
R920 VDD.n784 VDD.n782 4.5005
R921 VDD.n1162 VDD.n784 4.5005
R922 VDD.n701 VDD.n694 4.5005
R923 VDD.n1224 VDD.n701 4.5005
R924 VDD.n1221 VDD.n1220 4.5005
R925 VDD.n536 VDD.n535 4.5005
R926 VDD.n1334 VDD.n1333 4.5005
R927 VDD.n583 VDD.n582 4.5005
R928 VDD.n593 VDD.n591 4.5005
R929 VDD.n1337 VDD.n593 4.5005
R930 VDD.n1348 VDD.n1347 4.5005
R931 VDD.n567 VDD.n566 4.5005
R932 VDD.n577 VDD.n575 4.5005
R933 VDD.n1351 VDD.n577 4.5005
R934 VDD.n1360 VDD.n1359 4.5005
R935 VDD.n551 VDD.n550 4.5005
R936 VDD.n561 VDD.n559 4.5005
R937 VDD.n1363 VDD.n561 4.5005
R938 VDD.n545 VDD.n543 4.5005
R939 VDD.n1375 VDD.n545 4.5005
R940 VDD.n1372 VDD.n1371 4.5005
R941 VDD.n607 VDD.n605 4.5005
R942 VDD.n1325 VDD.n607 4.5005
R943 VDD.n524 VDD.n517 4.5005
R944 VDD.n1387 VDD.n524 4.5005
R945 VDD.n1384 VDD.n1383 4.5005
R946 VDD.n359 VDD.n358 4.5005
R947 VDD.n1497 VDD.n1496 4.5005
R948 VDD.n406 VDD.n405 4.5005
R949 VDD.n416 VDD.n414 4.5005
R950 VDD.n1500 VDD.n416 4.5005
R951 VDD.n1511 VDD.n1510 4.5005
R952 VDD.n390 VDD.n389 4.5005
R953 VDD.n400 VDD.n398 4.5005
R954 VDD.n1514 VDD.n400 4.5005
R955 VDD.n1523 VDD.n1522 4.5005
R956 VDD.n374 VDD.n373 4.5005
R957 VDD.n384 VDD.n382 4.5005
R958 VDD.n1526 VDD.n384 4.5005
R959 VDD.n368 VDD.n366 4.5005
R960 VDD.n1538 VDD.n368 4.5005
R961 VDD.n1535 VDD.n1534 4.5005
R962 VDD.n430 VDD.n428 4.5005
R963 VDD.n1488 VDD.n430 4.5005
R964 VDD.n347 VDD.n340 4.5005
R965 VDD.n1550 VDD.n347 4.5005
R966 VDD.n1547 VDD.n1546 4.5005
R967 VDD.n204 VDD.n153 4.5005
R968 VDD.n1660 VDD.n1659 4.5005
R969 VDD.n1669 VDD.n1668 4.5005
R970 VDD.n239 VDD.n223 4.5005
R971 VDD.n1663 VDD.n223 4.5005
R972 VDD.n221 VDD.n219 4.5005
R973 VDD.n1680 VDD.n1679 4.5005
R974 VDD.n231 VDD.n230 4.5005
R975 VDD.n231 VDD.n229 4.5005
R976 VDD.n1684 VDD.n1683 4.5005
R977 VDD.n1684 VDD.n152 4.5005
R978 VDD.n1682 VDD.n1681 4.5005
R979 VDD.n253 VDD.n251 4.5005
R980 VDD.n1651 VDD.n253 4.5005
R981 VDD.n166 VDD.n165 4.5005
R982 VDD.n167 VDD.n166 4.5005
R983 VDD.n184 VDD.n170 4.5005
R984 VDD.n1007 VDD.n1006 4.5005
R985 VDD.n962 VDD.n955 4.5005
R986 VDD.n885 VDD.n870 4.5005
R987 VDD.n904 VDD.n877 4.5005
R988 VDD.n888 VDD.n887 4.5005
R989 VDD.n924 VDD.n923 4.5005
R990 VDD.n897 VDD.n895 4.5005
R991 VDD.n943 VDD.n916 4.5005
R992 VDD.n927 VDD.n926 4.5005
R993 VDD.n1004 VDD.n1003 4.5005
R994 VDD.n936 VDD.n934 4.5005
R995 VDD.n954 VDD.n952 4.5005
R996 VDD.n956 VDD.n954 4.5005
R997 VDD.n876 VDD.n874 4.5005
R998 VDD.n878 VDD.n876 4.5005
R999 VDD.n1048 VDD.n1047 4.5005
R1000 VDD.n1048 VDD.n894 4.5005
R1001 VDD.n915 VDD.n913 4.5005
R1002 VDD.n917 VDD.n915 4.5005
R1003 VDD.n1027 VDD.n1026 4.5005
R1004 VDD.n1027 VDD.n933 4.5005
R1005 VDD.n27 VDD.n26 4.5005
R1006 VDD.n9 VDD.n6 4.5005
R1007 VDD.n10 VDD.n8 4.5005
R1008 VDD VDD.n108 4.28667
R1009 VDD.n1715 VDD.n1713 3.52129
R1010 VDD.n1724 VDD.n25 3.46788
R1011 VDD.n20 VDD.n19 3.46651
R1012 VDD.n46 VDD.n45 3.46323
R1013 VDD.n41 VDD.n35 3.46321
R1014 VDD.n1711 VDD.n30 3.45407
R1015 VDD.n989 VDD.n53 3.45407
R1016 VDD.n986 VDD.n57 3.45407
R1017 VDD.n983 VDD.n61 3.45407
R1018 VDD.n979 VDD.n65 3.45407
R1019 VDD.n31 VDD.n29 3.45149
R1020 VDD.n988 VDD.n51 3.45149
R1021 VDD.n985 VDD.n55 3.45149
R1022 VDD.n982 VDD.n59 3.45149
R1023 VDD.n978 VDD.n63 3.45149
R1024 VDD.n1068 VDD.n1067 3.42985
R1025 VDD.n13 VDD.n10 3.4257
R1026 VDD.n974 VDD.n959 3.42443
R1027 VDD.n1693 VDD.n1692 3.42376
R1028 VDD.n1070 VDD.n1069 3.42376
R1029 VDD.n37 VDD.n34 3.41853
R1030 VDD.n26 VDD.n11 3.41388
R1031 VDD.n1071 VDD.n1070 3.41326
R1032 VDD.n1694 VDD.n1693 3.41257
R1033 VDD.n46 VDD.n32 3.41218
R1034 VDD.n1707 VDD.n30 3.41218
R1035 VDD.n53 VDD.n50 3.41218
R1036 VDD.n57 VDD.n54 3.41218
R1037 VDD.n61 VDD.n58 3.41218
R1038 VDD.n65 VDD.n62 3.41218
R1039 VDD.n36 VDD.n33 3.41162
R1040 VDD.n186 VDD.n185 3.4105
R1041 VDD.n193 VDD.n192 3.4105
R1042 VDD.n270 VDD.n259 3.4105
R1043 VDD.n1633 VDD.n1632 3.4105
R1044 VDD.n1625 VDD.n1624 3.4105
R1045 VDD.n1599 VDD.n1598 3.4105
R1046 VDD.n1591 VDD.n1590 3.4105
R1047 VDD.n1565 VDD.n1564 3.4105
R1048 VDD.n342 VDD.n336 3.4105
R1049 VDD.n447 VDD.n436 3.4105
R1050 VDD.n1470 VDD.n1469 3.4105
R1051 VDD.n1462 VDD.n1461 3.4105
R1052 VDD.n1436 VDD.n1435 3.4105
R1053 VDD.n1428 VDD.n1427 3.4105
R1054 VDD.n1402 VDD.n1401 3.4105
R1055 VDD.n519 VDD.n513 3.4105
R1056 VDD.n624 VDD.n613 3.4105
R1057 VDD.n1307 VDD.n1306 3.4105
R1058 VDD.n1299 VDD.n1298 3.4105
R1059 VDD.n1273 VDD.n1272 3.4105
R1060 VDD.n1265 VDD.n1264 3.4105
R1061 VDD.n1239 VDD.n1238 3.4105
R1062 VDD.n696 VDD.n690 3.4105
R1063 VDD.n801 VDD.n790 3.4105
R1064 VDD.n1144 VDD.n1143 3.4105
R1065 VDD.n1136 VDD.n1135 3.4105
R1066 VDD.n1110 VDD.n1109 3.4105
R1067 VDD.n1102 VDD.n1101 3.4105
R1068 VDD.n1076 VDD.n1075 3.4105
R1069 VDD.n863 VDD.n862 3.4105
R1070 VDD.n1091 VDD.n843 3.4105
R1071 VDD.n838 VDD.n837 3.4105
R1072 VDD.n1125 VDD.n819 3.4105
R1073 VDD.n814 VDD.n813 3.4105
R1074 VDD.n1179 VDD.n769 3.4105
R1075 VDD.n1183 VDD.n1182 3.4105
R1076 VDD.n1191 VDD.n753 3.4105
R1077 VDD.n1195 VDD.n1194 3.4105
R1078 VDD.n1203 VDD.n737 3.4105
R1079 VDD.n1207 VDD.n1206 3.4105
R1080 VDD.n1215 VDD.n721 3.4105
R1081 VDD.n1219 VDD.n1218 3.4105
R1082 VDD.n1169 VDD.n1168 3.4105
R1083 VDD.n1165 VDD.n783 3.4105
R1084 VDD.n1227 VDD.n695 3.4105
R1085 VDD.n697 VDD.n689 3.4105
R1086 VDD.n685 VDD.n684 3.4105
R1087 VDD.n1254 VDD.n666 3.4105
R1088 VDD.n661 VDD.n660 3.4105
R1089 VDD.n1288 VDD.n642 3.4105
R1090 VDD.n637 VDD.n636 3.4105
R1091 VDD.n1342 VDD.n592 3.4105
R1092 VDD.n1346 VDD.n1345 3.4105
R1093 VDD.n1354 VDD.n576 3.4105
R1094 VDD.n1358 VDD.n1357 3.4105
R1095 VDD.n1366 VDD.n560 3.4105
R1096 VDD.n1370 VDD.n1369 3.4105
R1097 VDD.n1378 VDD.n544 3.4105
R1098 VDD.n1382 VDD.n1381 3.4105
R1099 VDD.n1332 VDD.n1331 3.4105
R1100 VDD.n1328 VDD.n606 3.4105
R1101 VDD.n1390 VDD.n518 3.4105
R1102 VDD.n520 VDD.n512 3.4105
R1103 VDD.n508 VDD.n507 3.4105
R1104 VDD.n1417 VDD.n489 3.4105
R1105 VDD.n484 VDD.n483 3.4105
R1106 VDD.n1451 VDD.n465 3.4105
R1107 VDD.n460 VDD.n459 3.4105
R1108 VDD.n1505 VDD.n415 3.4105
R1109 VDD.n1509 VDD.n1508 3.4105
R1110 VDD.n1517 VDD.n399 3.4105
R1111 VDD.n1521 VDD.n1520 3.4105
R1112 VDD.n1529 VDD.n383 3.4105
R1113 VDD.n1533 VDD.n1532 3.4105
R1114 VDD.n1541 VDD.n367 3.4105
R1115 VDD.n1545 VDD.n1544 3.4105
R1116 VDD.n1495 VDD.n1494 3.4105
R1117 VDD.n1491 VDD.n429 3.4105
R1118 VDD.n1553 VDD.n341 3.4105
R1119 VDD.n343 VDD.n335 3.4105
R1120 VDD.n331 VDD.n330 3.4105
R1121 VDD.n1580 VDD.n312 3.4105
R1122 VDD.n307 VDD.n306 3.4105
R1123 VDD.n1614 VDD.n288 3.4105
R1124 VDD.n283 VDD.n282 3.4105
R1125 VDD.n246 VDD.n222 3.4105
R1126 VDD.n1671 VDD.n1670 3.4105
R1127 VDD.n217 VDD.n158 3.4105
R1128 VDD.n159 VDD.n156 3.4105
R1129 VDD.n212 VDD.n154 3.4105
R1130 VDD.n206 VDD.n205 3.4105
R1131 VDD.n1658 VDD.n1657 3.4105
R1132 VDD.n1654 VDD.n252 3.4105
R1133 VDD.n176 VDD.n69 3.4105
R1134 VDD.n37 VDD.n36 3.4105
R1135 VDD.n42 VDD.n41 3.4105
R1136 VDD.n1696 VDD.n1695 3.4105
R1137 VDD.n1697 VDD.n1696 3.4105
R1138 VDD.n1699 VDD.n1698 3.4105
R1139 VDD.n1700 VDD.n1699 3.4105
R1140 VDD.n1702 VDD.n1701 3.4105
R1141 VDD.n1703 VDD.n1702 3.4105
R1142 VDD.n1705 VDD.n1704 3.4105
R1143 VDD.n1706 VDD.n1705 3.4105
R1144 VDD.n1709 VDD.n1708 3.4105
R1145 VDD.n1709 VDD.n49 3.4105
R1146 VDD.n48 VDD.n47 3.4105
R1147 VDD.n47 VDD.n43 3.4105
R1148 VDD.n67 VDD.n66 3.4105
R1149 VDD.n177 VDD.n173 3.4105
R1150 VDD.n164 VDD.n163 3.4105
R1151 VDD.n866 VDD.n856 3.4105
R1152 VDD.n1072 VDD.n857 3.4105
R1153 VDD.n865 VDD.n864 3.4105
R1154 VDD.n1103 VDD.n842 3.4105
R1155 VDD.n860 VDD.n859 3.4105
R1156 VDD.n1105 VDD.n1104 3.4105
R1157 VDD.n841 VDD.n831 3.4105
R1158 VDD.n1106 VDD.n832 3.4105
R1159 VDD.n840 VDD.n839 3.4105
R1160 VDD.n1137 VDD.n818 3.4105
R1161 VDD.n835 VDD.n834 3.4105
R1162 VDD.n1139 VDD.n1138 3.4105
R1163 VDD.n817 VDD.n798 3.4105
R1164 VDD.n1140 VDD.n799 3.4105
R1165 VDD.n816 VDD.n815 3.4105
R1166 VDD.n806 VDD.n805 3.4105
R1167 VDD.n809 VDD.n800 3.4105
R1168 VDD.n733 VDD.n732 3.4105
R1169 VDD.n718 VDD.n714 3.4105
R1170 VDD.n1217 VDD.n719 3.4105
R1171 VDD.n749 VDD.n748 3.4105
R1172 VDD.n734 VDD.n729 3.4105
R1173 VDD.n1205 VDD.n735 3.4105
R1174 VDD.n765 VDD.n764 3.4105
R1175 VDD.n750 VDD.n745 3.4105
R1176 VDD.n1193 VDD.n751 3.4105
R1177 VDD.n779 VDD.n778 3.4105
R1178 VDD.n766 VDD.n761 3.4105
R1179 VDD.n1181 VDD.n767 3.4105
R1180 VDD.n804 VDD.n803 3.4105
R1181 VDD.n780 VDD.n775 3.4105
R1182 VDD.n1167 VDD.n781 3.4105
R1183 VDD.n717 VDD.n716 3.4105
R1184 VDD.n1232 VDD.n1231 3.4105
R1185 VDD.n1230 VDD.n1229 3.4105
R1186 VDD.n1234 VDD.n1233 3.4105
R1187 VDD.n688 VDD.n678 3.4105
R1188 VDD.n1235 VDD.n679 3.4105
R1189 VDD.n687 VDD.n686 3.4105
R1190 VDD.n1266 VDD.n665 3.4105
R1191 VDD.n682 VDD.n681 3.4105
R1192 VDD.n1268 VDD.n1267 3.4105
R1193 VDD.n664 VDD.n654 3.4105
R1194 VDD.n1269 VDD.n655 3.4105
R1195 VDD.n663 VDD.n662 3.4105
R1196 VDD.n1300 VDD.n641 3.4105
R1197 VDD.n658 VDD.n657 3.4105
R1198 VDD.n1302 VDD.n1301 3.4105
R1199 VDD.n640 VDD.n621 3.4105
R1200 VDD.n1303 VDD.n622 3.4105
R1201 VDD.n639 VDD.n638 3.4105
R1202 VDD.n629 VDD.n628 3.4105
R1203 VDD.n632 VDD.n623 3.4105
R1204 VDD.n556 VDD.n555 3.4105
R1205 VDD.n541 VDD.n537 3.4105
R1206 VDD.n1380 VDD.n542 3.4105
R1207 VDD.n572 VDD.n571 3.4105
R1208 VDD.n557 VDD.n552 3.4105
R1209 VDD.n1368 VDD.n558 3.4105
R1210 VDD.n588 VDD.n587 3.4105
R1211 VDD.n573 VDD.n568 3.4105
R1212 VDD.n1356 VDD.n574 3.4105
R1213 VDD.n602 VDD.n601 3.4105
R1214 VDD.n589 VDD.n584 3.4105
R1215 VDD.n1344 VDD.n590 3.4105
R1216 VDD.n627 VDD.n626 3.4105
R1217 VDD.n603 VDD.n598 3.4105
R1218 VDD.n1330 VDD.n604 3.4105
R1219 VDD.n540 VDD.n539 3.4105
R1220 VDD.n1395 VDD.n1394 3.4105
R1221 VDD.n1393 VDD.n1392 3.4105
R1222 VDD.n1397 VDD.n1396 3.4105
R1223 VDD.n511 VDD.n501 3.4105
R1224 VDD.n1398 VDD.n502 3.4105
R1225 VDD.n510 VDD.n509 3.4105
R1226 VDD.n1429 VDD.n488 3.4105
R1227 VDD.n505 VDD.n504 3.4105
R1228 VDD.n1431 VDD.n1430 3.4105
R1229 VDD.n487 VDD.n477 3.4105
R1230 VDD.n1432 VDD.n478 3.4105
R1231 VDD.n486 VDD.n485 3.4105
R1232 VDD.n1463 VDD.n464 3.4105
R1233 VDD.n481 VDD.n480 3.4105
R1234 VDD.n1465 VDD.n1464 3.4105
R1235 VDD.n463 VDD.n444 3.4105
R1236 VDD.n1466 VDD.n445 3.4105
R1237 VDD.n462 VDD.n461 3.4105
R1238 VDD.n452 VDD.n451 3.4105
R1239 VDD.n455 VDD.n446 3.4105
R1240 VDD.n379 VDD.n378 3.4105
R1241 VDD.n364 VDD.n360 3.4105
R1242 VDD.n1543 VDD.n365 3.4105
R1243 VDD.n395 VDD.n394 3.4105
R1244 VDD.n380 VDD.n375 3.4105
R1245 VDD.n1531 VDD.n381 3.4105
R1246 VDD.n411 VDD.n410 3.4105
R1247 VDD.n396 VDD.n391 3.4105
R1248 VDD.n1519 VDD.n397 3.4105
R1249 VDD.n425 VDD.n424 3.4105
R1250 VDD.n412 VDD.n407 3.4105
R1251 VDD.n1507 VDD.n413 3.4105
R1252 VDD.n450 VDD.n449 3.4105
R1253 VDD.n426 VDD.n421 3.4105
R1254 VDD.n1493 VDD.n427 3.4105
R1255 VDD.n363 VDD.n362 3.4105
R1256 VDD.n1558 VDD.n1557 3.4105
R1257 VDD.n1556 VDD.n1555 3.4105
R1258 VDD.n1560 VDD.n1559 3.4105
R1259 VDD.n334 VDD.n324 3.4105
R1260 VDD.n1561 VDD.n325 3.4105
R1261 VDD.n333 VDD.n332 3.4105
R1262 VDD.n1592 VDD.n311 3.4105
R1263 VDD.n328 VDD.n327 3.4105
R1264 VDD.n1594 VDD.n1593 3.4105
R1265 VDD.n310 VDD.n300 3.4105
R1266 VDD.n1595 VDD.n301 3.4105
R1267 VDD.n309 VDD.n308 3.4105
R1268 VDD.n1626 VDD.n287 3.4105
R1269 VDD.n304 VDD.n303 3.4105
R1270 VDD.n1628 VDD.n1627 3.4105
R1271 VDD.n286 VDD.n267 3.4105
R1272 VDD.n1629 VDD.n268 3.4105
R1273 VDD.n285 VDD.n284 3.4105
R1274 VDD.n275 VDD.n274 3.4105
R1275 VDD.n278 VDD.n269 3.4105
R1276 VDD.n213 VDD.n161 3.4105
R1277 VDD.n208 VDD.n207 3.4105
R1278 VDD.n209 VDD.n162 3.4105
R1279 VDD.n1674 VDD.n1673 3.4105
R1280 VDD.n215 VDD.n214 3.4105
R1281 VDD.n1677 VDD.n1676 3.4105
R1282 VDD.n248 VDD.n247 3.4105
R1283 VDD.n1672 VDD.n216 3.4105
R1284 VDD.n243 VDD.n218 3.4105
R1285 VDD.n273 VDD.n272 3.4105
R1286 VDD.n249 VDD.n241 3.4105
R1287 VDD.n1656 VDD.n250 3.4105
R1288 VDD.n189 VDD.n172 3.4105
R1289 VDD.n188 VDD.n187 3.4105
R1290 VDD.n969 VDD.n968 3.4105
R1291 VDD.n1018 VDD.n949 3.4105
R1292 VDD.n948 VDD.n938 3.4105
R1293 VDD.n1020 VDD.n1019 3.4105
R1294 VDD.n947 VDD.n946 3.4105
R1295 VDD.n1039 VDD.n910 3.4105
R1296 VDD.n909 VDD.n899 3.4105
R1297 VDD.n1041 VDD.n1040 3.4105
R1298 VDD.n908 VDD.n907 3.4105
R1299 VDD.n1060 VDD.n872 3.4105
R1300 VDD.n1062 VDD.n1061 3.4105
R1301 VDD.n971 VDD.n970 3.4105
R1302 VDD.n960 VDD.n958 3.4105
R1303 VDD.n964 VDD.n963 3.4105
R1304 VDD.n1021 VDD.n939 3.4105
R1305 VDD.n942 VDD.n941 3.4105
R1306 VDD.n1042 VDD.n900 3.4105
R1307 VDD.n903 VDD.n902 3.4105
R1308 VDD.n1067 VDD.n1066 3.4105
R1309 VDD.n886 VDD.n871 3.4105
R1310 VDD.n1005 VDD.n950 3.4105
R1311 VDD.n1025 VDD.n1024 3.4105
R1312 VDD.n945 VDD.n944 3.4105
R1313 VDD.n1038 VDD.n1037 3.4105
R1314 VDD.n925 VDD.n911 3.4105
R1315 VDD.n1046 VDD.n1045 3.4105
R1316 VDD.n906 VDD.n905 3.4105
R1317 VDD.n1059 VDD.n1058 3.4105
R1318 VDD.n1064 VDD.n1063 3.4105
R1319 VDD.n967 VDD.n966 3.4105
R1320 VDD.n1017 VDD.n1016 3.4105
R1321 VDD.n1728 VDD.n1727 3.4105
R1322 VDD.n16 VDD.n15 3.4105
R1323 VDD.n18 VDD.n17 3.4105
R1324 VDD.n1726 VDD.n23 3.4105
R1325 VDD.n22 VDD.n21 3.4105
R1326 VDD.n1730 VDD.n1729 3.4105
R1327 VDD.n24 VDD.n22 3.4105
R1328 VDD.n1120 VDD.n106 3.38568
R1329 VDD.n1086 VDD.n107 3.38568
R1330 VDD.n1283 VDD.n97 3.38568
R1331 VDD.n1249 VDD.n98 3.38568
R1332 VDD.n703 VDD.n99 3.38568
R1333 VDD.n1446 VDD.n88 3.38568
R1334 VDD.n1412 VDD.n89 3.38568
R1335 VDD.n526 VDD.n90 3.38568
R1336 VDD.n1609 VDD.n79 3.38568
R1337 VDD.n1575 VDD.n80 3.38568
R1338 VDD.n349 VDD.n81 3.38568
R1339 VDD.n1013 VDD.n1012 3.38568
R1340 VDD.n1176 VDD.n104 3.38568
R1341 VDD.n1339 VDD.n95 3.38568
R1342 VDD.n1502 VDD.n86 3.38568
R1343 VDD.n1665 VDD.n77 3.38568
R1344 VDD.n180 VDD.n71 3.10353
R1345 VDD.n179 VDD.n169 3.10353
R1346 VDD.n199 VDD.n167 3.10353
R1347 VDD.n198 VDD.n151 3.10353
R1348 VDD.n224 VDD.n152 3.10353
R1349 VDD.n227 VDD.n225 3.10353
R1350 VDD.n233 VDD.n229 3.10353
R1351 VDD.n236 VDD.n235 3.10353
R1352 VDD.n1663 VDD.n1662 3.10353
R1353 VDD.n256 VDD.n237 3.10353
R1354 VDD.n1651 VDD.n1650 3.10353
R1355 VDD.n1643 VDD.n257 3.10353
R1356 VDD.n1641 VDD.n1638 3.10353
R1357 VDD.n1637 VDD.n262 3.10353
R1358 VDD.n1619 VDD.n1611 3.10353
R1359 VDD.n1618 VDD.n294 3.10353
R1360 VDD.n1607 VDD.n1604 3.10353
R1361 VDD.n1603 VDD.n295 3.10353
R1362 VDD.n1585 VDD.n1577 3.10353
R1363 VDD.n1584 VDD.n318 3.10353
R1364 VDD.n1573 VDD.n1570 3.10353
R1365 VDD.n1569 VDD.n319 3.10353
R1366 VDD.n352 VDD.n351 3.10353
R1367 VDD.n355 VDD.n353 3.10353
R1368 VDD.n1550 VDD.n1549 3.10353
R1369 VDD.n370 VDD.n357 3.10353
R1370 VDD.n1538 VDD.n1537 3.10353
R1371 VDD.n386 VDD.n372 3.10353
R1372 VDD.n1526 VDD.n1525 3.10353
R1373 VDD.n402 VDD.n388 3.10353
R1374 VDD.n1514 VDD.n1513 3.10353
R1375 VDD.n417 VDD.n404 3.10353
R1376 VDD.n1500 VDD.n1499 3.10353
R1377 VDD.n433 VDD.n418 3.10353
R1378 VDD.n1488 VDD.n1487 3.10353
R1379 VDD.n1480 VDD.n434 3.10353
R1380 VDD.n1478 VDD.n1475 3.10353
R1381 VDD.n1474 VDD.n439 3.10353
R1382 VDD.n1456 VDD.n1448 3.10353
R1383 VDD.n1455 VDD.n471 3.10353
R1384 VDD.n1444 VDD.n1441 3.10353
R1385 VDD.n1440 VDD.n472 3.10353
R1386 VDD.n1422 VDD.n1414 3.10353
R1387 VDD.n1421 VDD.n495 3.10353
R1388 VDD.n1410 VDD.n1407 3.10353
R1389 VDD.n1406 VDD.n496 3.10353
R1390 VDD.n529 VDD.n528 3.10353
R1391 VDD.n532 VDD.n530 3.10353
R1392 VDD.n1387 VDD.n1386 3.10353
R1393 VDD.n547 VDD.n534 3.10353
R1394 VDD.n1375 VDD.n1374 3.10353
R1395 VDD.n563 VDD.n549 3.10353
R1396 VDD.n1363 VDD.n1362 3.10353
R1397 VDD.n579 VDD.n565 3.10353
R1398 VDD.n1351 VDD.n1350 3.10353
R1399 VDD.n594 VDD.n581 3.10353
R1400 VDD.n1337 VDD.n1336 3.10353
R1401 VDD.n610 VDD.n595 3.10353
R1402 VDD.n1325 VDD.n1324 3.10353
R1403 VDD.n1317 VDD.n611 3.10353
R1404 VDD.n1315 VDD.n1312 3.10353
R1405 VDD.n1311 VDD.n616 3.10353
R1406 VDD.n1293 VDD.n1285 3.10353
R1407 VDD.n1292 VDD.n648 3.10353
R1408 VDD.n1281 VDD.n1278 3.10353
R1409 VDD.n1277 VDD.n649 3.10353
R1410 VDD.n1259 VDD.n1251 3.10353
R1411 VDD.n1258 VDD.n672 3.10353
R1412 VDD.n1247 VDD.n1244 3.10353
R1413 VDD.n1243 VDD.n673 3.10353
R1414 VDD.n706 VDD.n705 3.10353
R1415 VDD.n709 VDD.n707 3.10353
R1416 VDD.n1224 VDD.n1223 3.10353
R1417 VDD.n724 VDD.n711 3.10353
R1418 VDD.n1212 VDD.n1211 3.10353
R1419 VDD.n740 VDD.n726 3.10353
R1420 VDD.n1200 VDD.n1199 3.10353
R1421 VDD.n756 VDD.n742 3.10353
R1422 VDD.n1188 VDD.n1187 3.10353
R1423 VDD.n771 VDD.n758 3.10353
R1424 VDD.n1174 VDD.n1173 3.10353
R1425 VDD.n787 VDD.n772 3.10353
R1426 VDD.n1162 VDD.n1161 3.10353
R1427 VDD.n1154 VDD.n788 3.10353
R1428 VDD.n1152 VDD.n1149 3.10353
R1429 VDD.n1148 VDD.n793 3.10353
R1430 VDD.n1130 VDD.n1122 3.10353
R1431 VDD.n1129 VDD.n825 3.10353
R1432 VDD.n1118 VDD.n1115 3.10353
R1433 VDD.n1114 VDD.n826 3.10353
R1434 VDD.n1096 VDD.n1088 3.10353
R1435 VDD.n1095 VDD.n849 3.10353
R1436 VDD.n1084 VDD.n1081 3.10353
R1437 VDD.n1080 VDD.n850 3.10353
R1438 VDD.n891 VDD.n884 3.10353
R1439 VDD.n890 VDD.n878 3.10353
R1440 VDD.n1051 VDD.n879 3.10353
R1441 VDD.n1050 VDD.n894 3.10353
R1442 VDD.n930 VDD.n922 3.10353
R1443 VDD.n929 VDD.n917 3.10353
R1444 VDD.n1030 VDD.n918 3.10353
R1445 VDD.n1029 VDD.n933 3.10353
R1446 VDD.n1010 VDD.n1002 3.10353
R1447 VDD.n1009 VDD.n956 3.10353
R1448 VDD.n6 VDD.n5 3.03311
R1449 VDD VDD.n981 2.90898
R1450 VDD.n1736 VDD.n1735 2.64177
R1451 VDD.n881 VDD.n869 2.5429
R1452 VDD.n1720 VDD.n5 2.4386
R1453 VDD.n996 VDD.n957 2.28608
R1454 VDD.n1712 VDD.n29 2.24869
R1455 VDD.n990 VDD.n988 2.24869
R1456 VDD.n987 VDD.n985 2.24869
R1457 VDD.n984 VDD.n982 2.24869
R1458 VDD.n980 VDD.n978 2.24869
R1459 VDD.n996 VDD.n995 2.15377
R1460 VDD.n994 VDD.n993 1.99051
R1461 VDD.n976 VDD.n975 1.94045
R1462 VDD.n19 VDD.n0 1.94045
R1463 VDD.n1724 VDD.n1723 1.94045
R1464 VDD.n1121 VDD.n1120 1.76521
R1465 VDD.n1087 VDD.n1086 1.76521
R1466 VDD.n708 VDD.n118 1.76521
R1467 VDD.n723 VDD.n100 1.76521
R1468 VDD.n739 VDD.n116 1.76521
R1469 VDD.n755 VDD.n102 1.76521
R1470 VDD.n1176 VDD.n1175 1.76521
R1471 VDD.n1284 VDD.n1283 1.76521
R1472 VDD.n1250 VDD.n1249 1.76521
R1473 VDD.n704 VDD.n703 1.76521
R1474 VDD.n531 VDD.n129 1.76521
R1475 VDD.n546 VDD.n91 1.76521
R1476 VDD.n562 VDD.n127 1.76521
R1477 VDD.n578 VDD.n93 1.76521
R1478 VDD.n1339 VDD.n1338 1.76521
R1479 VDD.n1447 VDD.n1446 1.76521
R1480 VDD.n1413 VDD.n1412 1.76521
R1481 VDD.n527 VDD.n526 1.76521
R1482 VDD.n354 VDD.n140 1.76521
R1483 VDD.n369 VDD.n82 1.76521
R1484 VDD.n385 VDD.n138 1.76521
R1485 VDD.n401 VDD.n84 1.76521
R1486 VDD.n1502 VDD.n1501 1.76521
R1487 VDD.n1610 VDD.n1609 1.76521
R1488 VDD.n1576 VDD.n1575 1.76521
R1489 VDD.n350 VDD.n349 1.76521
R1490 VDD.n1687 VDD.n149 1.76521
R1491 VDD.n226 VDD.n75 1.76521
R1492 VDD.n1665 VDD.n1664 1.76521
R1493 VDD.n883 VDD.n882 1.76521
R1494 VDD.n1013 VDD.n998 1.76521
R1495 VDD.n981 VDD.t5 1.68435
R1496 VDD.n1054 VDD.n1053 1.66612
R1497 VDD.n920 VDD.n919 1.66612
R1498 VDD.n1033 VDD.n1032 1.66612
R1499 VDD.n1000 VDD.n999 1.66612
R1500 VDD.n1640 VDD.n147 1.66612
R1501 VDD.n1606 VDD.n145 1.66612
R1502 VDD.n1572 VDD.n143 1.66612
R1503 VDD.n1477 VDD.n136 1.66612
R1504 VDD.n1443 VDD.n134 1.66612
R1505 VDD.n1409 VDD.n132 1.66612
R1506 VDD.n1314 VDD.n125 1.66612
R1507 VDD.n1280 VDD.n123 1.66612
R1508 VDD.n1246 VDD.n121 1.66612
R1509 VDD.n1151 VDD.n114 1.66612
R1510 VDD.n1117 VDD.n112 1.66612
R1511 VDD.n1083 VDD.n110 1.66612
R1512 VDD.n786 VDD.n105 1.66612
R1513 VDD.n609 VDD.n96 1.66612
R1514 VDD.n432 VDD.n87 1.66612
R1515 VDD.n255 VDD.n78 1.66612
R1516 VDD.n168 VDD.n73 1.66612
R1517 VDD.n1016 VDD.n1015 1.35607
R1518 VDD.n194 VDD.n193 1.35607
R1519 VDD.n261 VDD.n259 1.35607
R1520 VDD.n1633 VDD.n264 1.35607
R1521 VDD.n1624 VDD.n1623 1.35607
R1522 VDD.n1599 VDD.n297 1.35607
R1523 VDD.n1590 VDD.n1589 1.35607
R1524 VDD.n1565 VDD.n321 1.35607
R1525 VDD.n438 VDD.n436 1.35607
R1526 VDD.n1470 VDD.n441 1.35607
R1527 VDD.n1461 VDD.n1460 1.35607
R1528 VDD.n1436 VDD.n474 1.35607
R1529 VDD.n1427 VDD.n1426 1.35607
R1530 VDD.n1402 VDD.n498 1.35607
R1531 VDD.n615 VDD.n613 1.35607
R1532 VDD.n1307 VDD.n618 1.35607
R1533 VDD.n1298 VDD.n1297 1.35607
R1534 VDD.n1273 VDD.n651 1.35607
R1535 VDD.n1264 VDD.n1263 1.35607
R1536 VDD.n1239 VDD.n675 1.35607
R1537 VDD.n792 VDD.n790 1.35607
R1538 VDD.n1144 VDD.n795 1.35607
R1539 VDD.n1135 VDD.n1134 1.35607
R1540 VDD.n1110 VDD.n828 1.35607
R1541 VDD.n1101 VDD.n1100 1.35607
R1542 VDD.n1076 VDD.n853 1.35607
R1543 VDD.n1179 VDD.n1178 1.35607
R1544 VDD.n1191 VDD.n1190 1.35607
R1545 VDD.n1203 VDD.n1202 1.35607
R1546 VDD.n1215 VDD.n1214 1.35607
R1547 VDD.n1165 VDD.n1164 1.35607
R1548 VDD.n1227 VDD.n1226 1.35607
R1549 VDD.n1342 VDD.n1341 1.35607
R1550 VDD.n1354 VDD.n1353 1.35607
R1551 VDD.n1366 VDD.n1365 1.35607
R1552 VDD.n1378 VDD.n1377 1.35607
R1553 VDD.n1328 VDD.n1327 1.35607
R1554 VDD.n1390 VDD.n1389 1.35607
R1555 VDD.n1505 VDD.n1504 1.35607
R1556 VDD.n1517 VDD.n1516 1.35607
R1557 VDD.n1529 VDD.n1528 1.35607
R1558 VDD.n1541 VDD.n1540 1.35607
R1559 VDD.n1491 VDD.n1490 1.35607
R1560 VDD.n1553 VDD.n1552 1.35607
R1561 VDD.n1667 VDD.n222 1.35607
R1562 VDD.n158 VDD.n157 1.35607
R1563 VDD.n1685 VDD.n154 1.35607
R1564 VDD.n1654 VDD.n1653 1.35607
R1565 VDD.n1691 VDD.n69 1.35607
R1566 VDD.n1025 VDD.n935 1.35607
R1567 VDD.n1037 VDD.n1036 1.35607
R1568 VDD.n1046 VDD.n896 1.35607
R1569 VDD.n1058 VDD.n1057 1.35607
R1570 VDD.n1732 VDD.n1731 1.35607
R1571 VDD.n44 VDD.n32 1.13981
R1572 VDD.n1074 VDD.n1073 1.13717
R1573 VDD.n68 VDD.n67 1.13717
R1574 VDD.n857 VDD.n855 1.13717
R1575 VDD.n858 VDD.n844 1.13717
R1576 VDD.n860 VDD.n846 1.13717
R1577 VDD.n1108 VDD.n1107 1.13717
R1578 VDD.n832 VDD.n830 1.13717
R1579 VDD.n833 VDD.n820 1.13717
R1580 VDD.n835 VDD.n822 1.13717
R1581 VDD.n1142 VDD.n1141 1.13717
R1582 VDD.n799 VDD.n797 1.13717
R1583 VDD.n808 VDD.n807 1.13717
R1584 VDD.n810 VDD.n809 1.13717
R1585 VDD.n731 VDD.n715 1.13717
R1586 VDD.n1217 VDD.n1216 1.13717
R1587 VDD.n747 VDD.n730 1.13717
R1588 VDD.n1205 VDD.n1204 1.13717
R1589 VDD.n763 VDD.n746 1.13717
R1590 VDD.n1193 VDD.n1192 1.13717
R1591 VDD.n777 VDD.n762 1.13717
R1592 VDD.n1181 VDD.n1180 1.13717
R1593 VDD.n802 VDD.n776 1.13717
R1594 VDD.n1167 VDD.n1166 1.13717
R1595 VDD.n692 VDD.n691 1.13717
R1596 VDD.n1229 VDD.n1228 1.13717
R1597 VDD.n1237 VDD.n1236 1.13717
R1598 VDD.n679 VDD.n677 1.13717
R1599 VDD.n680 VDD.n667 1.13717
R1600 VDD.n682 VDD.n669 1.13717
R1601 VDD.n1271 VDD.n1270 1.13717
R1602 VDD.n655 VDD.n653 1.13717
R1603 VDD.n656 VDD.n643 1.13717
R1604 VDD.n658 VDD.n645 1.13717
R1605 VDD.n1305 VDD.n1304 1.13717
R1606 VDD.n622 VDD.n620 1.13717
R1607 VDD.n631 VDD.n630 1.13717
R1608 VDD.n633 VDD.n632 1.13717
R1609 VDD.n554 VDD.n538 1.13717
R1610 VDD.n1380 VDD.n1379 1.13717
R1611 VDD.n570 VDD.n553 1.13717
R1612 VDD.n1368 VDD.n1367 1.13717
R1613 VDD.n586 VDD.n569 1.13717
R1614 VDD.n1356 VDD.n1355 1.13717
R1615 VDD.n600 VDD.n585 1.13717
R1616 VDD.n1344 VDD.n1343 1.13717
R1617 VDD.n625 VDD.n599 1.13717
R1618 VDD.n1330 VDD.n1329 1.13717
R1619 VDD.n515 VDD.n514 1.13717
R1620 VDD.n1392 VDD.n1391 1.13717
R1621 VDD.n1400 VDD.n1399 1.13717
R1622 VDD.n502 VDD.n500 1.13717
R1623 VDD.n503 VDD.n490 1.13717
R1624 VDD.n505 VDD.n492 1.13717
R1625 VDD.n1434 VDD.n1433 1.13717
R1626 VDD.n478 VDD.n476 1.13717
R1627 VDD.n479 VDD.n466 1.13717
R1628 VDD.n481 VDD.n468 1.13717
R1629 VDD.n1468 VDD.n1467 1.13717
R1630 VDD.n445 VDD.n443 1.13717
R1631 VDD.n454 VDD.n453 1.13717
R1632 VDD.n456 VDD.n455 1.13717
R1633 VDD.n377 VDD.n361 1.13717
R1634 VDD.n1543 VDD.n1542 1.13717
R1635 VDD.n393 VDD.n376 1.13717
R1636 VDD.n1531 VDD.n1530 1.13717
R1637 VDD.n409 VDD.n392 1.13717
R1638 VDD.n1519 VDD.n1518 1.13717
R1639 VDD.n423 VDD.n408 1.13717
R1640 VDD.n1507 VDD.n1506 1.13717
R1641 VDD.n448 VDD.n422 1.13717
R1642 VDD.n1493 VDD.n1492 1.13717
R1643 VDD.n338 VDD.n337 1.13717
R1644 VDD.n1555 VDD.n1554 1.13717
R1645 VDD.n1563 VDD.n1562 1.13717
R1646 VDD.n325 VDD.n323 1.13717
R1647 VDD.n326 VDD.n313 1.13717
R1648 VDD.n328 VDD.n315 1.13717
R1649 VDD.n1597 VDD.n1596 1.13717
R1650 VDD.n301 VDD.n299 1.13717
R1651 VDD.n302 VDD.n289 1.13717
R1652 VDD.n304 VDD.n291 1.13717
R1653 VDD.n1631 VDD.n1630 1.13717
R1654 VDD.n268 VDD.n266 1.13717
R1655 VDD.n277 VDD.n276 1.13717
R1656 VDD.n279 VDD.n278 1.13717
R1657 VDD.n211 VDD.n210 1.13717
R1658 VDD.n203 VDD.n162 1.13717
R1659 VDD.n1675 VDD.n160 1.13717
R1660 VDD.n1678 VDD.n1677 1.13717
R1661 VDD.n245 VDD.n244 1.13717
R1662 VDD.n220 VDD.n218 1.13717
R1663 VDD.n271 VDD.n242 1.13717
R1664 VDD.n1656 VDD.n1655 1.13717
R1665 VDD.n172 VDD.n171 1.13717
R1666 VDD.n191 VDD.n190 1.13717
R1667 VDD.n175 VDD.n174 1.13717
R1668 VDD.n965 VDD.n951 1.13717
R1669 VDD.n868 VDD.n867 1.13717
R1670 VDD.n901 VDD.n873 1.13717
R1671 VDD.n1044 VDD.n1043 1.13717
R1672 VDD.n940 VDD.n912 1.13717
R1673 VDD.n1023 VDD.n1022 1.13717
R1674 VDD.n939 VDD.n937 1.13717
R1675 VDD.n942 VDD.n914 1.13717
R1676 VDD.n900 VDD.n898 1.13717
R1677 VDD.n903 VDD.n875 1.13717
R1678 VDD.n1065 VDD.n1064 1.13717
R1679 VDD.n966 VDD.n953 1.13717
R1680 VDD.n1730 VDD.n12 1.13717
R1681 VDD.n63 VDD.n62 1.13462
R1682 VDD.n59 VDD.n58 1.13462
R1683 VDD.n55 VDD.n54 1.13462
R1684 VDD.n51 VDD.n50 1.13462
R1685 VDD.n1707 VDD.n31 1.13462
R1686 VDD.n41 VDD.n40 1.13005
R1687 VDD.n1712 VDD.n1711 1.04017
R1688 VDD.n990 VDD.n989 1.04017
R1689 VDD.n987 VDD.n986 1.04017
R1690 VDD.n984 VDD.n983 1.04017
R1691 VDD.n980 VDD.n979 1.04017
R1692 VDD.n1734 VDD.n5 1.01637
R1693 VDD.t5 VDD 0.918966
R1694 VDD.n25 VDD.n23 0.870766
R1695 VDD.n20 VDD.n18 0.870578
R1696 VDD.n34 VDD.n33 0.853291
R1697 VDD.n1696 VDD.n64 0.853
R1698 VDD.n1699 VDD.n60 0.853
R1699 VDD.n1702 VDD.n56 0.853
R1700 VDD.n1705 VDD.n52 0.853
R1701 VDD.n1710 VDD.n1709 0.853
R1702 VDD.n973 VDD.n972 0.853
R1703 VDD.n1731 VDD.n1730 0.853
R1704 VDD.n1066 VDD.n869 0.849366
R1705 VDD.n1718 VDD.n28 0.813198
R1706 VDD.n1736 VDD.n1734 0.813198
R1707 VDD.n45 VDD.n44 0.684595
R1708 VDD.n19 VDD.n14 0.682713
R1709 VDD.n1725 VDD.n1724 0.682713
R1710 VDD.n975 VDD.n974 0.682447
R1711 VDD.n994 VDD.t8 0.612811
R1712 VDD.n1688 VDD.n108 0.459733
R1713 VDD.t2 VDD.n1714 0.454532
R1714 VDD.n1714 VDD.t11 0.45205
R1715 VDD.n1743 VDD.n1742 0.406849
R1716 VDD.n43 VDD.n42 0.357419
R1717 VDD.n346 VDD.n345 0.314894
R1718 VDD.n523 VDD.n522 0.314894
R1719 VDD.n700 VDD.n699 0.314894
R1720 VDD.n1648 VDD.n258 0.30353
R1721 VDD.n1485 VDD.n435 0.30353
R1722 VDD.n1322 VDD.n612 0.30353
R1723 VDD.n1159 VDD.n789 0.30353
R1724 VDD.n1647 VDD.n1646 0.30353
R1725 VDD.n1484 VDD.n1483 0.30353
R1726 VDD.n1321 VDD.n1320 0.30353
R1727 VDD.n1158 VDD.n1157 0.30353
R1728 VDD.n343 VDD.n342 0.288379
R1729 VDD.n520 VDD.n519 0.288379
R1730 VDD.n697 VDD.n696 0.288379
R1731 VDD.n1690 VDD.n71 0.194439
R1732 VDD.n195 VDD.n169 0.194439
R1733 VDD.n195 VDD.n167 0.194439
R1734 VDD.n1686 VDD.n151 0.194439
R1735 VDD.n1686 VDD.n152 0.194439
R1736 VDD.n228 VDD.n227 0.194439
R1737 VDD.n229 VDD.n228 0.194439
R1738 VDD.n1666 VDD.n236 0.194439
R1739 VDD.n1666 VDD.n1663 0.194439
R1740 VDD.n1652 VDD.n256 0.194439
R1741 VDD.n1652 VDD.n1651 0.194439
R1742 VDD.n1643 VDD.n1642 0.194439
R1743 VDD.n1642 VDD.n1641 0.194439
R1744 VDD.n1608 VDD.n262 0.194439
R1745 VDD.n1611 VDD.n1608 0.194439
R1746 VDD.n1622 VDD.n294 0.194439
R1747 VDD.n1622 VDD.n1607 0.194439
R1748 VDD.n1574 VDD.n295 0.194439
R1749 VDD.n1577 VDD.n1574 0.194439
R1750 VDD.n1588 VDD.n318 0.194439
R1751 VDD.n1588 VDD.n1573 0.194439
R1752 VDD.n348 VDD.n319 0.194439
R1753 VDD.n351 VDD.n348 0.194439
R1754 VDD.n1551 VDD.n355 0.194439
R1755 VDD.n1551 VDD.n1550 0.194439
R1756 VDD.n1539 VDD.n370 0.194439
R1757 VDD.n1539 VDD.n1538 0.194439
R1758 VDD.n1527 VDD.n386 0.194439
R1759 VDD.n1527 VDD.n1526 0.194439
R1760 VDD.n1515 VDD.n402 0.194439
R1761 VDD.n1515 VDD.n1514 0.194439
R1762 VDD.n1503 VDD.n417 0.194439
R1763 VDD.n1503 VDD.n1500 0.194439
R1764 VDD.n1489 VDD.n433 0.194439
R1765 VDD.n1489 VDD.n1488 0.194439
R1766 VDD.n1480 VDD.n1479 0.194439
R1767 VDD.n1479 VDD.n1478 0.194439
R1768 VDD.n1445 VDD.n439 0.194439
R1769 VDD.n1448 VDD.n1445 0.194439
R1770 VDD.n1459 VDD.n471 0.194439
R1771 VDD.n1459 VDD.n1444 0.194439
R1772 VDD.n1411 VDD.n472 0.194439
R1773 VDD.n1414 VDD.n1411 0.194439
R1774 VDD.n1425 VDD.n495 0.194439
R1775 VDD.n1425 VDD.n1410 0.194439
R1776 VDD.n525 VDD.n496 0.194439
R1777 VDD.n528 VDD.n525 0.194439
R1778 VDD.n1388 VDD.n532 0.194439
R1779 VDD.n1388 VDD.n1387 0.194439
R1780 VDD.n1376 VDD.n547 0.194439
R1781 VDD.n1376 VDD.n1375 0.194439
R1782 VDD.n1364 VDD.n563 0.194439
R1783 VDD.n1364 VDD.n1363 0.194439
R1784 VDD.n1352 VDD.n579 0.194439
R1785 VDD.n1352 VDD.n1351 0.194439
R1786 VDD.n1340 VDD.n594 0.194439
R1787 VDD.n1340 VDD.n1337 0.194439
R1788 VDD.n1326 VDD.n610 0.194439
R1789 VDD.n1326 VDD.n1325 0.194439
R1790 VDD.n1317 VDD.n1316 0.194439
R1791 VDD.n1316 VDD.n1315 0.194439
R1792 VDD.n1282 VDD.n616 0.194439
R1793 VDD.n1285 VDD.n1282 0.194439
R1794 VDD.n1296 VDD.n648 0.194439
R1795 VDD.n1296 VDD.n1281 0.194439
R1796 VDD.n1248 VDD.n649 0.194439
R1797 VDD.n1251 VDD.n1248 0.194439
R1798 VDD.n1262 VDD.n672 0.194439
R1799 VDD.n1262 VDD.n1247 0.194439
R1800 VDD.n702 VDD.n673 0.194439
R1801 VDD.n705 VDD.n702 0.194439
R1802 VDD.n1225 VDD.n709 0.194439
R1803 VDD.n1225 VDD.n1224 0.194439
R1804 VDD.n1213 VDD.n724 0.194439
R1805 VDD.n1213 VDD.n1212 0.194439
R1806 VDD.n1201 VDD.n740 0.194439
R1807 VDD.n1201 VDD.n1200 0.194439
R1808 VDD.n1189 VDD.n756 0.194439
R1809 VDD.n1189 VDD.n1188 0.194439
R1810 VDD.n1177 VDD.n771 0.194439
R1811 VDD.n1177 VDD.n1174 0.194439
R1812 VDD.n1163 VDD.n787 0.194439
R1813 VDD.n1163 VDD.n1162 0.194439
R1814 VDD.n1154 VDD.n1153 0.194439
R1815 VDD.n1153 VDD.n1152 0.194439
R1816 VDD.n1119 VDD.n793 0.194439
R1817 VDD.n1122 VDD.n1119 0.194439
R1818 VDD.n1133 VDD.n825 0.194439
R1819 VDD.n1133 VDD.n1118 0.194439
R1820 VDD.n1085 VDD.n826 0.194439
R1821 VDD.n1088 VDD.n1085 0.194439
R1822 VDD.n1099 VDD.n849 0.194439
R1823 VDD.n1099 VDD.n1084 0.194439
R1824 VDD.n852 VDD.n850 0.194439
R1825 VDD.n884 VDD.n881 0.194439
R1826 VDD.n1056 VDD.n878 0.194439
R1827 VDD.n1056 VDD.n879 0.194439
R1828 VDD.n921 VDD.n894 0.194439
R1829 VDD.n922 VDD.n921 0.194439
R1830 VDD.n1035 VDD.n917 0.194439
R1831 VDD.n1035 VDD.n918 0.194439
R1832 VDD.n1001 VDD.n933 0.194439
R1833 VDD.n1002 VDD.n1001 0.194439
R1834 VDD.n1014 VDD.n956 0.194439
R1835 VDD.n1014 VDD.n957 0.194439
R1836 VDD.n977 VDD.n976 0.132407
R1837 VDD.n976 VDD.n955 0.127283
R1838 VDD.n1695 VDD 0.103754
R1839 VDD.n274 VDD.n273 0.102103
R1840 VDD.n451 VDD.n450 0.102103
R1841 VDD.n628 VDD.n627 0.102103
R1842 VDD.n805 VDD.n804 0.102103
R1843 VDD.n1559 VDD.n1558 0.100721
R1844 VDD.n1396 VDD.n1395 0.100721
R1845 VDD.n1233 VDD.n1232 0.100721
R1846 VDD VDD.n1068 0.100533
R1847 VDD.n1722 VDD.n27 0.0981562
R1848 VDD.n275 VDD.n272 0.0890769
R1849 VDD.n452 VDD.n449 0.0890769
R1850 VDD.n629 VDD.n626 0.0890769
R1851 VDD.n806 VDD.n803 0.0890769
R1852 VDD.n1132 VDD.n112 0.0847059
R1853 VDD.n1098 VDD.n110 0.0847059
R1854 VDD.n1295 VDD.n123 0.0847059
R1855 VDD.n1261 VDD.n121 0.0847059
R1856 VDD.n1458 VDD.n134 0.0847059
R1857 VDD.n1424 VDD.n132 0.0847059
R1858 VDD.n1621 VDD.n145 0.0847059
R1859 VDD.n1587 VDD.n143 0.0847059
R1860 VDD.n196 VDD.n73 0.0847059
R1861 VDD.n1055 VDD.n1054 0.0847059
R1862 VDD.n919 VDD.n893 0.0847059
R1863 VDD.n1034 VDD.n1033 0.0847059
R1864 VDD.n999 VDD.n932 0.0847059
R1865 VDD.n963 VDD.n958 0.0796667
R1866 VDD.n888 VDD.n885 0.0705758
R1867 VDD.n895 VDD.n877 0.0705758
R1868 VDD.n927 VDD.n923 0.0705758
R1869 VDD.n934 VDD.n916 0.0705758
R1870 VDD.n1007 VDD.n1003 0.0705758
R1871 VDD.n182 VDD.n170 0.0705758
R1872 VDD.n201 VDD.n153 0.0705758
R1873 VDD.n1681 VDD.n1680 0.0705758
R1874 VDD.n1668 VDD.n221 0.0705758
R1875 VDD.n1660 VDD.n238 0.0705758
R1876 VDD.n280 VDD.n263 0.0705758
R1877 VDD.n1616 VDD.n1612 0.0705758
R1878 VDD.n296 VDD.n293 0.0705758
R1879 VDD.n1582 VDD.n1578 0.0705758
R1880 VDD.n320 VDD.n317 0.0705758
R1881 VDD.n1547 VDD.n358 0.0705758
R1882 VDD.n1535 VDD.n373 0.0705758
R1883 VDD.n1523 VDD.n389 0.0705758
R1884 VDD.n1511 VDD.n405 0.0705758
R1885 VDD.n1497 VDD.n419 0.0705758
R1886 VDD.n457 VDD.n440 0.0705758
R1887 VDD.n1453 VDD.n1449 0.0705758
R1888 VDD.n473 VDD.n470 0.0705758
R1889 VDD.n1419 VDD.n1415 0.0705758
R1890 VDD.n497 VDD.n494 0.0705758
R1891 VDD.n1384 VDD.n535 0.0705758
R1892 VDD.n1372 VDD.n550 0.0705758
R1893 VDD.n1360 VDD.n566 0.0705758
R1894 VDD.n1348 VDD.n582 0.0705758
R1895 VDD.n1334 VDD.n596 0.0705758
R1896 VDD.n634 VDD.n617 0.0705758
R1897 VDD.n1290 VDD.n1286 0.0705758
R1898 VDD.n650 VDD.n647 0.0705758
R1899 VDD.n1256 VDD.n1252 0.0705758
R1900 VDD.n674 VDD.n671 0.0705758
R1901 VDD.n1221 VDD.n712 0.0705758
R1902 VDD.n1209 VDD.n727 0.0705758
R1903 VDD.n1197 VDD.n743 0.0705758
R1904 VDD.n1185 VDD.n759 0.0705758
R1905 VDD.n1171 VDD.n773 0.0705758
R1906 VDD.n811 VDD.n794 0.0705758
R1907 VDD.n1127 VDD.n1123 0.0705758
R1908 VDD.n827 VDD.n824 0.0705758
R1909 VDD.n1093 VDD.n1089 0.0705758
R1910 VDD.n851 VDD.n848 0.0705758
R1911 VDD.n1560 VDD 0.0619615
R1912 VDD.n1397 VDD 0.0619615
R1913 VDD.n1234 VDD 0.0619615
R1914 VDD.n1071 VDD 0.0619615
R1915 VDD.n7 VDD.n0 0.0616979
R1916 VDD VDD.n7 0.0603958
R1917 VDD.n1744 VDD.n0 0.0590938
R1918 VDD.n961 VDD 0.0579444
R1919 VDD.n1723 VDD.n1722 0.0577917
R1920 VDD.n185 VDD.n183 0.0573182
R1921 VDD.n205 VDD.n202 0.0573182
R1922 VDD.n1682 VDD.n156 0.0573182
R1923 VDD.n1670 VDD.n219 0.0573182
R1924 VDD.n1659 VDD.n1658 0.0573182
R1925 VDD.n282 VDD.n265 0.0573182
R1926 VDD.n1615 VDD.n1614 0.0573182
R1927 VDD.n306 VDD.n298 0.0573182
R1928 VDD.n1581 VDD.n1580 0.0573182
R1929 VDD.n330 VDD.n322 0.0573182
R1930 VDD.n1546 VDD.n1545 0.0573182
R1931 VDD.n1534 VDD.n1533 0.0573182
R1932 VDD.n1522 VDD.n1521 0.0573182
R1933 VDD.n1510 VDD.n1509 0.0573182
R1934 VDD.n1496 VDD.n1495 0.0573182
R1935 VDD.n459 VDD.n442 0.0573182
R1936 VDD.n1452 VDD.n1451 0.0573182
R1937 VDD.n483 VDD.n475 0.0573182
R1938 VDD.n1418 VDD.n1417 0.0573182
R1939 VDD.n507 VDD.n499 0.0573182
R1940 VDD.n1383 VDD.n1382 0.0573182
R1941 VDD.n1371 VDD.n1370 0.0573182
R1942 VDD.n1359 VDD.n1358 0.0573182
R1943 VDD.n1347 VDD.n1346 0.0573182
R1944 VDD.n1333 VDD.n1332 0.0573182
R1945 VDD.n636 VDD.n619 0.0573182
R1946 VDD.n1289 VDD.n1288 0.0573182
R1947 VDD.n660 VDD.n652 0.0573182
R1948 VDD.n1255 VDD.n1254 0.0573182
R1949 VDD.n684 VDD.n676 0.0573182
R1950 VDD.n1220 VDD.n1219 0.0573182
R1951 VDD.n1208 VDD.n1207 0.0573182
R1952 VDD.n1196 VDD.n1195 0.0573182
R1953 VDD.n1184 VDD.n1183 0.0573182
R1954 VDD.n1170 VDD.n1169 0.0573182
R1955 VDD.n813 VDD.n796 0.0573182
R1956 VDD.n1126 VDD.n1125 0.0573182
R1957 VDD.n837 VDD.n829 0.0573182
R1958 VDD.n1092 VDD.n1091 0.0573182
R1959 VDD.n862 VDD.n854 0.0573182
R1960 VDD.n887 VDD.n886 0.0573182
R1961 VDD.n905 VDD.n897 0.0573182
R1962 VDD.n926 VDD.n925 0.0573182
R1963 VDD.n944 VDD.n936 0.0573182
R1964 VDD.n1006 VDD.n1005 0.0573182
R1965 VDD.n1728 VDD.n23 0.0517727
R1966 VDD.n975 VDD.n958 0.0455
R1967 VDD.n18 VDD.n15 0.0438377
R1968 VDD.n885 VDD.n869 0.0429036
R1969 VDD.n1727 VDD.n1726 0.041625
R1970 VDD.n1723 VDD 0.0408646
R1971 VDD.n1057 VDD.n877 0.0402727
R1972 VDD.n923 VDD.n896 0.0402727
R1973 VDD.n1036 VDD.n916 0.0402727
R1974 VDD.n1003 VDD.n935 0.0402727
R1975 VDD.n1015 VDD.n955 0.0402727
R1976 VDD.n194 VDD.n170 0.0402727
R1977 VDD.n1685 VDD.n153 0.0402727
R1978 VDD.n1680 VDD.n157 0.0402727
R1979 VDD.n1668 VDD.n1667 0.0402727
R1980 VDD.n1653 VDD.n238 0.0402727
R1981 VDD.n280 VDD.n261 0.0402727
R1982 VDD.n1612 VDD.n264 0.0402727
R1983 VDD.n1623 VDD.n293 0.0402727
R1984 VDD.n1578 VDD.n297 0.0402727
R1985 VDD.n1589 VDD.n317 0.0402727
R1986 VDD.n345 VDD.n321 0.0402727
R1987 VDD.n1552 VDD.n346 0.0402727
R1988 VDD.n1540 VDD.n358 0.0402727
R1989 VDD.n1528 VDD.n373 0.0402727
R1990 VDD.n1516 VDD.n389 0.0402727
R1991 VDD.n1504 VDD.n405 0.0402727
R1992 VDD.n1490 VDD.n419 0.0402727
R1993 VDD.n457 VDD.n438 0.0402727
R1994 VDD.n1449 VDD.n441 0.0402727
R1995 VDD.n1460 VDD.n470 0.0402727
R1996 VDD.n1415 VDD.n474 0.0402727
R1997 VDD.n1426 VDD.n494 0.0402727
R1998 VDD.n522 VDD.n498 0.0402727
R1999 VDD.n1389 VDD.n523 0.0402727
R2000 VDD.n1377 VDD.n535 0.0402727
R2001 VDD.n1365 VDD.n550 0.0402727
R2002 VDD.n1353 VDD.n566 0.0402727
R2003 VDD.n1341 VDD.n582 0.0402727
R2004 VDD.n1327 VDD.n596 0.0402727
R2005 VDD.n634 VDD.n615 0.0402727
R2006 VDD.n1286 VDD.n618 0.0402727
R2007 VDD.n1297 VDD.n647 0.0402727
R2008 VDD.n1252 VDD.n651 0.0402727
R2009 VDD.n1263 VDD.n671 0.0402727
R2010 VDD.n699 VDD.n675 0.0402727
R2011 VDD.n1226 VDD.n700 0.0402727
R2012 VDD.n1214 VDD.n712 0.0402727
R2013 VDD.n1202 VDD.n727 0.0402727
R2014 VDD.n1190 VDD.n743 0.0402727
R2015 VDD.n1178 VDD.n759 0.0402727
R2016 VDD.n1164 VDD.n773 0.0402727
R2017 VDD.n811 VDD.n792 0.0402727
R2018 VDD.n1123 VDD.n795 0.0402727
R2019 VDD.n1134 VDD.n824 0.0402727
R2020 VDD.n1089 VDD.n828 0.0402727
R2021 VDD.n1100 VDD.n848 0.0402727
R2022 VDD.n183 VDD.n178 0.0402727
R2023 VDD.n202 VDD.n165 0.0402727
R2024 VDD.n1683 VDD.n1682 0.0402727
R2025 VDD.n230 VDD.n219 0.0402727
R2026 VDD.n1659 VDD.n239 0.0402727
R2027 VDD.n1647 VDD.n251 0.0402727
R2028 VDD.n1646 VDD.n1645 0.0402727
R2029 VDD.n1634 VDD.n265 0.0402727
R2030 VDD.n1615 VDD.n290 0.0402727
R2031 VDD.n1600 VDD.n298 0.0402727
R2032 VDD.n1581 VDD.n314 0.0402727
R2033 VDD.n1566 VDD.n322 0.0402727
R2034 VDD.n1546 VDD.n340 0.0402727
R2035 VDD.n1534 VDD.n366 0.0402727
R2036 VDD.n1522 VDD.n382 0.0402727
R2037 VDD.n1510 VDD.n398 0.0402727
R2038 VDD.n1496 VDD.n414 0.0402727
R2039 VDD.n1484 VDD.n428 0.0402727
R2040 VDD.n1483 VDD.n1482 0.0402727
R2041 VDD.n1471 VDD.n442 0.0402727
R2042 VDD.n1452 VDD.n467 0.0402727
R2043 VDD.n1437 VDD.n475 0.0402727
R2044 VDD.n1418 VDD.n491 0.0402727
R2045 VDD.n1403 VDD.n499 0.0402727
R2046 VDD.n1383 VDD.n517 0.0402727
R2047 VDD.n1371 VDD.n543 0.0402727
R2048 VDD.n1359 VDD.n559 0.0402727
R2049 VDD.n1347 VDD.n575 0.0402727
R2050 VDD.n1333 VDD.n591 0.0402727
R2051 VDD.n1321 VDD.n605 0.0402727
R2052 VDD.n1320 VDD.n1319 0.0402727
R2053 VDD.n1308 VDD.n619 0.0402727
R2054 VDD.n1289 VDD.n644 0.0402727
R2055 VDD.n1274 VDD.n652 0.0402727
R2056 VDD.n1255 VDD.n668 0.0402727
R2057 VDD.n1240 VDD.n676 0.0402727
R2058 VDD.n1220 VDD.n694 0.0402727
R2059 VDD.n1208 VDD.n720 0.0402727
R2060 VDD.n1196 VDD.n736 0.0402727
R2061 VDD.n1184 VDD.n752 0.0402727
R2062 VDD.n1170 VDD.n768 0.0402727
R2063 VDD.n1158 VDD.n782 0.0402727
R2064 VDD.n1157 VDD.n1156 0.0402727
R2065 VDD.n1145 VDD.n796 0.0402727
R2066 VDD.n1126 VDD.n821 0.0402727
R2067 VDD.n1111 VDD.n829 0.0402727
R2068 VDD.n1092 VDD.n845 0.0402727
R2069 VDD.n1077 VDD.n854 0.0402727
R2070 VDD.n887 VDD.n874 0.0402727
R2071 VDD.n1047 VDD.n897 0.0402727
R2072 VDD.n926 VDD.n913 0.0402727
R2073 VDD.n1026 VDD.n936 0.0402727
R2074 VDD.n1006 VDD.n952 0.0402727
R2075 VDD.n1692 VDD.n68 0.0364848
R2076 VDD.n184 VDD.n171 0.0364848
R2077 VDD.n204 VDD.n203 0.0364848
R2078 VDD.n1679 VDD.n1678 0.0364848
R2079 VDD.n1669 VDD.n220 0.0364848
R2080 VDD.n1655 VDD.n240 0.0364848
R2081 VDD.n281 VDD.n279 0.0364848
R2082 VDD.n1613 VDD.n266 0.0364848
R2083 VDD.n305 VDD.n291 0.0364848
R2084 VDD.n1579 VDD.n299 0.0364848
R2085 VDD.n329 VDD.n315 0.0364848
R2086 VDD.n344 VDD.n323 0.0364848
R2087 VDD.n1554 VDD.n339 0.0364848
R2088 VDD.n1542 VDD.n359 0.0364848
R2089 VDD.n1530 VDD.n374 0.0364848
R2090 VDD.n1518 VDD.n390 0.0364848
R2091 VDD.n1506 VDD.n406 0.0364848
R2092 VDD.n1492 VDD.n420 0.0364848
R2093 VDD.n458 VDD.n456 0.0364848
R2094 VDD.n1450 VDD.n443 0.0364848
R2095 VDD.n482 VDD.n468 0.0364848
R2096 VDD.n1416 VDD.n476 0.0364848
R2097 VDD.n506 VDD.n492 0.0364848
R2098 VDD.n521 VDD.n500 0.0364848
R2099 VDD.n1391 VDD.n516 0.0364848
R2100 VDD.n1379 VDD.n536 0.0364848
R2101 VDD.n1367 VDD.n551 0.0364848
R2102 VDD.n1355 VDD.n567 0.0364848
R2103 VDD.n1343 VDD.n583 0.0364848
R2104 VDD.n1329 VDD.n597 0.0364848
R2105 VDD.n635 VDD.n633 0.0364848
R2106 VDD.n1287 VDD.n620 0.0364848
R2107 VDD.n659 VDD.n645 0.0364848
R2108 VDD.n1253 VDD.n653 0.0364848
R2109 VDD.n683 VDD.n669 0.0364848
R2110 VDD.n698 VDD.n677 0.0364848
R2111 VDD.n1228 VDD.n693 0.0364848
R2112 VDD.n1216 VDD.n713 0.0364848
R2113 VDD.n1204 VDD.n728 0.0364848
R2114 VDD.n1192 VDD.n744 0.0364848
R2115 VDD.n1180 VDD.n760 0.0364848
R2116 VDD.n1166 VDD.n774 0.0364848
R2117 VDD.n812 VDD.n810 0.0364848
R2118 VDD.n1124 VDD.n797 0.0364848
R2119 VDD.n836 VDD.n822 0.0364848
R2120 VDD.n1090 VDD.n830 0.0364848
R2121 VDD.n861 VDD.n846 0.0364848
R2122 VDD.n1069 VDD.n855 0.0364848
R2123 VDD.n1065 VDD.n870 0.0364848
R2124 VDD.n904 VDD.n875 0.0364848
R2125 VDD.n924 VDD.n898 0.0364848
R2126 VDD.n943 VDD.n914 0.0364848
R2127 VDD.n1004 VDD.n937 0.0364848
R2128 VDD.n962 VDD.n953 0.0364848
R2129 VDD.n17 VDD.n16 0.0351948
R2130 VDD.n1731 VDD.n10 0.0309054
R2131 VDD.n889 VDD.n876 0.030803
R2132 VDD.n1049 VDD.n1048 0.030803
R2133 VDD.n928 VDD.n915 0.030803
R2134 VDD.n1028 VDD.n1027 0.030803
R2135 VDD.n1008 VDD.n954 0.030803
R2136 VDD.n181 VDD.n70 0.030803
R2137 VDD.n200 VDD.n166 0.030803
R2138 VDD.n1684 VDD.n155 0.030803
R2139 VDD.n232 VDD.n231 0.030803
R2140 VDD.n1661 VDD.n223 0.030803
R2141 VDD.n1649 VDD.n253 0.030803
R2142 VDD.n1644 VDD.n260 0.030803
R2143 VDD.n1636 VDD.n1635 0.030803
R2144 VDD.n1617 VDD.n292 0.030803
R2145 VDD.n1602 VDD.n1601 0.030803
R2146 VDD.n1583 VDD.n316 0.030803
R2147 VDD.n1568 VDD.n1567 0.030803
R2148 VDD.n1548 VDD.n347 0.030803
R2149 VDD.n1536 VDD.n368 0.030803
R2150 VDD.n1524 VDD.n384 0.030803
R2151 VDD.n1512 VDD.n400 0.030803
R2152 VDD.n1498 VDD.n416 0.030803
R2153 VDD.n1486 VDD.n430 0.030803
R2154 VDD.n1481 VDD.n437 0.030803
R2155 VDD.n1473 VDD.n1472 0.030803
R2156 VDD.n1454 VDD.n469 0.030803
R2157 VDD.n1439 VDD.n1438 0.030803
R2158 VDD.n1420 VDD.n493 0.030803
R2159 VDD.n1405 VDD.n1404 0.030803
R2160 VDD.n1385 VDD.n524 0.030803
R2161 VDD.n1373 VDD.n545 0.030803
R2162 VDD.n1361 VDD.n561 0.030803
R2163 VDD.n1349 VDD.n577 0.030803
R2164 VDD.n1335 VDD.n593 0.030803
R2165 VDD.n1323 VDD.n607 0.030803
R2166 VDD.n1318 VDD.n614 0.030803
R2167 VDD.n1310 VDD.n1309 0.030803
R2168 VDD.n1291 VDD.n646 0.030803
R2169 VDD.n1276 VDD.n1275 0.030803
R2170 VDD.n1257 VDD.n670 0.030803
R2171 VDD.n1242 VDD.n1241 0.030803
R2172 VDD.n1222 VDD.n701 0.030803
R2173 VDD.n1210 VDD.n722 0.030803
R2174 VDD.n1198 VDD.n738 0.030803
R2175 VDD.n1186 VDD.n754 0.030803
R2176 VDD.n1172 VDD.n770 0.030803
R2177 VDD.n1160 VDD.n784 0.030803
R2178 VDD.n1155 VDD.n791 0.030803
R2179 VDD.n1147 VDD.n1146 0.030803
R2180 VDD.n1128 VDD.n823 0.030803
R2181 VDD.n1113 VDD.n1112 0.030803
R2182 VDD.n1094 VDD.n847 0.030803
R2183 VDD.n1079 VDD.n1078 0.030803
R2184 VDD.n26 VDD.n9 0.0292162
R2185 VDD.n49 VDD.n48 0.0273994
R2186 VDD.n8 VDD 0.0265417
R2187 VDD.n1710 VDD.n29 0.0242893
R2188 VDD.n988 VDD.n52 0.0242893
R2189 VDD.n985 VDD.n56 0.0242893
R2190 VDD.n982 VDD.n60 0.0242893
R2191 VDD.n978 VDD.n64 0.0242893
R2192 VDD.n1732 VDD.n8 0.0239375
R2193 VDD.n39 VDD.n38 0.0234759
R2194 VDD VDD.n1744 0.0226354
R2195 VDD.n970 VDD.n969 0.0206084
R2196 VDD.n177 VDD.n176 0.0205441
R2197 VDD.n192 VDD.n164 0.0205441
R2198 VDD.n213 VDD.n212 0.0205441
R2199 VDD.n1673 VDD.n217 0.0205441
R2200 VDD.n247 VDD.n246 0.0205441
R2201 VDD.n273 VDD.n252 0.0205441
R2202 VDD.n362 VDD.n341 0.0205441
R2203 VDD.n378 VDD.n367 0.0205441
R2204 VDD.n394 VDD.n383 0.0205441
R2205 VDD.n410 VDD.n399 0.0205441
R2206 VDD.n424 VDD.n415 0.0205441
R2207 VDD.n450 VDD.n429 0.0205441
R2208 VDD.n539 VDD.n518 0.0205441
R2209 VDD.n555 VDD.n544 0.0205441
R2210 VDD.n571 VDD.n560 0.0205441
R2211 VDD.n587 VDD.n576 0.0205441
R2212 VDD.n601 VDD.n592 0.0205441
R2213 VDD.n627 VDD.n606 0.0205441
R2214 VDD.n716 VDD.n695 0.0205441
R2215 VDD.n732 VDD.n721 0.0205441
R2216 VDD.n748 VDD.n737 0.0205441
R2217 VDD.n764 VDD.n753 0.0205441
R2218 VDD.n778 VDD.n769 0.0205441
R2219 VDD.n804 VDD.n783 0.0205441
R2220 VDD.n274 VDD.n270 0.0198529
R2221 VDD.n1632 VDD.n267 0.0198529
R2222 VDD.n1626 VDD.n1625 0.0198529
R2223 VDD.n1598 VDD.n300 0.0198529
R2224 VDD.n1592 VDD.n1591 0.0198529
R2225 VDD.n1564 VDD.n324 0.0198529
R2226 VDD.n451 VDD.n447 0.0198529
R2227 VDD.n1469 VDD.n444 0.0198529
R2228 VDD.n1463 VDD.n1462 0.0198529
R2229 VDD.n1435 VDD.n477 0.0198529
R2230 VDD.n1429 VDD.n1428 0.0198529
R2231 VDD.n1401 VDD.n501 0.0198529
R2232 VDD.n628 VDD.n624 0.0198529
R2233 VDD.n1306 VDD.n621 0.0198529
R2234 VDD.n1300 VDD.n1299 0.0198529
R2235 VDD.n1272 VDD.n654 0.0198529
R2236 VDD.n1266 VDD.n1265 0.0198529
R2237 VDD.n1238 VDD.n678 0.0198529
R2238 VDD.n805 VDD.n801 0.0198529
R2239 VDD.n1143 VDD.n798 0.0198529
R2240 VDD.n1137 VDD.n1136 0.0198529
R2241 VDD.n1109 VDD.n831 0.0198529
R2242 VDD.n1103 VDD.n1102 0.0198529
R2243 VDD.n1075 VDD.n856 0.0198529
R2244 VDD.n1060 VDD.n1059 0.0198529
R2245 VDD.n1045 VDD.n899 0.0198529
R2246 VDD.n1039 VDD.n1038 0.0198529
R2247 VDD.n1024 VDD.n938 0.0198529
R2248 VDD.n1018 VDD.n1017 0.0198529
R2249 VDD.n1728 VDD.n12 0.0188117
R2250 VDD.n15 VDD.n12 0.0188117
R2251 VDD.n174 VDD.n173 0.0185769
R2252 VDD.n190 VDD.n163 0.0185769
R2253 VDD.n210 VDD.n161 0.0185769
R2254 VDD.n1675 VDD.n1674 0.0185769
R2255 VDD.n248 VDD.n244 0.0185769
R2256 VDD.n272 VDD.n271 0.0185769
R2257 VDD.n285 VDD.n269 0.0185769
R2258 VDD.n1629 VDD.n1628 0.0185769
R2259 VDD.n309 VDD.n303 0.0185769
R2260 VDD.n1595 VDD.n1594 0.0185769
R2261 VDD.n333 VDD.n327 0.0185769
R2262 VDD.n1561 VDD.n1560 0.0185769
R2263 VDD.n363 VDD.n337 0.0185769
R2264 VDD.n379 VDD.n377 0.0185769
R2265 VDD.n395 VDD.n393 0.0185769
R2266 VDD.n411 VDD.n409 0.0185769
R2267 VDD.n425 VDD.n423 0.0185769
R2268 VDD.n449 VDD.n448 0.0185769
R2269 VDD.n462 VDD.n446 0.0185769
R2270 VDD.n1466 VDD.n1465 0.0185769
R2271 VDD.n486 VDD.n480 0.0185769
R2272 VDD.n1432 VDD.n1431 0.0185769
R2273 VDD.n510 VDD.n504 0.0185769
R2274 VDD.n1398 VDD.n1397 0.0185769
R2275 VDD.n540 VDD.n514 0.0185769
R2276 VDD.n556 VDD.n554 0.0185769
R2277 VDD.n572 VDD.n570 0.0185769
R2278 VDD.n588 VDD.n586 0.0185769
R2279 VDD.n602 VDD.n600 0.0185769
R2280 VDD.n626 VDD.n625 0.0185769
R2281 VDD.n639 VDD.n623 0.0185769
R2282 VDD.n1303 VDD.n1302 0.0185769
R2283 VDD.n663 VDD.n657 0.0185769
R2284 VDD.n1269 VDD.n1268 0.0185769
R2285 VDD.n687 VDD.n681 0.0185769
R2286 VDD.n1235 VDD.n1234 0.0185769
R2287 VDD.n717 VDD.n691 0.0185769
R2288 VDD.n733 VDD.n731 0.0185769
R2289 VDD.n749 VDD.n747 0.0185769
R2290 VDD.n765 VDD.n763 0.0185769
R2291 VDD.n779 VDD.n777 0.0185769
R2292 VDD.n803 VDD.n802 0.0185769
R2293 VDD.n816 VDD.n800 0.0185769
R2294 VDD.n1140 VDD.n1139 0.0185769
R2295 VDD.n840 VDD.n834 0.0185769
R2296 VDD.n1106 VDD.n1105 0.0185769
R2297 VDD.n865 VDD.n859 0.0185769
R2298 VDD.n1072 VDD.n1071 0.0185769
R2299 VDD.n971 VDD.n961 0.0185349
R2300 VDD.n1693 VDD.n67 0.0184706
R2301 VDD.n186 VDD.n172 0.0184706
R2302 VDD.n206 VDD.n162 0.0184706
R2303 VDD.n1677 VDD.n159 0.0184706
R2304 VDD.n1671 VDD.n218 0.0184706
R2305 VDD.n1657 VDD.n1656 0.0184706
R2306 VDD.n283 VDD.n278 0.0184706
R2307 VDD.n288 VDD.n268 0.0184706
R2308 VDD.n307 VDD.n304 0.0184706
R2309 VDD.n312 VDD.n301 0.0184706
R2310 VDD.n331 VDD.n328 0.0184706
R2311 VDD.n335 VDD.n325 0.0184706
R2312 VDD.n1555 VDD.n336 0.0184706
R2313 VDD.n1544 VDD.n1543 0.0184706
R2314 VDD.n1532 VDD.n1531 0.0184706
R2315 VDD.n1520 VDD.n1519 0.0184706
R2316 VDD.n1508 VDD.n1507 0.0184706
R2317 VDD.n1494 VDD.n1493 0.0184706
R2318 VDD.n460 VDD.n455 0.0184706
R2319 VDD.n465 VDD.n445 0.0184706
R2320 VDD.n484 VDD.n481 0.0184706
R2321 VDD.n489 VDD.n478 0.0184706
R2322 VDD.n508 VDD.n505 0.0184706
R2323 VDD.n512 VDD.n502 0.0184706
R2324 VDD.n1392 VDD.n513 0.0184706
R2325 VDD.n1381 VDD.n1380 0.0184706
R2326 VDD.n1369 VDD.n1368 0.0184706
R2327 VDD.n1357 VDD.n1356 0.0184706
R2328 VDD.n1345 VDD.n1344 0.0184706
R2329 VDD.n1331 VDD.n1330 0.0184706
R2330 VDD.n637 VDD.n632 0.0184706
R2331 VDD.n642 VDD.n622 0.0184706
R2332 VDD.n661 VDD.n658 0.0184706
R2333 VDD.n666 VDD.n655 0.0184706
R2334 VDD.n685 VDD.n682 0.0184706
R2335 VDD.n689 VDD.n679 0.0184706
R2336 VDD.n1229 VDD.n690 0.0184706
R2337 VDD.n1218 VDD.n1217 0.0184706
R2338 VDD.n1206 VDD.n1205 0.0184706
R2339 VDD.n1194 VDD.n1193 0.0184706
R2340 VDD.n1182 VDD.n1181 0.0184706
R2341 VDD.n1168 VDD.n1167 0.0184706
R2342 VDD.n814 VDD.n809 0.0184706
R2343 VDD.n819 VDD.n799 0.0184706
R2344 VDD.n838 VDD.n835 0.0184706
R2345 VDD.n843 VDD.n832 0.0184706
R2346 VDD.n863 VDD.n860 0.0184706
R2347 VDD.n1070 VDD.n857 0.0184706
R2348 VDD.n1064 VDD.n871 0.0184706
R2349 VDD.n906 VDD.n903 0.0184706
R2350 VDD.n911 VDD.n900 0.0184706
R2351 VDD.n945 VDD.n942 0.0184706
R2352 VDD.n950 VDD.n939 0.0184706
R2353 VDD.n966 VDD.n964 0.0184706
R2354 VDD.n1694 VDD.n66 0.0179744
R2355 VDD.n189 VDD.n188 0.0179744
R2356 VDD.n209 VDD.n208 0.0179744
R2357 VDD.n1676 VDD.n215 0.0179744
R2358 VDD.n243 VDD.n216 0.0179744
R2359 VDD.n250 VDD.n249 0.0179744
R2360 VDD.n276 VDD.n275 0.0179744
R2361 VDD.n1630 VDD.n286 0.0179744
R2362 VDD.n302 VDD.n287 0.0179744
R2363 VDD.n1596 VDD.n310 0.0179744
R2364 VDD.n326 VDD.n311 0.0179744
R2365 VDD.n1562 VDD.n334 0.0179744
R2366 VDD.n1557 VDD.n1556 0.0179744
R2367 VDD.n365 VDD.n364 0.0179744
R2368 VDD.n381 VDD.n380 0.0179744
R2369 VDD.n397 VDD.n396 0.0179744
R2370 VDD.n413 VDD.n412 0.0179744
R2371 VDD.n427 VDD.n426 0.0179744
R2372 VDD.n453 VDD.n452 0.0179744
R2373 VDD.n1467 VDD.n463 0.0179744
R2374 VDD.n479 VDD.n464 0.0179744
R2375 VDD.n1433 VDD.n487 0.0179744
R2376 VDD.n503 VDD.n488 0.0179744
R2377 VDD.n1399 VDD.n511 0.0179744
R2378 VDD.n1394 VDD.n1393 0.0179744
R2379 VDD.n542 VDD.n541 0.0179744
R2380 VDD.n558 VDD.n557 0.0179744
R2381 VDD.n574 VDD.n573 0.0179744
R2382 VDD.n590 VDD.n589 0.0179744
R2383 VDD.n604 VDD.n603 0.0179744
R2384 VDD.n630 VDD.n629 0.0179744
R2385 VDD.n1304 VDD.n640 0.0179744
R2386 VDD.n656 VDD.n641 0.0179744
R2387 VDD.n1270 VDD.n664 0.0179744
R2388 VDD.n680 VDD.n665 0.0179744
R2389 VDD.n1236 VDD.n688 0.0179744
R2390 VDD.n1231 VDD.n1230 0.0179744
R2391 VDD.n719 VDD.n718 0.0179744
R2392 VDD.n735 VDD.n734 0.0179744
R2393 VDD.n751 VDD.n750 0.0179744
R2394 VDD.n767 VDD.n766 0.0179744
R2395 VDD.n781 VDD.n780 0.0179744
R2396 VDD.n807 VDD.n806 0.0179744
R2397 VDD.n1141 VDD.n817 0.0179744
R2398 VDD.n833 VDD.n818 0.0179744
R2399 VDD.n1107 VDD.n841 0.0179744
R2400 VDD.n858 VDD.n842 0.0179744
R2401 VDD.n1073 VDD.n866 0.0179744
R2402 VDD.n1063 VDD.n1062 0.0179074
R2403 VDD.n908 VDD.n902 0.0179074
R2404 VDD.n1042 VDD.n1041 0.0179074
R2405 VDD.n947 VDD.n941 0.0179074
R2406 VDD.n1021 VDD.n1020 0.0179074
R2407 VDD.n968 VDD.n967 0.0179074
R2408 VDD.n1068 VDD.n867 0.0173272
R2409 VDD.n901 VDD.n872 0.0173272
R2410 VDD.n1043 VDD.n909 0.0173272
R2411 VDD.n940 VDD.n910 0.0173272
R2412 VDD.n1022 VDD.n948 0.0173272
R2413 VDD.n965 VDD.n949 0.0173272
R2414 VDD.n42 VDD.n33 0.0172857
R2415 VDD.n972 VDD.n971 0.0168953
R2416 VDD.n972 VDD.n959 0.0168953
R2417 VDD.n1704 VDD.n1703 0.0167579
R2418 VDD.n1719 VDD.n6 0.016125
R2419 VDD.n47 VDD.n46 0.0156071
R2420 VDD.n1709 VDD.n30 0.0156071
R2421 VDD.n1705 VDD.n53 0.0156071
R2422 VDD.n1702 VDD.n57 0.0156071
R2423 VDD.n1699 VDD.n61 0.0156071
R2424 VDD.n1696 VDD.n65 0.0156071
R2425 VDD.n973 VDD.n960 0.0152558
R2426 VDD.n40 VDD.n37 0.0148621
R2427 VDD.n1708 VDD.n1706 0.0148365
R2428 VDD.n187 VDD.n177 0.0143235
R2429 VDD.n207 VDD.n164 0.0143235
R2430 VDD.n214 VDD.n213 0.0143235
R2431 VDD.n1673 VDD.n1672 0.0143235
R2432 VDD.n247 VDD.n241 0.0143235
R2433 VDD.n284 VDD.n267 0.0143235
R2434 VDD.n1627 VDD.n1626 0.0143235
R2435 VDD.n308 VDD.n300 0.0143235
R2436 VDD.n1593 VDD.n1592 0.0143235
R2437 VDD.n332 VDD.n324 0.0143235
R2438 VDD.n362 VDD.n360 0.0143235
R2439 VDD.n378 VDD.n375 0.0143235
R2440 VDD.n394 VDD.n391 0.0143235
R2441 VDD.n410 VDD.n407 0.0143235
R2442 VDD.n424 VDD.n421 0.0143235
R2443 VDD.n461 VDD.n444 0.0143235
R2444 VDD.n1464 VDD.n1463 0.0143235
R2445 VDD.n485 VDD.n477 0.0143235
R2446 VDD.n1430 VDD.n1429 0.0143235
R2447 VDD.n509 VDD.n501 0.0143235
R2448 VDD.n539 VDD.n537 0.0143235
R2449 VDD.n555 VDD.n552 0.0143235
R2450 VDD.n571 VDD.n568 0.0143235
R2451 VDD.n587 VDD.n584 0.0143235
R2452 VDD.n601 VDD.n598 0.0143235
R2453 VDD.n638 VDD.n621 0.0143235
R2454 VDD.n1301 VDD.n1300 0.0143235
R2455 VDD.n662 VDD.n654 0.0143235
R2456 VDD.n1267 VDD.n1266 0.0143235
R2457 VDD.n686 VDD.n678 0.0143235
R2458 VDD.n716 VDD.n714 0.0143235
R2459 VDD.n732 VDD.n729 0.0143235
R2460 VDD.n748 VDD.n745 0.0143235
R2461 VDD.n764 VDD.n761 0.0143235
R2462 VDD.n778 VDD.n775 0.0143235
R2463 VDD.n815 VDD.n798 0.0143235
R2464 VDD.n1138 VDD.n1137 0.0143235
R2465 VDD.n839 VDD.n831 0.0143235
R2466 VDD.n1104 VDD.n1103 0.0143235
R2467 VDD.n864 VDD.n856 0.0143235
R2468 VDD.n1061 VDD.n1060 0.0143235
R2469 VDD.n907 VDD.n899 0.0143235
R2470 VDD.n1040 VDD.n1039 0.0143235
R2471 VDD.n946 VDD.n938 0.0143235
R2472 VDD.n1019 VDD.n1018 0.0143235
R2473 VDD.n1701 VDD.n1700 0.0140975
R2474 VDD.n1731 VDD.n9 0.0140135
R2475 VDD.n185 VDD.n184 0.0137576
R2476 VDD.n205 VDD.n204 0.0137576
R2477 VDD.n1679 VDD.n156 0.0137576
R2478 VDD.n1670 VDD.n1669 0.0137576
R2479 VDD.n1658 VDD.n240 0.0137576
R2480 VDD.n282 VDD.n281 0.0137576
R2481 VDD.n1614 VDD.n1613 0.0137576
R2482 VDD.n306 VDD.n305 0.0137576
R2483 VDD.n1580 VDD.n1579 0.0137576
R2484 VDD.n330 VDD.n329 0.0137576
R2485 VDD.n344 VDD.n343 0.0137576
R2486 VDD.n342 VDD.n339 0.0137576
R2487 VDD.n1545 VDD.n359 0.0137576
R2488 VDD.n1533 VDD.n374 0.0137576
R2489 VDD.n1521 VDD.n390 0.0137576
R2490 VDD.n1509 VDD.n406 0.0137576
R2491 VDD.n1495 VDD.n420 0.0137576
R2492 VDD.n459 VDD.n458 0.0137576
R2493 VDD.n1451 VDD.n1450 0.0137576
R2494 VDD.n483 VDD.n482 0.0137576
R2495 VDD.n1417 VDD.n1416 0.0137576
R2496 VDD.n507 VDD.n506 0.0137576
R2497 VDD.n521 VDD.n520 0.0137576
R2498 VDD.n519 VDD.n516 0.0137576
R2499 VDD.n1382 VDD.n536 0.0137576
R2500 VDD.n1370 VDD.n551 0.0137576
R2501 VDD.n1358 VDD.n567 0.0137576
R2502 VDD.n1346 VDD.n583 0.0137576
R2503 VDD.n1332 VDD.n597 0.0137576
R2504 VDD.n636 VDD.n635 0.0137576
R2505 VDD.n1288 VDD.n1287 0.0137576
R2506 VDD.n660 VDD.n659 0.0137576
R2507 VDD.n1254 VDD.n1253 0.0137576
R2508 VDD.n684 VDD.n683 0.0137576
R2509 VDD.n698 VDD.n697 0.0137576
R2510 VDD.n696 VDD.n693 0.0137576
R2511 VDD.n1219 VDD.n713 0.0137576
R2512 VDD.n1207 VDD.n728 0.0137576
R2513 VDD.n1195 VDD.n744 0.0137576
R2514 VDD.n1183 VDD.n760 0.0137576
R2515 VDD.n1169 VDD.n774 0.0137576
R2516 VDD.n813 VDD.n812 0.0137576
R2517 VDD.n1125 VDD.n1124 0.0137576
R2518 VDD.n837 VDD.n836 0.0137576
R2519 VDD.n1091 VDD.n1090 0.0137576
R2520 VDD.n862 VDD.n861 0.0137576
R2521 VDD.n886 VDD.n870 0.0137576
R2522 VDD.n905 VDD.n904 0.0137576
R2523 VDD.n925 VDD.n924 0.0137576
R2524 VDD.n944 VDD.n943 0.0137576
R2525 VDD.n1005 VDD.n1004 0.0137576
R2526 VDD.n963 VDD.n962 0.0137576
R2527 VDD.n39 VDD.n35 0.0137243
R2528 VDD.n1730 VDD.n11 0.0137188
R2529 VDD.n1730 VDD.n13 0.0137188
R2530 VDD.n1726 VDD.n1725 0.0130393
R2531 VDD.n17 VDD.n14 0.0130393
R2532 VDD.n1698 VDD.n1697 0.0129151
R2533 VDD.n188 VDD.n173 0.0125513
R2534 VDD.n208 VDD.n163 0.0125513
R2535 VDD.n215 VDD.n161 0.0125513
R2536 VDD.n1674 VDD.n216 0.0125513
R2537 VDD.n249 VDD.n248 0.0125513
R2538 VDD.n286 VDD.n285 0.0125513
R2539 VDD.n1628 VDD.n287 0.0125513
R2540 VDD.n310 VDD.n309 0.0125513
R2541 VDD.n1594 VDD.n311 0.0125513
R2542 VDD.n334 VDD.n333 0.0125513
R2543 VDD.n364 VDD.n363 0.0125513
R2544 VDD.n380 VDD.n379 0.0125513
R2545 VDD.n396 VDD.n395 0.0125513
R2546 VDD.n412 VDD.n411 0.0125513
R2547 VDD.n426 VDD.n425 0.0125513
R2548 VDD.n463 VDD.n462 0.0125513
R2549 VDD.n1465 VDD.n464 0.0125513
R2550 VDD.n487 VDD.n486 0.0125513
R2551 VDD.n1431 VDD.n488 0.0125513
R2552 VDD.n511 VDD.n510 0.0125513
R2553 VDD.n541 VDD.n540 0.0125513
R2554 VDD.n557 VDD.n556 0.0125513
R2555 VDD.n573 VDD.n572 0.0125513
R2556 VDD.n589 VDD.n588 0.0125513
R2557 VDD.n603 VDD.n602 0.0125513
R2558 VDD.n640 VDD.n639 0.0125513
R2559 VDD.n1302 VDD.n641 0.0125513
R2560 VDD.n664 VDD.n663 0.0125513
R2561 VDD.n1268 VDD.n665 0.0125513
R2562 VDD.n688 VDD.n687 0.0125513
R2563 VDD.n718 VDD.n717 0.0125513
R2564 VDD.n734 VDD.n733 0.0125513
R2565 VDD.n750 VDD.n749 0.0125513
R2566 VDD.n766 VDD.n765 0.0125513
R2567 VDD.n780 VDD.n779 0.0125513
R2568 VDD.n817 VDD.n816 0.0125513
R2569 VDD.n1139 VDD.n818 0.0125513
R2570 VDD.n841 VDD.n840 0.0125513
R2571 VDD.n1105 VDD.n842 0.0125513
R2572 VDD.n866 VDD.n865 0.0125513
R2573 VDD.n1062 VDD.n872 0.0121049
R2574 VDD.n909 VDD.n908 0.0121049
R2575 VDD.n1041 VDD.n910 0.0121049
R2576 VDD.n948 VDD.n947 0.0121049
R2577 VDD.n1020 VDD.n949 0.0121049
R2578 VDD.n41 VDD.n36 0.0105714
R2579 VDD.n1711 VDD.n1710 0.0103794
R2580 VDD.n989 VDD.n52 0.0103794
R2581 VDD.n986 VDD.n56 0.0103794
R2582 VDD.n983 VDD.n60 0.0103794
R2583 VDD.n979 VDD.n64 0.0103794
R2584 VDD.n889 VDD.n888 0.0099697
R2585 VDD.n1049 VDD.n895 0.0099697
R2586 VDD.n928 VDD.n927 0.0099697
R2587 VDD.n1028 VDD.n934 0.0099697
R2588 VDD.n1008 VDD.n1007 0.0099697
R2589 VDD.n182 VDD.n181 0.0099697
R2590 VDD.n201 VDD.n200 0.0099697
R2591 VDD.n1681 VDD.n155 0.0099697
R2592 VDD.n232 VDD.n221 0.0099697
R2593 VDD.n1661 VDD.n1660 0.0099697
R2594 VDD.n1649 VDD.n1648 0.0099697
R2595 VDD.n260 VDD.n258 0.0099697
R2596 VDD.n1636 VDD.n263 0.0099697
R2597 VDD.n1617 VDD.n1616 0.0099697
R2598 VDD.n1602 VDD.n296 0.0099697
R2599 VDD.n1583 VDD.n1582 0.0099697
R2600 VDD.n1568 VDD.n320 0.0099697
R2601 VDD.n1548 VDD.n1547 0.0099697
R2602 VDD.n1536 VDD.n1535 0.0099697
R2603 VDD.n1524 VDD.n1523 0.0099697
R2604 VDD.n1512 VDD.n1511 0.0099697
R2605 VDD.n1498 VDD.n1497 0.0099697
R2606 VDD.n1486 VDD.n1485 0.0099697
R2607 VDD.n437 VDD.n435 0.0099697
R2608 VDD.n1473 VDD.n440 0.0099697
R2609 VDD.n1454 VDD.n1453 0.0099697
R2610 VDD.n1439 VDD.n473 0.0099697
R2611 VDD.n1420 VDD.n1419 0.0099697
R2612 VDD.n1405 VDD.n497 0.0099697
R2613 VDD.n1385 VDD.n1384 0.0099697
R2614 VDD.n1373 VDD.n1372 0.0099697
R2615 VDD.n1361 VDD.n1360 0.0099697
R2616 VDD.n1349 VDD.n1348 0.0099697
R2617 VDD.n1335 VDD.n1334 0.0099697
R2618 VDD.n1323 VDD.n1322 0.0099697
R2619 VDD.n614 VDD.n612 0.0099697
R2620 VDD.n1310 VDD.n617 0.0099697
R2621 VDD.n1291 VDD.n1290 0.0099697
R2622 VDD.n1276 VDD.n650 0.0099697
R2623 VDD.n1257 VDD.n1256 0.0099697
R2624 VDD.n1242 VDD.n674 0.0099697
R2625 VDD.n1222 VDD.n1221 0.0099697
R2626 VDD.n1210 VDD.n1209 0.0099697
R2627 VDD.n1198 VDD.n1197 0.0099697
R2628 VDD.n1186 VDD.n1185 0.0099697
R2629 VDD.n1172 VDD.n1171 0.0099697
R2630 VDD.n1160 VDD.n1159 0.0099697
R2631 VDD.n791 VDD.n789 0.0099697
R2632 VDD.n1147 VDD.n794 0.0099697
R2633 VDD.n1128 VDD.n1127 0.0099697
R2634 VDD.n1113 VDD.n827 0.0099697
R2635 VDD.n1094 VDD.n1093 0.0099697
R2636 VDD.n1079 VDD.n851 0.0099697
R2637 VDD.n1719 VDD.n27 0.00701042
R2638 VDD.n1733 VDD.n6 0.00701042
R2639 VDD.n1709 VDD.n31 0.00635126
R2640 VDD.n1705 VDD.n51 0.00635126
R2641 VDD.n1702 VDD.n55 0.00635126
R2642 VDD.n1699 VDD.n59 0.00635126
R2643 VDD.n1696 VDD.n63 0.00635126
R2644 VDD.n1695 VDD.n62 0.00493396
R2645 VDD.n1697 VDD.n62 0.00493396
R2646 VDD.n1698 VDD.n58 0.00493396
R2647 VDD.n1700 VDD.n58 0.00493396
R2648 VDD.n1701 VDD.n54 0.00493396
R2649 VDD.n1703 VDD.n54 0.00493396
R2650 VDD.n1704 VDD.n50 0.00493396
R2651 VDD.n1706 VDD.n50 0.00493396
R2652 VDD.n1708 VDD.n1707 0.00493396
R2653 VDD.n1707 VDD.n49 0.00493396
R2654 VDD.n48 VDD.n32 0.00493396
R2655 VDD.n43 VDD.n32 0.00493396
R2656 VDD.n25 VDD.n24 0.00490305
R2657 VDD.n1733 VDD.n1732 0.00440625
R2658 VDD.n1714 VDD.t17 0.00429204
R2659 VDD.n69 VDD.n68 0.00428788
R2660 VDD.n193 VDD.n171 0.00428788
R2661 VDD.n203 VDD.n154 0.00428788
R2662 VDD.n1678 VDD.n158 0.00428788
R2663 VDD.n222 VDD.n220 0.00428788
R2664 VDD.n1655 VDD.n1654 0.00428788
R2665 VDD.n279 VDD.n259 0.00428788
R2666 VDD.n1633 VDD.n266 0.00428788
R2667 VDD.n1624 VDD.n291 0.00428788
R2668 VDD.n1599 VDD.n299 0.00428788
R2669 VDD.n1590 VDD.n315 0.00428788
R2670 VDD.n1565 VDD.n323 0.00428788
R2671 VDD.n1554 VDD.n1553 0.00428788
R2672 VDD.n1542 VDD.n1541 0.00428788
R2673 VDD.n1530 VDD.n1529 0.00428788
R2674 VDD.n1518 VDD.n1517 0.00428788
R2675 VDD.n1506 VDD.n1505 0.00428788
R2676 VDD.n1492 VDD.n1491 0.00428788
R2677 VDD.n456 VDD.n436 0.00428788
R2678 VDD.n1470 VDD.n443 0.00428788
R2679 VDD.n1461 VDD.n468 0.00428788
R2680 VDD.n1436 VDD.n476 0.00428788
R2681 VDD.n1427 VDD.n492 0.00428788
R2682 VDD.n1402 VDD.n500 0.00428788
R2683 VDD.n1391 VDD.n1390 0.00428788
R2684 VDD.n1379 VDD.n1378 0.00428788
R2685 VDD.n1367 VDD.n1366 0.00428788
R2686 VDD.n1355 VDD.n1354 0.00428788
R2687 VDD.n1343 VDD.n1342 0.00428788
R2688 VDD.n1329 VDD.n1328 0.00428788
R2689 VDD.n633 VDD.n613 0.00428788
R2690 VDD.n1307 VDD.n620 0.00428788
R2691 VDD.n1298 VDD.n645 0.00428788
R2692 VDD.n1273 VDD.n653 0.00428788
R2693 VDD.n1264 VDD.n669 0.00428788
R2694 VDD.n1239 VDD.n677 0.00428788
R2695 VDD.n1228 VDD.n1227 0.00428788
R2696 VDD.n1216 VDD.n1215 0.00428788
R2697 VDD.n1204 VDD.n1203 0.00428788
R2698 VDD.n1192 VDD.n1191 0.00428788
R2699 VDD.n1180 VDD.n1179 0.00428788
R2700 VDD.n1166 VDD.n1165 0.00428788
R2701 VDD.n810 VDD.n790 0.00428788
R2702 VDD.n1144 VDD.n797 0.00428788
R2703 VDD.n1135 VDD.n822 0.00428788
R2704 VDD.n1110 VDD.n830 0.00428788
R2705 VDD.n1101 VDD.n846 0.00428788
R2706 VDD.n1076 VDD.n855 0.00428788
R2707 VDD.n1066 VDD.n1065 0.00428788
R2708 VDD.n1058 VDD.n875 0.00428788
R2709 VDD.n1046 VDD.n898 0.00428788
R2710 VDD.n1037 VDD.n914 0.00428788
R2711 VDD.n1025 VDD.n937 0.00428788
R2712 VDD.n1016 VDD.n953 0.00428788
R2713 VDD.n21 VDD.n20 0.00428087
R2714 VDD.n974 VDD.n973 0.00391036
R2715 VDD.n959 VDD 0.00377907
R2716 VDD.n1725 VDD.n24 0.00360776
R2717 VDD.n21 VDD.n14 0.00360776
R2718 VDD.n41 VDD.n34 0.00351641
R2719 VDD.n284 VDD.n283 0.00326471
R2720 VDD.n1627 VDD.n288 0.00326471
R2721 VDD.n308 VDD.n307 0.00326471
R2722 VDD.n1593 VDD.n312 0.00326471
R2723 VDD.n332 VDD.n331 0.00326471
R2724 VDD.n1559 VDD.n335 0.00326471
R2725 VDD.n461 VDD.n460 0.00326471
R2726 VDD.n1464 VDD.n465 0.00326471
R2727 VDD.n485 VDD.n484 0.00326471
R2728 VDD.n1430 VDD.n489 0.00326471
R2729 VDD.n509 VDD.n508 0.00326471
R2730 VDD.n1396 VDD.n512 0.00326471
R2731 VDD.n638 VDD.n637 0.00326471
R2732 VDD.n1301 VDD.n642 0.00326471
R2733 VDD.n662 VDD.n661 0.00326471
R2734 VDD.n1267 VDD.n666 0.00326471
R2735 VDD.n686 VDD.n685 0.00326471
R2736 VDD.n1233 VDD.n689 0.00326471
R2737 VDD.n815 VDD.n814 0.00326471
R2738 VDD.n1138 VDD.n819 0.00326471
R2739 VDD.n839 VDD.n838 0.00326471
R2740 VDD.n1104 VDD.n843 0.00326471
R2741 VDD.n864 VDD.n863 0.00326471
R2742 VDD.n1061 VDD.n871 0.00326471
R2743 VDD.n907 VDD.n906 0.00326471
R2744 VDD.n1040 VDD.n911 0.00326471
R2745 VDD.n946 VDD.n945 0.00326471
R2746 VDD.n1019 VDD.n950 0.00326471
R2747 VDD.n969 VDD.n964 0.00326471
R2748 VDD.n187 VDD.n186 0.00257353
R2749 VDD.n207 VDD.n206 0.00257353
R2750 VDD.n214 VDD.n159 0.00257353
R2751 VDD.n1672 VDD.n1671 0.00257353
R2752 VDD.n1657 VDD.n241 0.00257353
R2753 VDD.n1558 VDD.n336 0.00257353
R2754 VDD.n1544 VDD.n360 0.00257353
R2755 VDD.n1532 VDD.n375 0.00257353
R2756 VDD.n1520 VDD.n391 0.00257353
R2757 VDD.n1508 VDD.n407 0.00257353
R2758 VDD.n1494 VDD.n421 0.00257353
R2759 VDD.n1395 VDD.n513 0.00257353
R2760 VDD.n1381 VDD.n537 0.00257353
R2761 VDD.n1369 VDD.n552 0.00257353
R2762 VDD.n1357 VDD.n568 0.00257353
R2763 VDD.n1345 VDD.n584 0.00257353
R2764 VDD.n1331 VDD.n598 0.00257353
R2765 VDD.n1232 VDD.n690 0.00257353
R2766 VDD.n1218 VDD.n714 0.00257353
R2767 VDD.n1206 VDD.n729 0.00257353
R2768 VDD.n1194 VDD.n745 0.00257353
R2769 VDD.n1182 VDD.n761 0.00257353
R2770 VDD.n1168 VDD.n775 0.00257353
R2771 VDD.n1057 VDD.n876 0.00239394
R2772 VDD.n1048 VDD.n896 0.00239394
R2773 VDD.n1036 VDD.n915 0.00239394
R2774 VDD.n1027 VDD.n935 0.00239394
R2775 VDD.n1015 VDD.n954 0.00239394
R2776 VDD.n1691 VDD.n70 0.00239394
R2777 VDD.n194 VDD.n166 0.00239394
R2778 VDD.n1685 VDD.n1684 0.00239394
R2779 VDD.n231 VDD.n157 0.00239394
R2780 VDD.n1667 VDD.n223 0.00239394
R2781 VDD.n1653 VDD.n253 0.00239394
R2782 VDD.n1644 VDD.n261 0.00239394
R2783 VDD.n1635 VDD.n264 0.00239394
R2784 VDD.n1623 VDD.n292 0.00239394
R2785 VDD.n1601 VDD.n297 0.00239394
R2786 VDD.n1589 VDD.n316 0.00239394
R2787 VDD.n1567 VDD.n321 0.00239394
R2788 VDD.n1552 VDD.n347 0.00239394
R2789 VDD.n1540 VDD.n368 0.00239394
R2790 VDD.n1528 VDD.n384 0.00239394
R2791 VDD.n1516 VDD.n400 0.00239394
R2792 VDD.n1504 VDD.n416 0.00239394
R2793 VDD.n1490 VDD.n430 0.00239394
R2794 VDD.n1481 VDD.n438 0.00239394
R2795 VDD.n1472 VDD.n441 0.00239394
R2796 VDD.n1460 VDD.n469 0.00239394
R2797 VDD.n1438 VDD.n474 0.00239394
R2798 VDD.n1426 VDD.n493 0.00239394
R2799 VDD.n1404 VDD.n498 0.00239394
R2800 VDD.n1389 VDD.n524 0.00239394
R2801 VDD.n1377 VDD.n545 0.00239394
R2802 VDD.n1365 VDD.n561 0.00239394
R2803 VDD.n1353 VDD.n577 0.00239394
R2804 VDD.n1341 VDD.n593 0.00239394
R2805 VDD.n1327 VDD.n607 0.00239394
R2806 VDD.n1318 VDD.n615 0.00239394
R2807 VDD.n1309 VDD.n618 0.00239394
R2808 VDD.n1297 VDD.n646 0.00239394
R2809 VDD.n1275 VDD.n651 0.00239394
R2810 VDD.n1263 VDD.n670 0.00239394
R2811 VDD.n1241 VDD.n675 0.00239394
R2812 VDD.n1226 VDD.n701 0.00239394
R2813 VDD.n1214 VDD.n722 0.00239394
R2814 VDD.n1202 VDD.n738 0.00239394
R2815 VDD.n1190 VDD.n754 0.00239394
R2816 VDD.n1178 VDD.n770 0.00239394
R2817 VDD.n1164 VDD.n784 0.00239394
R2818 VDD.n1155 VDD.n792 0.00239394
R2819 VDD.n1146 VDD.n795 0.00239394
R2820 VDD.n1134 VDD.n823 0.00239394
R2821 VDD.n1112 VDD.n828 0.00239394
R2822 VDD.n1100 VDD.n847 0.00239394
R2823 VDD.n1078 VDD.n853 0.00239394
R2824 VDD.n178 VDD.n69 0.00239394
R2825 VDD.n193 VDD.n165 0.00239394
R2826 VDD.n1683 VDD.n154 0.00239394
R2827 VDD.n230 VDD.n158 0.00239394
R2828 VDD.n239 VDD.n222 0.00239394
R2829 VDD.n1654 VDD.n251 0.00239394
R2830 VDD.n1645 VDD.n259 0.00239394
R2831 VDD.n1634 VDD.n1633 0.00239394
R2832 VDD.n1624 VDD.n290 0.00239394
R2833 VDD.n1600 VDD.n1599 0.00239394
R2834 VDD.n1590 VDD.n314 0.00239394
R2835 VDD.n1566 VDD.n1565 0.00239394
R2836 VDD.n1553 VDD.n340 0.00239394
R2837 VDD.n1541 VDD.n366 0.00239394
R2838 VDD.n1529 VDD.n382 0.00239394
R2839 VDD.n1517 VDD.n398 0.00239394
R2840 VDD.n1505 VDD.n414 0.00239394
R2841 VDD.n1491 VDD.n428 0.00239394
R2842 VDD.n1482 VDD.n436 0.00239394
R2843 VDD.n1471 VDD.n1470 0.00239394
R2844 VDD.n1461 VDD.n467 0.00239394
R2845 VDD.n1437 VDD.n1436 0.00239394
R2846 VDD.n1427 VDD.n491 0.00239394
R2847 VDD.n1403 VDD.n1402 0.00239394
R2848 VDD.n1390 VDD.n517 0.00239394
R2849 VDD.n1378 VDD.n543 0.00239394
R2850 VDD.n1366 VDD.n559 0.00239394
R2851 VDD.n1354 VDD.n575 0.00239394
R2852 VDD.n1342 VDD.n591 0.00239394
R2853 VDD.n1328 VDD.n605 0.00239394
R2854 VDD.n1319 VDD.n613 0.00239394
R2855 VDD.n1308 VDD.n1307 0.00239394
R2856 VDD.n1298 VDD.n644 0.00239394
R2857 VDD.n1274 VDD.n1273 0.00239394
R2858 VDD.n1264 VDD.n668 0.00239394
R2859 VDD.n1240 VDD.n1239 0.00239394
R2860 VDD.n1227 VDD.n694 0.00239394
R2861 VDD.n1215 VDD.n720 0.00239394
R2862 VDD.n1203 VDD.n736 0.00239394
R2863 VDD.n1191 VDD.n752 0.00239394
R2864 VDD.n1179 VDD.n768 0.00239394
R2865 VDD.n1165 VDD.n782 0.00239394
R2866 VDD.n1156 VDD.n790 0.00239394
R2867 VDD.n1145 VDD.n1144 0.00239394
R2868 VDD.n1135 VDD.n821 0.00239394
R2869 VDD.n1111 VDD.n1110 0.00239394
R2870 VDD.n1101 VDD.n845 0.00239394
R2871 VDD.n1077 VDD.n1076 0.00239394
R2872 VDD.n1058 VDD.n874 0.00239394
R2873 VDD.n1047 VDD.n1046 0.00239394
R2874 VDD.n1037 VDD.n913 0.00239394
R2875 VDD.n1026 VDD.n1025 0.00239394
R2876 VDD.n1016 VDD.n952 0.00239394
R2877 VDD.n968 VDD.n961 0.00224074
R2878 VDD.n47 VDD.n44 0.0021514
R2879 VDD.n970 VDD.n960 0.00213953
R2880 VDD.n1727 VDD.n11 0.00196875
R2881 VDD.n16 VDD.n13 0.00196875
R2882 VDD VDD.n1694 0.00170513
R2883 VDD.n1557 VDD 0.00170513
R2884 VDD.n1394 VDD 0.00170513
R2885 VDD.n1231 VDD 0.00170513
R2886 VDD.n175 VDD.n67 0.00119118
R2887 VDD.n176 VDD.n175 0.00119118
R2888 VDD.n191 VDD.n172 0.00119118
R2889 VDD.n192 VDD.n191 0.00119118
R2890 VDD.n211 VDD.n162 0.00119118
R2891 VDD.n212 VDD.n211 0.00119118
R2892 VDD.n1677 VDD.n160 0.00119118
R2893 VDD.n217 VDD.n160 0.00119118
R2894 VDD.n245 VDD.n218 0.00119118
R2895 VDD.n246 VDD.n245 0.00119118
R2896 VDD.n1656 VDD.n242 0.00119118
R2897 VDD.n252 VDD.n242 0.00119118
R2898 VDD.n277 VDD.n270 0.00119118
R2899 VDD.n278 VDD.n277 0.00119118
R2900 VDD.n1632 VDD.n1631 0.00119118
R2901 VDD.n1631 VDD.n268 0.00119118
R2902 VDD.n1625 VDD.n289 0.00119118
R2903 VDD.n304 VDD.n289 0.00119118
R2904 VDD.n1598 VDD.n1597 0.00119118
R2905 VDD.n1597 VDD.n301 0.00119118
R2906 VDD.n1591 VDD.n313 0.00119118
R2907 VDD.n328 VDD.n313 0.00119118
R2908 VDD.n1564 VDD.n1563 0.00119118
R2909 VDD.n1563 VDD.n325 0.00119118
R2910 VDD.n1555 VDD.n338 0.00119118
R2911 VDD.n341 VDD.n338 0.00119118
R2912 VDD.n1543 VDD.n361 0.00119118
R2913 VDD.n367 VDD.n361 0.00119118
R2914 VDD.n1531 VDD.n376 0.00119118
R2915 VDD.n383 VDD.n376 0.00119118
R2916 VDD.n1519 VDD.n392 0.00119118
R2917 VDD.n399 VDD.n392 0.00119118
R2918 VDD.n1507 VDD.n408 0.00119118
R2919 VDD.n415 VDD.n408 0.00119118
R2920 VDD.n1493 VDD.n422 0.00119118
R2921 VDD.n429 VDD.n422 0.00119118
R2922 VDD.n454 VDD.n447 0.00119118
R2923 VDD.n455 VDD.n454 0.00119118
R2924 VDD.n1469 VDD.n1468 0.00119118
R2925 VDD.n1468 VDD.n445 0.00119118
R2926 VDD.n1462 VDD.n466 0.00119118
R2927 VDD.n481 VDD.n466 0.00119118
R2928 VDD.n1435 VDD.n1434 0.00119118
R2929 VDD.n1434 VDD.n478 0.00119118
R2930 VDD.n1428 VDD.n490 0.00119118
R2931 VDD.n505 VDD.n490 0.00119118
R2932 VDD.n1401 VDD.n1400 0.00119118
R2933 VDD.n1400 VDD.n502 0.00119118
R2934 VDD.n1392 VDD.n515 0.00119118
R2935 VDD.n518 VDD.n515 0.00119118
R2936 VDD.n1380 VDD.n538 0.00119118
R2937 VDD.n544 VDD.n538 0.00119118
R2938 VDD.n1368 VDD.n553 0.00119118
R2939 VDD.n560 VDD.n553 0.00119118
R2940 VDD.n1356 VDD.n569 0.00119118
R2941 VDD.n576 VDD.n569 0.00119118
R2942 VDD.n1344 VDD.n585 0.00119118
R2943 VDD.n592 VDD.n585 0.00119118
R2944 VDD.n1330 VDD.n599 0.00119118
R2945 VDD.n606 VDD.n599 0.00119118
R2946 VDD.n631 VDD.n624 0.00119118
R2947 VDD.n632 VDD.n631 0.00119118
R2948 VDD.n1306 VDD.n1305 0.00119118
R2949 VDD.n1305 VDD.n622 0.00119118
R2950 VDD.n1299 VDD.n643 0.00119118
R2951 VDD.n658 VDD.n643 0.00119118
R2952 VDD.n1272 VDD.n1271 0.00119118
R2953 VDD.n1271 VDD.n655 0.00119118
R2954 VDD.n1265 VDD.n667 0.00119118
R2955 VDD.n682 VDD.n667 0.00119118
R2956 VDD.n1238 VDD.n1237 0.00119118
R2957 VDD.n1237 VDD.n679 0.00119118
R2958 VDD.n1229 VDD.n692 0.00119118
R2959 VDD.n695 VDD.n692 0.00119118
R2960 VDD.n1217 VDD.n715 0.00119118
R2961 VDD.n721 VDD.n715 0.00119118
R2962 VDD.n1205 VDD.n730 0.00119118
R2963 VDD.n737 VDD.n730 0.00119118
R2964 VDD.n1193 VDD.n746 0.00119118
R2965 VDD.n753 VDD.n746 0.00119118
R2966 VDD.n1181 VDD.n762 0.00119118
R2967 VDD.n769 VDD.n762 0.00119118
R2968 VDD.n1167 VDD.n776 0.00119118
R2969 VDD.n783 VDD.n776 0.00119118
R2970 VDD.n808 VDD.n801 0.00119118
R2971 VDD.n809 VDD.n808 0.00119118
R2972 VDD.n1143 VDD.n1142 0.00119118
R2973 VDD.n1142 VDD.n799 0.00119118
R2974 VDD.n1136 VDD.n820 0.00119118
R2975 VDD.n835 VDD.n820 0.00119118
R2976 VDD.n1109 VDD.n1108 0.00119118
R2977 VDD.n1108 VDD.n832 0.00119118
R2978 VDD.n1102 VDD.n844 0.00119118
R2979 VDD.n860 VDD.n844 0.00119118
R2980 VDD.n1075 VDD.n1074 0.00119118
R2981 VDD.n1074 VDD.n857 0.00119118
R2982 VDD.n1067 VDD.n868 0.00119118
R2983 VDD.n1064 VDD.n868 0.00119118
R2984 VDD.n1059 VDD.n873 0.00119118
R2985 VDD.n903 VDD.n873 0.00119118
R2986 VDD.n1045 VDD.n1044 0.00119118
R2987 VDD.n1044 VDD.n900 0.00119118
R2988 VDD.n1038 VDD.n912 0.00119118
R2989 VDD.n942 VDD.n912 0.00119118
R2990 VDD.n1024 VDD.n1023 0.00119118
R2991 VDD.n1023 VDD.n939 0.00119118
R2992 VDD.n1017 VDD.n951 0.00119118
R2993 VDD.n966 VDD.n951 0.00119118
R2994 VDD.n37 VDD.n35 0.0011215
R2995 VDD.n174 VDD.n66 0.00110256
R2996 VDD.n190 VDD.n189 0.00110256
R2997 VDD.n210 VDD.n209 0.00110256
R2998 VDD.n1676 VDD.n1675 0.00110256
R2999 VDD.n244 VDD.n243 0.00110256
R3000 VDD.n271 VDD.n250 0.00110256
R3001 VDD.n276 VDD.n269 0.00110256
R3002 VDD.n1630 VDD.n1629 0.00110256
R3003 VDD.n303 VDD.n302 0.00110256
R3004 VDD.n1596 VDD.n1595 0.00110256
R3005 VDD.n327 VDD.n326 0.00110256
R3006 VDD.n1562 VDD.n1561 0.00110256
R3007 VDD.n1556 VDD.n337 0.00110256
R3008 VDD.n377 VDD.n365 0.00110256
R3009 VDD.n393 VDD.n381 0.00110256
R3010 VDD.n409 VDD.n397 0.00110256
R3011 VDD.n423 VDD.n413 0.00110256
R3012 VDD.n448 VDD.n427 0.00110256
R3013 VDD.n453 VDD.n446 0.00110256
R3014 VDD.n1467 VDD.n1466 0.00110256
R3015 VDD.n480 VDD.n479 0.00110256
R3016 VDD.n1433 VDD.n1432 0.00110256
R3017 VDD.n504 VDD.n503 0.00110256
R3018 VDD.n1399 VDD.n1398 0.00110256
R3019 VDD.n1393 VDD.n514 0.00110256
R3020 VDD.n554 VDD.n542 0.00110256
R3021 VDD.n570 VDD.n558 0.00110256
R3022 VDD.n586 VDD.n574 0.00110256
R3023 VDD.n600 VDD.n590 0.00110256
R3024 VDD.n625 VDD.n604 0.00110256
R3025 VDD.n630 VDD.n623 0.00110256
R3026 VDD.n1304 VDD.n1303 0.00110256
R3027 VDD.n657 VDD.n656 0.00110256
R3028 VDD.n1270 VDD.n1269 0.00110256
R3029 VDD.n681 VDD.n680 0.00110256
R3030 VDD.n1236 VDD.n1235 0.00110256
R3031 VDD.n1230 VDD.n691 0.00110256
R3032 VDD.n731 VDD.n719 0.00110256
R3033 VDD.n747 VDD.n735 0.00110256
R3034 VDD.n763 VDD.n751 0.00110256
R3035 VDD.n777 VDD.n767 0.00110256
R3036 VDD.n802 VDD.n781 0.00110256
R3037 VDD.n807 VDD.n800 0.00110256
R3038 VDD.n1141 VDD.n1140 0.00110256
R3039 VDD.n834 VDD.n833 0.00110256
R3040 VDD.n1107 VDD.n1106 0.00110256
R3041 VDD.n859 VDD.n858 0.00110256
R3042 VDD.n1073 VDD.n1072 0.00110256
R3043 VDD.n1063 VDD.n867 0.00108025
R3044 VDD.n902 VDD.n901 0.00108025
R3045 VDD.n1043 VDD.n1042 0.00108025
R3046 VDD.n941 VDD.n940 0.00108025
R3047 VDD.n1022 VDD.n1021 0.00108025
R3048 VDD.n967 VDD.n965 0.00108025
R3049 VDD.n1729 VDD.n1728 0.000837321
R3050 VDD VDD.n22 0.00072488
R3051 VDD.n1729 VDD.n22 0.00061244
R3052 code[2] code[2].t1 140.387
R3053 code[2].n1 code[2].t2 140.34
R3054 code[2].n0 code[2].t0 140.34
R3055 code[2].n2 code[2].t3 140.34
R3056 code[2].n2 code[2] 2.82659
R3057 code[2].n1 code[2] 0.285826
R3058 code[2].n2 code[2].n0 0.264087
R3059 code[2].n0 code[2] 0.0466957
R3060 code[2] code[2].n1 0.0466957
R3061 code[2] code[2].n2 0.0371379
R3062 VSS.n616 VSS.n615 1272.41
R3063 VSS.n663 VSS 1043.16
R3064 VSS.n689 VSS.t11 641.946
R3065 VSS.n617 VSS.n616 626.532
R3066 VSS.n616 VSS.t3 621.635
R3067 VSS.n566 VSS.t1 359.05
R3068 VSS.n689 VSS 320.974
R3069 VSS.n691 VSS.n690 292.5
R3070 VSS.n690 VSS.n689 292.5
R3071 VSS.t3 VSS.t4 233.113
R3072 VSS.n641 VSS.n640 200.608
R3073 VSS.n665 VSS.n664 173.861
R3074 VSS.n665 VSS.t7 147.113
R3075 VSS.n567 VSS.n566 126.269
R3076 VSS.t1 VSS.t9 112.822
R3077 VSS.n691 VSS.t12 107.195
R3078 VSS.n658 VSS.t8 107.195
R3079 VSS.n642 VSS.n638 93.0283
R3080 VSS.n530 VSS.t6 77.3934
R3081 VSS.n530 VSS.t5 77.3934
R3082 VSS.n666 VSS.n662 71.1394
R3083 VSS.n664 VSS.n663 53.4959
R3084 VSS.n541 VSS.t2 43.7547
R3085 VSS.n617 VSS.t10 41.4448
R3086 VSS.n640 VSS.n639 26.7482
R3087 VSS.n662 VSS.n661 21.8894
R3088 VSS.n45 VSS.n44 17.6402
R3089 VSS.n256 VSS.n59 17.6402
R3090 VSS.n89 VSS.n88 17.6402
R3091 VSS.n329 VSS.n328 17.6402
R3092 VSS.n198 VSS.n52 17.6397
R3093 VSS.n74 VSS.n73 17.6397
R3094 VSS.n289 VSS.n288 17.6397
R3095 VSS.n429 VSS.n428 17.6397
R3096 VSS.n557 VSS.n556 17.6348
R3097 VSS.n481 VSS.n454 17.6348
R3098 VSS.n399 VSS.n314 17.6348
R3099 VSS.n667 VSS.n666 9.3005
R3100 VSS.n666 VSS.n665 9.3005
R3101 VSS.n655 VSS.n654 9.3005
R3102 VSS.n653 VSS.n652 9.3005
R3103 VSS.n561 VSS.n560 9.15497
R3104 VSS.n51 VSS.n50 9.15497
R3105 VSS.n36 VSS.n35 9.15497
R3106 VSS.n65 VSS.n64 9.15497
R3107 VSS.n58 VSS.n57 9.15497
R3108 VSS.n95 VSS.n94 9.15497
R3109 VSS.n80 VSS.n79 9.15497
R3110 VSS.n29 VSS.n28 9.15497
R3111 VSS.n303 VSS.n302 9.15497
R3112 VSS.n558 VSS.n303 9.15497
R3113 VSS.n313 VSS.n312 9.15497
R3114 VSS.n335 VSS.n334 9.15497
R3115 VSS.n320 VSS.n319 9.15497
R3116 VSS.n22 VSS.n21 9.15497
R3117 VSS.n443 VSS.n442 9.15497
R3118 VSS.n558 VSS.n443 9.15497
R3119 VSS.n453 VSS.n452 9.15497
R3120 VSS.n15 VSS.n14 9.15497
R3121 VSS.n501 VSS.n500 9.15497
R3122 VSS.n558 VSS.n501 9.15497
R3123 VSS.n511 VSS.n510 9.15497
R3124 VSS.n569 VSS.n568 9.15497
R3125 VSS.n568 VSS.n567 9.15497
R3126 VSS.n614 VSS.n613 9.15497
R3127 VSS.n615 VSS.n614 9.15497
R3128 VSS.n643 VSS.n642 9.01392
R3129 VSS.n642 VSS.n641 9.01392
R3130 VSS.n314 VSS.n313 8.61509
R3131 VSS.n454 VSS.n453 8.61509
R3132 VSS.n557 VSS.n511 8.61509
R3133 VSS.n52 VSS.n51 8.48617
R3134 VSS.n74 VSS.n65 8.48617
R3135 VSS.n289 VSS.n95 8.48617
R3136 VSS.n429 VSS.n335 8.48617
R3137 VSS.n45 VSS.n36 8.48574
R3138 VSS.n59 VSS.n58 8.48574
R3139 VSS.n89 VSS.n80 8.48574
R3140 VSS.n329 VSS.n320 8.48574
R3141 VSS.n560 VSS.n559 8.48521
R3142 VSS VSS.n691 7.93155
R3143 VSS.n659 VSS.n658 7.52991
R3144 VSS.n558 VSS.n30 6.48513
R3145 VSS.n558 VSS.n23 6.48513
R3146 VSS.n558 VSS.n16 6.48513
R3147 VSS.n633 VSS.n632 4.6505
R3148 VSS.n669 VSS.n668 4.5005
R3149 VSS.n668 VSS.n657 3.76521
R3150 VSS.n643 VSS.n637 3.45447
R3151 VSS.n660 VSS.n659 3.38874
R3152 VSS.n644 VSS.n636 3.25129
R3153 VSS.n400 VSS.n399 3.03311
R3154 VSS.n94 VSS.n93 3.03311
R3155 VSS.n64 VSS.n63 3.03311
R3156 VSS.n50 VSS.n49 3.03311
R3157 VSS.n482 VSS.n481 3.03311
R3158 VSS.n334 VSS.n333 3.03311
R3159 VSS.n556 VSS.n555 3.03311
R3160 VSS.n156 VSS.n153 3.03311
R3161 VSS.n562 VSS.n561 3.03311
R3162 VSS.n35 VSS.n34 3.03311
R3163 VSS.n44 VSS.n43 3.03311
R3164 VSS.n199 VSS.n198 3.03311
R3165 VSS.n57 VSS.n56 3.03311
R3166 VSS.n257 VSS.n256 3.03311
R3167 VSS.n73 VSS.n72 3.03311
R3168 VSS.n79 VSS.n78 3.03311
R3169 VSS.n88 VSS.n87 3.03311
R3170 VSS.n288 VSS.n287 3.03311
R3171 VSS.n28 VSS.n27 3.03311
R3172 VSS.n302 VSS.n301 3.03311
R3173 VSS.n312 VSS.n311 3.03311
R3174 VSS.n319 VSS.n318 3.03311
R3175 VSS.n328 VSS.n327 3.03311
R3176 VSS.n428 VSS.n427 3.03311
R3177 VSS.n21 VSS.n20 3.03311
R3178 VSS.n442 VSS.n441 3.03311
R3179 VSS.n452 VSS.n451 3.03311
R3180 VSS.n14 VSS.n13 3.03311
R3181 VSS.n500 VSS.n499 3.03311
R3182 VSS.n510 VSS.n509 3.03311
R3183 VSS.n570 VSS.n569 3.03311
R3184 VSS.n613 VSS.n612 3.03311
R3185 VSS.n645 VSS.n644 3.03311
R3186 VSS.n667 VSS.n660 3.01226
R3187 VSS.n16 VSS.n15 2.56987
R3188 VSS.n23 VSS.n22 2.56987
R3189 VSS.n30 VSS.n29 2.56987
R3190 VSS.n620 VSS.n619 2.24031
R3191 VSS.n621 VSS 1.94963
R3192 VSS.n668 VSS.n667 1.50638
R3193 VSS.n650 VSS.n649 1.35607
R3194 VSS.n674 VSS.n673 1.35607
R3195 VSS.n42 VSS.n41 1.35607
R3196 VSS.n71 VSS.n70 1.35607
R3197 VSS.n86 VSS.n85 1.35607
R3198 VSS.n310 VSS.n309 1.35607
R3199 VSS.n404 VSS.n403 1.35607
R3200 VSS.n326 VSS.n325 1.35607
R3201 VSS.n450 VSS.n449 1.35607
R3202 VSS.n486 VSS.n485 1.35607
R3203 VSS.n508 VSS.n507 1.35607
R3204 VSS.n554 VSS.n553 1.35607
R3205 VSS.n611 VSS.n610 1.35607
R3206 VSS.n688 VSS.n687 1.35607
R3207 VSS.n543 VSS.n542 1.13981
R3208 VSS.n301 VSS.n300 1.04008
R3209 VSS.n258 VSS.n257 1.04008
R3210 VSS.n441 VSS.n440 1.04008
R3211 VSS.n499 VSS.n498 1.04008
R3212 VSS.n157 VSS.n156 1.03985
R3213 VSS.n287 VSS.n285 1.03985
R3214 VSS.n200 VSS.n199 1.03985
R3215 VSS.n427 VSS.n425 1.03985
R3216 VSS.n497 VSS.n496 0.853
R3217 VSS.n535 VSS.n533 0.853
R3218 VSS.n496 VSS.n495 0.853
R3219 VSS.n553 VSS.n552 0.853
R3220 VSS.n552 VSS.n551 0.853
R3221 VSS.n491 VSS.n486 0.853
R3222 VSS.n423 VSS.n422 0.853
R3223 VSS.n424 VSS.n423 0.853
R3224 VSS.n388 VSS.n387 0.853
R3225 VSS.n492 VSS.n491 0.853
R3226 VSS.n409 VSS.n404 0.853
R3227 VSS.n218 VSS.n217 0.853
R3228 VSS.n217 VSS.n216 0.853
R3229 VSS.n261 VSS.n260 0.853
R3230 VSS.n260 VSS.n259 0.853
R3231 VSS.n283 VSS.n282 0.853
R3232 VSS.n284 VSS.n283 0.853
R3233 VSS.n149 VSS.n148 0.853
R3234 VSS.n410 VSS.n409 0.853
R3235 VSS.n623 VSS.n621 0.853
R3236 VSS.n624 VSS.n623 0.853
R3237 VSS.n609 VSS.n608 0.853
R3238 VSS.n166 VSS.n165 0.853
R3239 VSS.n167 VSS.n166 0.853
R3240 VSS.n610 VSS.n609 0.853
R3241 VSS.n676 VSS.n674 0.853
R3242 VSS.n687 VSS.n686 0.853
R3243 VSS.t9 VSS.t0 0.824007
R3244 VSS.n629 VSS.n628 0.699777
R3245 VSS.n537 VSS.n536 0.698382
R3246 VSS.n542 VSS.n541 0.684595
R3247 VSS.n538 VSS.n537 0.352759
R3248 VSS.n558 VSS.n314 0.341248
R3249 VSS.n558 VSS.n454 0.341248
R3250 VSS.n558 VSS.n557 0.341248
R3251 VSS.n558 VSS.n45 0.33661
R3252 VSS.n558 VSS.n59 0.33661
R3253 VSS.n558 VSS.n89 0.33661
R3254 VSS.n558 VSS.n329 0.33661
R3255 VSS.n559 VSS.n558 0.336142
R3256 VSS.n558 VSS.n52 0.336142
R3257 VSS.n558 VSS.n74 0.336142
R3258 VSS.n558 VSS.n289 0.336142
R3259 VSS.n558 VSS.n429 0.336142
R3260 VSS.n545 VSS.n544 0.280638
R3261 VSS.n146 VSS.n145 0.212
R3262 VSS.n385 VSS.n384 0.212
R3263 VSS.n644 VSS.n643 0.203675
R3264 VSS VSS.n6 0.177439
R3265 VSS.n627 VSS.n626 0.17525
R3266 VSS VSS.n493 0.148517
R3267 VSS VSS.n411 0.147312
R3268 VSS VSS.n168 0.147312
R3269 VSS.n626 VSS.n625 0.129277
R3270 VSS.n494 VSS 0.111158
R3271 VSS VSS.n389 0.111158
R3272 VSS.n412 VSS 0.111158
R3273 VSS VSS.n150 0.111158
R3274 VSS.n272 VSS 0.111158
R3275 VSS.n220 VSS 0.111158
R3276 VSS.n169 VSS 0.111158
R3277 VSS.n607 VSS 0.111158
R3278 VSS.n618 VSS 0.104812
R3279 VSS.n634 VSS.n633 0.0929479
R3280 VSS.n672 VSS.n671 0.0734167
R3281 VSS.n390 VSS 0.0718924
R3282 VSS.n151 VSS 0.0718924
R3283 VSS VSS.n271 0.0718924
R3284 VSS VSS.n219 0.0718924
R3285 VSS.n402 VSS.n401 0.0685147
R3286 VSS.n305 VSS.n304 0.0685147
R3287 VSS.n25 VSS.n24 0.0685147
R3288 VSS.n484 VSS.n483 0.0685147
R3289 VSS.n445 VSS.n444 0.0685147
R3290 VSS.n18 VSS.n17 0.0685147
R3291 VSS.n513 VSS.n512 0.0685147
R3292 VSS.n503 VSS.n502 0.0685147
R3293 VSS.n11 VSS.n10 0.0685147
R3294 VSS.n155 VSS.n154 0.0685147
R3295 VSS.n564 VSS.n563 0.0685147
R3296 VSS.n572 VSS.n571 0.0685147
R3297 VSS.n633 VSS.n0 0.0643021
R3298 VSS.n653 VSS 0.0512812
R3299 VSS.n628 VSS.n627 0.0498797
R3300 VSS.n162 VSS.n161 0.0482941
R3301 VSS.n575 VSS.n574 0.0482941
R3302 VSS.n581 VSS.n580 0.0482941
R3303 VSS.n397 VSS.n396 0.0482941
R3304 VSS.n296 VSS.n295 0.0482941
R3305 VSS.n108 VSS.n107 0.0482941
R3306 VSS.n102 VSS.n101 0.0482941
R3307 VSS.n246 VSS.n245 0.0482941
R3308 VSS.n252 VSS.n251 0.0482941
R3309 VSS.n213 VSS.n212 0.0482941
R3310 VSS.n207 VSS.n206 0.0482941
R3311 VSS.n479 VSS.n478 0.0482941
R3312 VSS.n436 VSS.n435 0.0482941
R3313 VSS.n348 VSS.n347 0.0482941
R3314 VSS.n342 VSS.n341 0.0482941
R3315 VSS.n517 VSS.n516 0.0482941
R3316 VSS.n461 VSS.n460 0.0482941
R3317 VSS.n687 VSS.n1 0.0427297
R3318 VSS.n533 VSS.n529 0.0415156
R3319 VSS.n621 VSS.n8 0.0415156
R3320 VSS.n684 VSS.n683 0.0411354
R3321 VSS.n164 VSS.n163 0.0391029
R3322 VSS.n160 VSS.n159 0.0391029
R3323 VSS.n577 VSS.n576 0.0391029
R3324 VSS.n579 VSS.n578 0.0391029
R3325 VSS.n610 VSS.n582 0.0391029
R3326 VSS.n403 VSS.n402 0.0391029
R3327 VSS.n310 VSS.n305 0.0391029
R3328 VSS.n26 VSS.n25 0.0391029
R3329 VSS.n404 VSS.n398 0.0391029
R3330 VSS.n309 VSS.n308 0.0391029
R3331 VSS.n292 VSS.n291 0.0391029
R3332 VSS.n294 VSS.n293 0.0391029
R3333 VSS.n298 VSS.n297 0.0391029
R3334 VSS.n287 VSS.n286 0.0391029
R3335 VSS.n91 VSS.n90 0.0391029
R3336 VSS.n93 VSS.n92 0.0391029
R3337 VSS.n76 VSS.n75 0.0391029
R3338 VSS.n78 VSS.n77 0.0391029
R3339 VSS.n86 VSS.n81 0.0391029
R3340 VSS.n110 VSS.n109 0.0391029
R3341 VSS.n106 VSS.n105 0.0391029
R3342 VSS.n104 VSS.n103 0.0391029
R3343 VSS.n100 VSS.n99 0.0391029
R3344 VSS.n98 VSS.n97 0.0391029
R3345 VSS.n85 VSS.n83 0.0391029
R3346 VSS.n71 VSS.n66 0.0391029
R3347 VSS.n63 VSS.n60 0.0391029
R3348 VSS.n62 VSS.n61 0.0391029
R3349 VSS.n56 VSS.n53 0.0391029
R3350 VSS.n55 VSS.n54 0.0391029
R3351 VSS.n257 VSS.n255 0.0391029
R3352 VSS.n70 VSS.n69 0.0391029
R3353 VSS.n242 VSS.n241 0.0391029
R3354 VSS.n244 VSS.n243 0.0391029
R3355 VSS.n248 VSS.n247 0.0391029
R3356 VSS.n250 VSS.n249 0.0391029
R3357 VSS.n254 VSS.n253 0.0391029
R3358 VSS.n199 VSS.n197 0.0391029
R3359 VSS.n47 VSS.n46 0.0391029
R3360 VSS.n49 VSS.n48 0.0391029
R3361 VSS.n32 VSS.n31 0.0391029
R3362 VSS.n34 VSS.n33 0.0391029
R3363 VSS.n42 VSS.n37 0.0391029
R3364 VSS.n215 VSS.n214 0.0391029
R3365 VSS.n211 VSS.n210 0.0391029
R3366 VSS.n209 VSS.n208 0.0391029
R3367 VSS.n205 VSS.n204 0.0391029
R3368 VSS.n203 VSS.n202 0.0391029
R3369 VSS.n41 VSS.n39 0.0391029
R3370 VSS.n485 VSS.n484 0.0391029
R3371 VSS.n450 VSS.n445 0.0391029
R3372 VSS.n19 VSS.n18 0.0391029
R3373 VSS.n486 VSS.n480 0.0391029
R3374 VSS.n449 VSS.n448 0.0391029
R3375 VSS.n432 VSS.n431 0.0391029
R3376 VSS.n434 VSS.n433 0.0391029
R3377 VSS.n438 VSS.n437 0.0391029
R3378 VSS.n427 VSS.n426 0.0391029
R3379 VSS.n331 VSS.n330 0.0391029
R3380 VSS.n333 VSS.n332 0.0391029
R3381 VSS.n316 VSS.n315 0.0391029
R3382 VSS.n318 VSS.n317 0.0391029
R3383 VSS.n326 VSS.n321 0.0391029
R3384 VSS.n350 VSS.n349 0.0391029
R3385 VSS.n346 VSS.n345 0.0391029
R3386 VSS.n344 VSS.n343 0.0391029
R3387 VSS.n340 VSS.n339 0.0391029
R3388 VSS.n338 VSS.n337 0.0391029
R3389 VSS.n325 VSS.n323 0.0391029
R3390 VSS.n554 VSS.n513 0.0391029
R3391 VSS.n508 VSS.n503 0.0391029
R3392 VSS.n12 VSS.n11 0.0391029
R3393 VSS.n553 VSS.n518 0.0391029
R3394 VSS.n507 VSS.n506 0.0391029
R3395 VSS.n457 VSS.n456 0.0391029
R3396 VSS.n459 VSS.n458 0.0391029
R3397 VSS.n463 VSS.n462 0.0391029
R3398 VSS.n156 VSS.n155 0.0391029
R3399 VSS.n154 VSS.n9 0.0391029
R3400 VSS.n563 VSS.n562 0.0391029
R3401 VSS.n565 VSS.n564 0.0391029
R3402 VSS.n571 VSS.n570 0.0391029
R3403 VSS.n611 VSS.n572 0.0391029
R3404 VSS.n4 VSS.n3 0.0361962
R3405 VSS.n647 VSS.n646 0.035973
R3406 VSS.n649 VSS.n648 0.035973
R3407 VSS VSS.n688 0.0330521
R3408 VSS.n674 VSS.n630 0.0325946
R3409 VSS VSS.n651 0.03175
R3410 VSS.n679 VSS.n678 0.029875
R3411 VSS.n651 VSS.n650 0.0278438
R3412 VSS.n619 VSS.n618 0.0257686
R3413 VSS.n531 VSS.n530 0.024008
R3414 VSS.n671 VSS 0.0226354
R3415 VSS.n621 VSS.n620 0.0223823
R3416 VSS.n610 VSS.n583 0.0219755
R3417 VSS.n404 VSS.n394 0.0219755
R3418 VSS.n85 VSS.n84 0.0219755
R3419 VSS.n70 VSS.n67 0.0219755
R3420 VSS.n41 VSS.n40 0.0219755
R3421 VSS.n486 VSS.n476 0.0219755
R3422 VSS.n325 VSS.n324 0.0219755
R3423 VSS.n553 VSS.n514 0.0219755
R3424 VSS.n645 VSS.n635 0.0213333
R3425 VSS.n673 VSS.n670 0.0200312
R3426 VSS.n409 VSS.n393 0.0191618
R3427 VSS.n409 VSS.n408 0.0191618
R3428 VSS.n136 VSS.n135 0.0191618
R3429 VSS.n140 VSS.n139 0.0191618
R3430 VSS.n141 VSS.n140 0.0191618
R3431 VSS.n148 VSS.n144 0.0191618
R3432 VSS.n148 VSS.n147 0.0191618
R3433 VSS.n283 VSS.n111 0.0191618
R3434 VSS.n283 VSS.n128 0.0191618
R3435 VSS.n125 VSS.n124 0.0191618
R3436 VSS.n124 VSS.n123 0.0191618
R3437 VSS.n120 VSS.n119 0.0191618
R3438 VSS.n119 VSS.n118 0.0191618
R3439 VSS.n115 VSS.n114 0.0191618
R3440 VSS.n114 VSS.n113 0.0191618
R3441 VSS.n223 VSS.n222 0.0191618
R3442 VSS.n224 VSS.n223 0.0191618
R3443 VSS.n228 VSS.n227 0.0191618
R3444 VSS.n229 VSS.n228 0.0191618
R3445 VSS.n233 VSS.n232 0.0191618
R3446 VSS.n234 VSS.n233 0.0191618
R3447 VSS.n260 VSS.n237 0.0191618
R3448 VSS.n260 VSS.n239 0.0191618
R3449 VSS.n217 VSS.n180 0.0191618
R3450 VSS.n217 VSS.n196 0.0191618
R3451 VSS.n193 VSS.n192 0.0191618
R3452 VSS.n192 VSS.n191 0.0191618
R3453 VSS.n188 VSS.n187 0.0191618
R3454 VSS.n187 VSS.n186 0.0191618
R3455 VSS.n183 VSS.n182 0.0191618
R3456 VSS.n182 VSS.n181 0.0191618
R3457 VSS.n491 VSS.n475 0.0191618
R3458 VSS.n491 VSS.n490 0.0191618
R3459 VSS.n375 VSS.n374 0.0191618
R3460 VSS.n379 VSS.n378 0.0191618
R3461 VSS.n380 VSS.n379 0.0191618
R3462 VSS.n387 VSS.n383 0.0191618
R3463 VSS.n387 VSS.n386 0.0191618
R3464 VSS.n423 VSS.n351 0.0191618
R3465 VSS.n423 VSS.n367 0.0191618
R3466 VSS.n364 VSS.n363 0.0191618
R3467 VSS.n363 VSS.n362 0.0191618
R3468 VSS.n359 VSS.n358 0.0191618
R3469 VSS.n358 VSS.n357 0.0191618
R3470 VSS.n354 VSS.n353 0.0191618
R3471 VSS.n353 VSS.n352 0.0191618
R3472 VSS.n552 VSS.n519 0.0191618
R3473 VSS.n552 VSS.n528 0.0191618
R3474 VSS.n525 VSS.n524 0.0191618
R3475 VSS.n524 VSS.n523 0.0191618
R3476 VSS.n465 VSS.n464 0.0191618
R3477 VSS.n496 VSS.n468 0.0191618
R3478 VSS.n496 VSS.n469 0.0191618
R3479 VSS.n166 VSS.n152 0.0191618
R3480 VSS.n588 VSS.n587 0.0191618
R3481 VSS.n589 VSS.n588 0.0191618
R3482 VSS.n593 VSS.n592 0.0191618
R3483 VSS.n594 VSS.n593 0.0191618
R3484 VSS.n609 VSS.n597 0.0191618
R3485 VSS.n609 VSS.n598 0.0191618
R3486 VSS.n551 VSS.n545 0.0183481
R3487 VSS.n551 VSS.n550 0.0183481
R3488 VSS.n549 VSS.n548 0.0183481
R3489 VSS.n548 VSS.n547 0.0183481
R3490 VSS.n471 VSS.n470 0.0183481
R3491 VSS.n495 VSS.n472 0.0183481
R3492 VSS.n495 VSS.n494 0.0183481
R3493 VSS.n493 VSS.n492 0.0183481
R3494 VSS.n492 VSS.n474 0.0183481
R3495 VSS.n369 VSS.n368 0.0183481
R3496 VSS.n371 VSS.n370 0.0183481
R3497 VSS.n372 VSS.n371 0.0183481
R3498 VSS.n388 VSS.n373 0.0183481
R3499 VSS.n389 VSS.n388 0.0183481
R3500 VSS.n422 VSS.n390 0.0183481
R3501 VSS.n422 VSS.n421 0.0183481
R3502 VSS.n420 VSS.n419 0.0183481
R3503 VSS.n419 VSS.n418 0.0183481
R3504 VSS.n417 VSS.n416 0.0183481
R3505 VSS.n416 VSS.n415 0.0183481
R3506 VSS.n414 VSS.n413 0.0183481
R3507 VSS.n413 VSS.n412 0.0183481
R3508 VSS.n411 VSS.n410 0.0183481
R3509 VSS.n410 VSS.n392 0.0183481
R3510 VSS.n130 VSS.n129 0.0183481
R3511 VSS.n132 VSS.n131 0.0183481
R3512 VSS.n133 VSS.n132 0.0183481
R3513 VSS.n149 VSS.n134 0.0183481
R3514 VSS.n150 VSS.n149 0.0183481
R3515 VSS.n282 VSS.n151 0.0183481
R3516 VSS.n282 VSS.n281 0.0183481
R3517 VSS.n280 VSS.n279 0.0183481
R3518 VSS.n279 VSS.n278 0.0183481
R3519 VSS.n277 VSS.n276 0.0183481
R3520 VSS.n276 VSS.n275 0.0183481
R3521 VSS.n274 VSS.n273 0.0183481
R3522 VSS.n273 VSS.n272 0.0183481
R3523 VSS.n271 VSS.n270 0.0183481
R3524 VSS.n270 VSS.n269 0.0183481
R3525 VSS.n268 VSS.n267 0.0183481
R3526 VSS.n267 VSS.n266 0.0183481
R3527 VSS.n265 VSS.n264 0.0183481
R3528 VSS.n264 VSS.n263 0.0183481
R3529 VSS.n262 VSS.n261 0.0183481
R3530 VSS.n261 VSS.n220 0.0183481
R3531 VSS.n219 VSS.n218 0.0183481
R3532 VSS.n218 VSS.n178 0.0183481
R3533 VSS.n177 VSS.n176 0.0183481
R3534 VSS.n176 VSS.n175 0.0183481
R3535 VSS.n174 VSS.n173 0.0183481
R3536 VSS.n173 VSS.n172 0.0183481
R3537 VSS.n171 VSS.n170 0.0183481
R3538 VSS.n170 VSS.n169 0.0183481
R3539 VSS.n168 VSS.n167 0.0183481
R3540 VSS.n601 VSS.n600 0.0183481
R3541 VSS.n602 VSS.n601 0.0183481
R3542 VSS.n604 VSS.n603 0.0183481
R3543 VSS.n605 VSS.n604 0.0183481
R3544 VSS.n608 VSS.n606 0.0183481
R3545 VSS.n608 VSS.n607 0.0183481
R3546 VSS.n627 VSS.n5 0.0183481
R3547 VSS.n5 VSS.n4 0.0183481
R3548 VSS.n624 VSS.n6 0.0172857
R3549 VSS.n625 VSS.n624 0.0172857
R3550 VSS.n540 VSS.n539 0.0156071
R3551 VSS.n535 VSS.n534 0.0156071
R3552 VSS.n623 VSS.n7 0.0156071
R3553 VSS.n623 VSS.n622 0.0156071
R3554 VSS.n407 VSS.n406 0.0143235
R3555 VSS.n138 VSS.n137 0.0143235
R3556 VSS.n143 VSS.n142 0.0143235
R3557 VSS.n127 VSS.n126 0.0143235
R3558 VSS.n122 VSS.n121 0.0143235
R3559 VSS.n117 VSS.n116 0.0143235
R3560 VSS.n226 VSS.n225 0.0143235
R3561 VSS.n231 VSS.n230 0.0143235
R3562 VSS.n236 VSS.n235 0.0143235
R3563 VSS.n195 VSS.n194 0.0143235
R3564 VSS.n190 VSS.n189 0.0143235
R3565 VSS.n185 VSS.n184 0.0143235
R3566 VSS.n489 VSS.n488 0.0143235
R3567 VSS.n377 VSS.n376 0.0143235
R3568 VSS.n382 VSS.n381 0.0143235
R3569 VSS.n366 VSS.n365 0.0143235
R3570 VSS.n361 VSS.n360 0.0143235
R3571 VSS.n356 VSS.n355 0.0143235
R3572 VSS.n527 VSS.n526 0.0143235
R3573 VSS.n522 VSS.n521 0.0143235
R3574 VSS.n467 VSS.n466 0.0143235
R3575 VSS.n586 VSS.n585 0.0143235
R3576 VSS.n591 VSS.n590 0.0143235
R3577 VSS.n596 VSS.n595 0.0143235
R3578 VSS.n618 VSS.n617 0.0142993
R3579 VSS.n532 VSS.n531 0.0137243
R3580 VSS.n686 VSS.n685 0.0137188
R3581 VSS.n682 VSS.n681 0.0137188
R3582 VSS.n681 VSS.n680 0.0137188
R3583 VSS.n677 VSS.n676 0.0137188
R3584 VSS.n669 VSS.n656 0.0135208
R3585 VSS.n550 VSS.n549 0.0123987
R3586 VSS.n547 VSS.n546 0.0123987
R3587 VSS.n472 VSS.n471 0.0123987
R3588 VSS.n474 VSS.n473 0.0123987
R3589 VSS.n370 VSS.n369 0.0123987
R3590 VSS.n373 VSS.n372 0.0123987
R3591 VSS.n421 VSS.n420 0.0123987
R3592 VSS.n418 VSS.n417 0.0123987
R3593 VSS.n415 VSS.n414 0.0123987
R3594 VSS.n392 VSS.n391 0.0123987
R3595 VSS.n131 VSS.n130 0.0123987
R3596 VSS.n134 VSS.n133 0.0123987
R3597 VSS.n281 VSS.n280 0.0123987
R3598 VSS.n278 VSS.n277 0.0123987
R3599 VSS.n275 VSS.n274 0.0123987
R3600 VSS.n269 VSS.n268 0.0123987
R3601 VSS.n266 VSS.n265 0.0123987
R3602 VSS.n263 VSS.n262 0.0123987
R3603 VSS.n178 VSS.n177 0.0123987
R3604 VSS.n175 VSS.n174 0.0123987
R3605 VSS.n172 VSS.n171 0.0123987
R3606 VSS.n600 VSS.n599 0.0123987
R3607 VSS.n603 VSS.n602 0.0123987
R3608 VSS.n606 VSS.n605 0.0123987
R3609 VSS.n674 VSS.n631 0.0123243
R3610 VSS.n619 VSS 0.0121822
R3611 VSS.n161 VSS.n160 0.0115294
R3612 VSS.n576 VSS.n575 0.0115294
R3613 VSS.n582 VSS.n581 0.0115294
R3614 VSS.n398 VSS.n397 0.0115294
R3615 VSS.n308 VSS.n307 0.0115294
R3616 VSS.n295 VSS.n294 0.0115294
R3617 VSS.n107 VSS.n106 0.0115294
R3618 VSS.n101 VSS.n100 0.0115294
R3619 VSS.n83 VSS.n82 0.0115294
R3620 VSS.n69 VSS.n68 0.0115294
R3621 VSS.n245 VSS.n244 0.0115294
R3622 VSS.n251 VSS.n250 0.0115294
R3623 VSS.n212 VSS.n211 0.0115294
R3624 VSS.n206 VSS.n205 0.0115294
R3625 VSS.n39 VSS.n38 0.0115294
R3626 VSS.n480 VSS.n479 0.0115294
R3627 VSS.n448 VSS.n447 0.0115294
R3628 VSS.n435 VSS.n434 0.0115294
R3629 VSS.n347 VSS.n346 0.0115294
R3630 VSS.n341 VSS.n340 0.0115294
R3631 VSS.n323 VSS.n322 0.0115294
R3632 VSS.n518 VSS.n517 0.0115294
R3633 VSS.n506 VSS.n505 0.0115294
R3634 VSS.n460 VSS.n459 0.0115294
R3635 VSS.n300 VSS.n299 0.0104679
R3636 VSS.n259 VSS.n258 0.0104679
R3637 VSS.n440 VSS.n439 0.0104679
R3638 VSS.n498 VSS.n497 0.0104679
R3639 VSS.n165 VSS.n157 0.0098203
R3640 VSS.n216 VSS.n200 0.0098203
R3641 VSS.n285 VSS.n284 0.0098203
R3642 VSS.n425 VSS.n424 0.0098203
R3643 VSS.n163 VSS.n162 0.00969118
R3644 VSS.n574 VSS.n573 0.00969118
R3645 VSS.n580 VSS.n579 0.00969118
R3646 VSS.n396 VSS.n395 0.00969118
R3647 VSS.n291 VSS.n290 0.00969118
R3648 VSS.n297 VSS.n296 0.00969118
R3649 VSS.n109 VSS.n108 0.00969118
R3650 VSS.n103 VSS.n102 0.00969118
R3651 VSS.n97 VSS.n96 0.00969118
R3652 VSS.n241 VSS.n240 0.00969118
R3653 VSS.n247 VSS.n246 0.00969118
R3654 VSS.n253 VSS.n252 0.00969118
R3655 VSS.n214 VSS.n213 0.00969118
R3656 VSS.n208 VSS.n207 0.00969118
R3657 VSS.n202 VSS.n201 0.00969118
R3658 VSS.n478 VSS.n477 0.00969118
R3659 VSS.n431 VSS.n430 0.00969118
R3660 VSS.n437 VSS.n436 0.00969118
R3661 VSS.n349 VSS.n348 0.00969118
R3662 VSS.n343 VSS.n342 0.00969118
R3663 VSS.n337 VSS.n336 0.00969118
R3664 VSS.n516 VSS.n515 0.00969118
R3665 VSS.n456 VSS.n455 0.00969118
R3666 VSS.n462 VSS.n461 0.00969118
R3667 VSS.n673 VSS.n672 0.00961458
R3668 VSS.n635 VSS.n634 0.00701042
R3669 VSS.n655 VSS.n653 0.00570833
R3670 VSS.n670 VSS.n669 0.00570833
R3671 VSS.n626 VSS 0.005375
R3672 VSS.n543 VSS.n538 0.00493396
R3673 VSS.n544 VSS.n543 0.00493396
R3674 VSS.n536 VSS.n535 0.00489326
R3675 VSS.n686 VSS.n629 0.00451955
R3676 VSS.n656 VSS.n655 0.00440625
R3677 VSS.n676 VSS.n675 0.00362372
R3678 VSS.n408 VSS.n407 0.00257353
R3679 VSS.n406 VSS.n405 0.00257353
R3680 VSS.n137 VSS.n136 0.00257353
R3681 VSS.n139 VSS.n138 0.00257353
R3682 VSS.n142 VSS.n141 0.00257353
R3683 VSS.n144 VSS.n143 0.00257353
R3684 VSS.n147 VSS.n146 0.00257353
R3685 VSS.n145 VSS.n111 0.00257353
R3686 VSS.n128 VSS.n127 0.00257353
R3687 VSS.n126 VSS.n125 0.00257353
R3688 VSS.n123 VSS.n122 0.00257353
R3689 VSS.n121 VSS.n120 0.00257353
R3690 VSS.n118 VSS.n117 0.00257353
R3691 VSS.n116 VSS.n115 0.00257353
R3692 VSS.n113 VSS.n112 0.00257353
R3693 VSS.n222 VSS.n221 0.00257353
R3694 VSS.n225 VSS.n224 0.00257353
R3695 VSS.n227 VSS.n226 0.00257353
R3696 VSS.n230 VSS.n229 0.00257353
R3697 VSS.n232 VSS.n231 0.00257353
R3698 VSS.n235 VSS.n234 0.00257353
R3699 VSS.n237 VSS.n236 0.00257353
R3700 VSS.n239 VSS.n238 0.00257353
R3701 VSS.n180 VSS.n179 0.00257353
R3702 VSS.n196 VSS.n195 0.00257353
R3703 VSS.n194 VSS.n193 0.00257353
R3704 VSS.n191 VSS.n190 0.00257353
R3705 VSS.n189 VSS.n188 0.00257353
R3706 VSS.n186 VSS.n185 0.00257353
R3707 VSS.n184 VSS.n183 0.00257353
R3708 VSS.n490 VSS.n489 0.00257353
R3709 VSS.n488 VSS.n487 0.00257353
R3710 VSS.n376 VSS.n375 0.00257353
R3711 VSS.n378 VSS.n377 0.00257353
R3712 VSS.n381 VSS.n380 0.00257353
R3713 VSS.n383 VSS.n382 0.00257353
R3714 VSS.n386 VSS.n385 0.00257353
R3715 VSS.n384 VSS.n351 0.00257353
R3716 VSS.n367 VSS.n366 0.00257353
R3717 VSS.n365 VSS.n364 0.00257353
R3718 VSS.n362 VSS.n361 0.00257353
R3719 VSS.n360 VSS.n359 0.00257353
R3720 VSS.n357 VSS.n356 0.00257353
R3721 VSS.n355 VSS.n354 0.00257353
R3722 VSS.n528 VSS.n527 0.00257353
R3723 VSS.n526 VSS.n525 0.00257353
R3724 VSS.n523 VSS.n522 0.00257353
R3725 VSS.n521 VSS.n520 0.00257353
R3726 VSS.n466 VSS.n465 0.00257353
R3727 VSS.n468 VSS.n467 0.00257353
R3728 VSS.n585 VSS.n584 0.00257353
R3729 VSS.n587 VSS.n586 0.00257353
R3730 VSS.n590 VSS.n589 0.00257353
R3731 VSS.n592 VSS.n591 0.00257353
R3732 VSS.n595 VSS.n594 0.00257353
R3733 VSS.n597 VSS.n596 0.00257353
R3734 VSS.n165 VSS.n164 0.00233824
R3735 VSS.n159 VSS.n158 0.00233824
R3736 VSS.n578 VSS.n577 0.00233824
R3737 VSS.n403 VSS.n400 0.00233824
R3738 VSS.n311 VSS.n310 0.00233824
R3739 VSS.n27 VSS.n26 0.00233824
R3740 VSS.n309 VSS.n306 0.00233824
R3741 VSS.n293 VSS.n292 0.00233824
R3742 VSS.n299 VSS.n298 0.00233824
R3743 VSS.n93 VSS.n91 0.00233824
R3744 VSS.n78 VSS.n76 0.00233824
R3745 VSS.n87 VSS.n86 0.00233824
R3746 VSS.n284 VSS.n110 0.00233824
R3747 VSS.n105 VSS.n104 0.00233824
R3748 VSS.n99 VSS.n98 0.00233824
R3749 VSS.n72 VSS.n71 0.00233824
R3750 VSS.n63 VSS.n62 0.00233824
R3751 VSS.n56 VSS.n55 0.00233824
R3752 VSS.n243 VSS.n242 0.00233824
R3753 VSS.n249 VSS.n248 0.00233824
R3754 VSS.n259 VSS.n254 0.00233824
R3755 VSS.n49 VSS.n47 0.00233824
R3756 VSS.n34 VSS.n32 0.00233824
R3757 VSS.n43 VSS.n42 0.00233824
R3758 VSS.n216 VSS.n215 0.00233824
R3759 VSS.n210 VSS.n209 0.00233824
R3760 VSS.n204 VSS.n203 0.00233824
R3761 VSS.n485 VSS.n482 0.00233824
R3762 VSS.n451 VSS.n450 0.00233824
R3763 VSS.n20 VSS.n19 0.00233824
R3764 VSS.n449 VSS.n446 0.00233824
R3765 VSS.n433 VSS.n432 0.00233824
R3766 VSS.n439 VSS.n438 0.00233824
R3767 VSS.n333 VSS.n331 0.00233824
R3768 VSS.n318 VSS.n316 0.00233824
R3769 VSS.n327 VSS.n326 0.00233824
R3770 VSS.n424 VSS.n350 0.00233824
R3771 VSS.n345 VSS.n344 0.00233824
R3772 VSS.n339 VSS.n338 0.00233824
R3773 VSS.n555 VSS.n554 0.00233824
R3774 VSS.n509 VSS.n508 0.00233824
R3775 VSS.n13 VSS.n12 0.00233824
R3776 VSS.n507 VSS.n504 0.00233824
R3777 VSS.n458 VSS.n457 0.00233824
R3778 VSS.n497 VSS.n463 0.00233824
R3779 VSS.n562 VSS.n9 0.00233824
R3780 VSS.n570 VSS.n565 0.00233824
R3781 VSS.n612 VSS.n611 0.00233824
R3782 VSS.n649 VSS.n647 0.00218919
R3783 VSS.n687 VSS.n2 0.00218919
R3784 VSS.n542 VSS.n540 0.0021514
R3785 VSS.n685 VSS.n684 0.00196875
R3786 VSS.n683 VSS.n682 0.00196875
R3787 VSS.n680 VSS.n679 0.00196875
R3788 VSS.n678 VSS.n677 0.00196875
R3789 VSS.n688 VSS.n0 0.00180208
R3790 VSS.n650 VSS.n645 0.00180208
R3791 VSS.n533 VSS.n532 0.0011215
R3792 code_offset.n2 code_offset.t1 230.016
R3793 code_offset.n1 code_offset.t2 153.665
R3794 code_offset.n2 code_offset 153.601
R3795 code_offset code_offset.t0 140.379
R3796 code_offset.n3 code_offset.n2 9.3005
R3797 code_offset.n2 code_offset.n1 4.91671
R3798 code_offset.n5 code_offset.n3 4.9013
R3799 code_offset.n4 code_offset 4.22092
R3800 code_offset code_offset.n0 2.4005
R3801 code_offset.n4 code_offset 1.01229
R3802 code_offset.n5 code_offset.n4 0.726043
R3803 code_offset.n3 code_offset.n0 0.533833
R3804 code_offset.n6 code_offset.n5 0.421696
R3805 code_offset code_offset.n6 0.0195217
R3806 code_offset.n6 code_offset 0.0170094
R3807 OUT.n2 OUT.t5 107.647
R3808 OUT.n1 OUT.t4 107.647
R3809 OUT.n2 OUT.t3 91.5805
R3810 OUT.n1 OUT.t2 91.5805
R3811 OUT.n0 OUT.t1 68.3658
R3812 OUT.n2 OUT.n1 58.5727
R3813 OUT.n0 OUT.t0 41.7552
R3814 OUT OUT.n2 13.4931
R3815 OUT OUT.n0 0.422914
R3816 code[1] code[1].t0 140.387
R3817 code[1].n0 code[1].t1 140.34
R3818 code[1].n0 code[1] 0.201587
R3819 code[1] code[1].n0 0.0371379
R3820 IN.t4 IN.t17 221.72
R3821 IN.t7 IN.t4 221.72
R3822 IN.t14 IN.t7 221.72
R3823 IN.t2 IN.t14 221.72
R3824 IN.t12 IN.t2 221.72
R3825 IN.t5 IN.t9 221.72
R3826 IN.t18 IN.t5 221.72
R3827 IN.t11 IN.t18 221.72
R3828 IN.t0 IN.t11 221.72
R3829 IN.t21 IN.t0 221.72
R3830 IN.t16 IN.t21 221.72
R3831 IN.t10 IN.t16 221.72
R3832 IN.t1 IN.t6 221.72
R3833 IN.t13 IN.t1 221.72
R3834 IN.t8 IN.t13 221.72
R3835 IN.t20 IN.t8 221.72
R3836 IN.t3 IN.t20 221.72
R3837 IN.t19 IN.t3 221.72
R3838 IN.t15 IN.t19 221.72
R3839 IN.n5 IN.t12 154.8
R3840 IN.n0 IN 89.9738
R3841 IN.n1 IN.t10 78.7272
R3842 IN.n0 IN.t15 74.6592
R3843 IN.n2 IN 40.1672
R3844 IN.n3 IN.n1 32.1338
R3845 IN IN.n1 21.4227
R3846 IN.n4 IN.n0 21.3547
R3847 IN.n4 IN.n3 17.8279
R3848 IN.n5 IN.n4 13.4163
R3849 IN.n2 IN 11.8854
R3850 IN.n3 IN.n2 3.96214
R3851 IN.n6 IN 1.64944
R3852 IN.n6 IN 0.10169
R3853 IN IN.n6 0.00215441
R3854 IN.n6 IN.n5 0.00197059
R3855 code[3].n0 code[3].t0 229.971
R3856 code[3].n0 code[3].t1 158.35
R3857 code[3].n1 code[3].n0 8.50845
R3858 code[3].n1 code[3] 3.95275
R3859 code[3].n2 code[3].n1 1.73287
R3860 code[3].n3 code[3] 0.474765
R3861 code[3] code[3].n3 0.366977
R3862 code[3].n2 code[3] 0.339042
R3863 code[3].n3 code[3].n2 0.00334091
R3864 code[0] code[0].t0 140.376
C0 a_9893_327# a_9805_327# 0.0022f
C1 VDD x2.floating 0.0334f
C2 x5[7].floating a_9830_2130# 2.76e-19
C3 code[2] x3[1].floating 0.00115f
C4 x6.SW a_9805_327# 3.1e-20
C5 x6.floating code_offset 0.0624f
C6 x10.Y x2.floating 0.00202f
C7 a_9805_1155# x6.SW 0.00179f
C8 x7.floating x6.SW 9.72e-19
C9 code[0] x5[7].floating 0.00119f
C10 VDD a_9893_1293# 1.29e-19
C11 IN a_9805_603# 0.0136f
C12 IN code[3] 0.00346f
C13 code[1] x4[3].floating 0.00929f
C14 a_15703_1681# x9.output_stack 0.00887f
C15 a_9965_1017# x6.SW 2.44e-19
C16 a_9830_2682# x6.floating 0.00578f
C17 a_15703_1681# OUT 0.137f
C18 a_9805_879# a_9965_741# 0.0388f
C19 VDD a_9830_2130# 0.103f
C20 code_offset a_9893_879# 4.7e-19
C21 x10.Y a_9830_2130# 0.039f
C22 a_9805_879# x10.Y 6.65e-20
C23 IN x6.floating 0.0299f
C24 code[0] VDD 0.00321f
C25 a_9805_1155# a_9893_1293# 0.00227f
C26 x7.floating a_9893_1293# 8.52e-19
C27 a_9918_2268# a_9830_2130# 0.0704f
C28 x4[3].floating x9.output_stack 0.636f
C29 code[0] x10.Y 0.0124f
C30 code_offset a_9965_465# 3.98e-19
C31 a_9805_879# a_9805_1155# 0.0316f
C32 x5[7].floating code_offset 0.00308f
C33 x7.floating a_9805_879# 0.00409f
C34 x6.floating code[3] 0.00519f
C35 a_9918_2544# code_offset 1.9e-19
C36 IN a_9893_879# 5.05e-19
C37 a_9965_1017# a_9805_879# 0.0388f
C38 a_9830_2682# x5[7].floating 2.14e-19
C39 VDD code_offset 0.2f
C40 code_offset a_9965_741# 8.34e-19
C41 a_9830_2682# a_9918_2544# 0.0704f
C42 IN a_9965_465# 0.0135f
C43 a_15703_1681# a_15703_1340# 0.0158f
C44 IN x5[7].floating 0.00127f
C45 code[1] x9.output_stack 0.0622f
C46 x4[3].floating x3[1].floating 1.19f
C47 code_offset a_9893_741# 3.54e-19
C48 code_offset x10.Y 0.0402f
C49 code[1] OUT 5.47e-22
C50 IN a_9918_2544# 0.00847f
C51 code_offset a_9805_327# 2.98e-19
C52 a_9830_2682# VDD 0.109f
C53 a_9918_2268# code_offset 3.64e-19
C54 a_9965_465# a_9805_603# 0.0388f
C55 a_9830_2682# x10.Y 1.02e-19
C56 code_offset a_9805_1155# 0.0165f
C57 x7.floating code_offset 0.17f
C58 IN VDD 0.323f
C59 IN a_9965_741# 0.0135f
C60 a_9965_1017# code_offset 0.00297f
C61 OUT x9.output_stack 0.127f
C62 IN a_9893_741# 3.4e-19
C63 IN x10.Y 0.0967f
C64 x6.floating a_9965_465# 0.00109f
C65 code[2] code_offset 0.00739f
C66 x6.floating x5[7].floating 1.18f
C67 code[1] x3[1].floating 0.219f
C68 IN a_9805_327# 0.0127f
C69 a_9965_741# a_9805_603# 0.0388f
C70 VDD code[3] 0.126f
C71 IN a_9918_2268# 0.00921f
C72 x6.floating a_9918_2544# 0.0191f
C73 code_offset a_9893_603# 2.7e-19
C74 IN a_9805_1155# 0.0217f
C75 a_9805_603# a_9893_741# 0.00227f
C76 x10.Y a_9805_603# 4.07e-20
C77 IN x7.floating 0.0241f
C78 x10.Y code[3] 0.0519f
C79 code_offset a_9893_465# 2.1e-19
C80 a_9805_327# a_9805_603# 0.0316f
C81 code[1] a_15703_1340# 3.4e-20
C82 IN a_9965_1017# 0.0135f
C83 x6.floating VDD 5.72f
C84 x6.floating a_9965_741# 0.00167f
C85 x3[1].floating x9.output_stack 0.341f
C86 x7.floating a_9805_603# 0.00409f
C87 x4[3].floating a_9805_879# 1.17e-19
C88 a_9805_879# a_9893_1017# 0.00227f
C89 x6.floating x10.Y 0.0881f
C90 IN a_9893_603# 2.42e-19
C91 code[1] x2.floating 0.0027f
C92 x6.floating a_9918_2268# 0.0194f
C93 code[0] x4[3].floating 2.28e-21
C94 IN a_9893_465# 1.8e-19
C95 a_9893_879# a_9965_741# 0.00227f
C96 x6.floating x7.floating 0.202f
C97 a_15703_1340# x9.output_stack 0.00892f
C98 x5[7].floating a_9918_2544# 0.00154f
C99 OUT a_15703_1340# 0.141f
C100 x6.SW x9.output_stack 0.164f
C101 a_9805_603# a_9893_603# 0.00227f
C102 x6.floating a_9965_1017# 0.00278f
C103 a_9965_741# a_9965_465# 0.0316f
C104 x5[7].floating VDD 43.9f
C105 x2.floating x9.output_stack 0.193f
C106 OUT x2.floating 0.0191f
C107 x7.floating a_9893_879# 8.52e-19
C108 x5[7].floating x10.Y 1.01f
C109 a_9918_2544# VDD 0.128f
C110 x4[3].floating code_offset 0.00402f
C111 code[1] code[0] 0.0619f
C112 code_offset a_9893_1017# 6.22e-19
C113 a_9965_465# a_9805_327# 0.0388f
C114 a_9893_1293# x9.output_stack 0.00227f
C115 a_9918_2544# x10.Y 1.49e-19
C116 x5[7].floating a_9918_2268# 0.00169f
C117 x3[1].floating a_15703_1340# 3.09e-19
C118 x7.floating a_9965_465# 0.00925f
C119 x5[7].floating x7.floating 0.182f
C120 a_9830_2130# x9.output_stack 0.0702f
C121 a_9918_2544# a_9918_2268# 0.0316f
C122 a_9965_741# a_9893_741# 0.00227f
C123 VDD x10.Y 2.7f
C124 x3[1].floating x2.floating 1.17f
C125 a_9830_2406# x6.SW 9.98e-20
C126 code[0] x9.output_stack 0.0232f
C127 x5[7].floating code[2] 0.0056f
C128 IN x4[3].floating 6.65e-19
C129 a_9918_2268# VDD 0.0732f
C130 IN a_9893_1017# 7.93e-19
C131 code[0] OUT 8.53e-20
C132 x10.Y a_9805_327# 2.2e-20
C133 a_9965_465# a_9893_603# 0.00227f
C134 VDD a_9805_1155# 0.00115f
C135 x7.floating a_9965_741# 0.00959f
C136 x7.floating VDD 0.0282f
C137 a_9918_2268# x10.Y 4.2e-19
C138 a_9965_465# a_9893_465# 0.00227f
C139 x10.Y a_9805_1155# 1.69e-19
C140 x4[3].floating a_9805_603# 1.17e-19
C141 x7.floating a_9893_741# 8.52e-19
C142 x7.floating x10.Y 0.00345f
C143 x2.floating a_15703_1340# 0.0104f
C144 a_9965_1017# a_9965_741# 0.0316f
C145 code[2] VDD 0.0372f
C146 x7.floating a_9805_327# 0.00218f
C147 code[2] x10.Y 0.00201f
C148 x7.floating a_9805_1155# 0.00409f
C149 code_offset x9.output_stack 0.255f
C150 code[0] x3[1].floating 0.0326f
C151 a_9830_2406# a_9830_2130# 0.0316f
C152 a_9965_1017# a_9805_1155# 0.0388f
C153 x7.floating a_9965_1017# 0.00959f
C154 a_9830_2130# x6.SW 0.00707f
C155 a_9805_879# x6.SW 8.11e-20
C156 x7.floating code[2] 0.0056f
C157 a_9893_1155# code_offset 7.9e-19
C158 a_15703_1681# x5[7].floating 0.0132f
C159 code[0] a_15703_1340# 0.00169f
C160 a_9805_327# a_9893_465# 0.00227f
C161 x7.floating a_9893_603# 8.52e-19
C162 IN x9.output_stack 0.37f
C163 x7.floating a_9893_465# 8.52e-19
C164 code[0] x2.floating 0.161f
C165 x4[3].floating a_9965_465# 7.47e-19
C166 x5[7].floating x4[3].floating 1.55f
C167 IN a_9893_1155# 0.0013f
C168 a_15703_1681# VDD 0.211f
C169 a_9830_2406# code_offset 6.38e-19
C170 a_15703_1681# x10.Y 0.00127f
C171 code_offset a_9893_327# 1.6e-19
C172 code_offset x6.SW 0.19f
C173 x6.floating x9.output_stack 0.229f
C174 a_9830_2682# a_9830_2406# 0.0316f
C175 x4[3].floating VDD 0.0565f
C176 x4[3].floating a_9965_741# 8.29e-19
C177 x4[3].floating x10.Y 0.00668f
C178 a_9830_2682# x6.SW 5.11e-20
C179 IN a_9830_2406# 0.00866f
C180 code[1] x5[7].floating 0.0022f
C181 x4[3].floating a_9805_327# 7.17e-20
C182 IN a_9893_327# 1.34e-19
C183 code_offset a_9893_1293# 9.08e-19
C184 IN x6.SW 0.0928f
C185 x4[3].floating a_9805_1155# 1.17e-19
C186 x7.floating x4[3].floating 1.18f
C187 x7.floating a_9893_1017# 8.52e-19
C188 code_offset a_9830_2130# 0.00273f
C189 a_9805_879# code_offset 0.0014f
C190 x4[3].floating a_9965_1017# 8.29e-19
C191 code[1] VDD 0.0181f
C192 a_9965_1017# a_9893_1017# 0.00227f
C193 x9.output_stack a_9965_465# 8.05e-20
C194 x5[7].floating x9.output_stack 1.19f
C195 x6.SW a_9805_603# 4.74e-20
C196 code[3] x6.SW 0.00466f
C197 x4[3].floating code[2] 0.518f
C198 x5[7].floating OUT 0.0199f
C199 code[1] x10.Y 6.64e-19
C200 x6.floating a_9830_2406# 0.00996f
C201 a_9918_2544# x9.output_stack 1.5e-19
C202 IN a_9893_1293# 0.00196f
C203 x6.floating x6.SW 0.13f
C204 IN a_9830_2130# 0.0175f
C205 IN a_9805_879# 0.0136f
C206 VDD x9.output_stack 0.594f
C207 a_9965_741# x9.output_stack 1.74e-19
C208 OUT VDD 0.239f
C209 x10.Y x9.output_stack 1.01f
C210 OUT x10.Y 1.13e-19
C211 x5[7].floating x3[1].floating 0.8f
C212 code[1] code[2] 0.00401f
C213 a_9830_2130# code[3] 2.69e-19
C214 a_9805_879# a_9805_603# 0.0316f
C215 a_9918_2268# x9.output_stack 0.032f
C216 a_9805_1155# x9.output_stack 0.0388f
C217 x7.floating x9.output_stack 0.185f
C218 x5[7].floating a_9830_2406# 2.76e-19
C219 a_9830_2682# code_offset 3.28e-19
C220 x6.floating a_9830_2130# 0.00996f
C221 a_9965_1017# x9.output_stack 0.032f
C222 a_9918_2544# a_9830_2406# 0.0704f
C223 x6.SW a_9965_465# 7.9e-20
C224 VDD x3[1].floating 0.0301f
C225 x5[7].floating x6.SW 0.00138f
C226 code[2] x9.output_stack 0.322f
C227 a_9893_1155# a_9805_1155# 0.00227f
C228 x7.floating a_9893_1155# 8.52e-19
C229 x10.Y x3[1].floating 0.00302f
C230 IN code_offset 0.239f
C231 a_9830_2406# VDD 0.0313f
C232 x5[7].floating x2.floating 0.441f
C233 a_9893_1155# a_9965_1017# 0.00227f
C234 VDD a_15703_1340# 0.235f
C235 a_9805_879# a_9893_879# 0.00227f
C236 a_9830_2406# x10.Y 2.35e-19
C237 IN a_9830_2682# 0.00832f
C238 VDD x6.SW 0.423f
C239 a_9965_741# x6.SW 1.28e-19
C240 code_offset a_9805_603# 5.57e-19
C241 code_offset code[3] 0.0293f
C242 a_9830_2406# a_9918_2268# 0.0704f
C243 x10.Y x6.SW 0.788f
C244 OUT VSS 0.422f
C245 a_9893_327# VSS 0.00426f
C246 a_9893_465# VSS 9.21e-19
C247 a_9805_327# VSS 0.177f
C248 a_9965_465# VSS 0.164f
C249 a_9893_603# VSS 8.65e-19
C250 a_9893_741# VSS 8.09e-19
C251 a_9805_603# VSS 0.114f
C252 a_9965_741# VSS 0.114f
C253 a_9893_879# VSS 7.57e-19
C254 a_9893_1017# VSS 7.1e-19
C255 a_9805_879# VSS 0.114f
C256 a_9965_1017# VSS 0.111f
C257 a_9893_1155# VSS 6.69e-19
C258 a_9893_1293# VSS 6.32e-19
C259 a_9805_1155# VSS 0.119f
C260 a_15703_1340# VSS 0.293f
C261 x2.floating VSS 6.42f
C262 x3[1].floating VSS 10.9f
C263 x4[3].floating VSS 21.7f
C264 x7.floating VSS 5.91f
C265 code[0] VSS 0.761f
C266 code[1] VSS 0.911f
C267 code[2] VSS 1.61f
C268 x5[7].floating VSS 0.107p
C269 x6.floating VSS 0.412f
C270 a_15703_1681# VSS 0.32f
C271 x9.output_stack VSS 1.56f
C272 x6.SW VSS 0.299f
C273 x10.Y VSS 2.76f
C274 code_offset VSS 1.11f
C275 code[3] VSS 0.267f
C276 a_9830_2130# VSS 0.0147f
C277 a_9918_2268# VSS 0.0402f
C278 a_9830_2406# VSS 0.0815f
C279 a_9918_2544# VSS 0.032f
C280 a_9830_2682# VSS 0.0953f
C281 IN VSS 1.42f
C282 VDD VSS 37.6f
C283 VDD.n0 VSS 0.0243f
C284 VDD.t13 VSS 0.0585f
C285 VDD.n1 VSS 0.0114f
C286 VDD.n2 VSS 0.0143f
C287 VDD.n3 VSS 0.105f
C288 VDD.n4 VSS 0.016f
C289 VDD.n5 VSS 0.00294f
C290 VDD.n6 VSS 0.00448f
C291 VDD.n7 VSS 0.0245f
C292 VDD.n8 VSS 0.01f
C293 VDD.n9 VSS 0.00508f
C294 VDD.n10 VSS 0.00772f
C295 VDD.n11 VSS 0.00792f
C296 VDD.n12 VSS 0.0127f
C297 VDD.n13 VSS 0.00792f
C298 VDD.n14 VSS 9.36e-19
C299 VDD.n15 VSS 0.0214f
C300 VDD.n16 VSS 0.0196f
C301 VDD.n17 VSS 0.0266f
C302 VDD.n18 VSS 0.047f
C303 VDD.n19 VSS 0.0227f
C304 VDD.n20 VSS 0.0183f
C305 VDD.n21 VSS 0.0142f
C306 VDD.n22 VSS 0.00345f
C307 VDD.n23 VSS 0.0695f
C308 VDD.n24 VSS 0.0142f
C309 VDD.n25 VSS 0.0315f
C310 VDD.n26 VSS 0.00468f
C311 VDD.n27 VSS 0.0211f
C312 VDD.t10 VSS 0.0585f
C313 VDD.n28 VSS 0.0644f
C314 VDD.t16 VSS 2.68f
C315 VDD.n29 VSS 0.00954f
C316 VDD.n30 VSS 0.0229f
C317 VDD.n31 VSS 0.0228f
C318 VDD.n32 VSS 0.0526f
C319 VDD.n33 VSS 0.0221f
C320 VDD.n34 VSS 0.0197f
C321 VDD.n35 VSS 0.00902f
C322 VDD.n36 VSS 0.0193f
C323 VDD.n37 VSS 0.00761f
C324 VDD.t15 VSS 0.00762f
C325 VDD.t3 VSS 0.00762f
C326 VDD.n38 VSS 0.0187f
C327 VDD.n39 VSS 0.0554f
C328 VDD.n40 VSS 0.00925f
C329 VDD.n41 VSS 0.0189f
C330 VDD.n42 VSS 0.115f
C331 VDD.n43 VSS 0.129f
C332 VDD.n44 VSS 0.0228f
C333 VDD.t1 VSS 0.0108f
C334 VDD.n45 VSS 0.157f
C335 VDD.n46 VSS 0.023f
C336 VDD.n47 VSS 0.0125f
C337 VDD.n48 VSS 0.185f
C338 VDD.n49 VSS 0.185f
C339 VDD.n50 VSS 0.0524f
C340 VDD.n51 VSS 0.0228f
C341 VDD.n52 VSS 0.00728f
C342 VDD.n53 VSS 0.0229f
C343 VDD.n54 VSS 0.0524f
C344 VDD.n55 VSS 0.0228f
C345 VDD.n56 VSS 0.00728f
C346 VDD.n57 VSS 0.0229f
C347 VDD.n58 VSS 0.0524f
C348 VDD.n59 VSS 0.0228f
C349 VDD.n60 VSS 0.00728f
C350 VDD.n61 VSS 0.0229f
C351 VDD.n62 VSS 0.0524f
C352 VDD.n63 VSS 0.0228f
C353 VDD.n64 VSS 0.00728f
C354 VDD.n65 VSS 0.0229f
C355 VDD.n66 VSS 0.00643f
C356 VDD.n67 VSS 0.00505f
C357 VDD.n68 VSS 0.00381f
C358 VDD.n69 VSS 5.44e-19
C359 VDD.n70 VSS 0.00308f
C360 VDD.n71 VSS 0.00308f
C361 VDD.n72 VSS 0.0148f
C362 VDD.n75 VSS 0.012f
C363 VDD.n78 VSS 0.0269f
C364 VDD.n82 VSS 0.012f
C365 VDD.n84 VSS 0.012f
C366 VDD.n87 VSS 0.0269f
C367 VDD.n91 VSS 0.012f
C368 VDD.n93 VSS 0.012f
C369 VDD.n96 VSS 0.0269f
C370 VDD.n100 VSS 0.012f
C371 VDD.n102 VSS 0.012f
C372 VDD.n105 VSS 0.0269f
C373 VDD.n108 VSS 0.529f
C374 VDD.n109 VSS 0.0232f
C375 VDD.n114 VSS 0.0269f
C376 VDD.n116 VSS 0.012f
C377 VDD.n118 VSS 0.012f
C378 VDD.n119 VSS 0.0199f
C379 VDD.n120 VSS 0.0199f
C380 VDD.n125 VSS 0.0269f
C381 VDD.n127 VSS 0.012f
C382 VDD.n129 VSS 0.012f
C383 VDD.n130 VSS 0.0199f
C384 VDD.n131 VSS 0.0199f
C385 VDD.n136 VSS 0.0269f
C386 VDD.n138 VSS 0.012f
C387 VDD.n140 VSS 0.012f
C388 VDD.n141 VSS 0.0199f
C389 VDD.n142 VSS 0.0199f
C390 VDD.n147 VSS 0.0269f
C391 VDD.n149 VSS 0.00318f
C392 VDD.n150 VSS 0.0148f
C393 VDD.n151 VSS 0.00308f
C394 VDD.n152 VSS 0.00308f
C395 VDD.n153 VSS 0.0105f
C396 VDD.n154 VSS 5.44e-19
C397 VDD.n155 VSS 0.00381f
C398 VDD.n156 VSS 0.00671f
C399 VDD.n157 VSS 0.00399f
C400 VDD.n158 VSS 5.44e-19
C401 VDD.n159 VSS 0.00542f
C402 VDD.n160 VSS 3.74e-19
C403 VDD.n161 VSS 0.0107f
C404 VDD.n162 VSS -0.0864f
C405 VDD.n163 VSS 0.0107f
C406 VDD.n164 VSS 0.00916f
C407 VDD.n165 VSS 0.00399f
C408 VDD.n166 VSS 0.00308f
C409 VDD.n167 VSS 0.00308f
C410 VDD.n168 VSS 0.00318f
C411 VDD.n169 VSS 0.00308f
C412 VDD.n170 VSS 0.0105f
C413 VDD.n171 VSS 0.00381f
C414 VDD.n172 VSS 0.00505f
C415 VDD.n173 VSS -0.216f
C416 VDD.n174 VSS -0.107f
C417 VDD.n175 VSS 3.74e-19
C418 VDD.n176 VSS 0.00561f
C419 VDD.n177 VSS 0.00916f
C420 VDD.n178 VSS 0.00399f
C421 VDD.n179 VSS 0.0112f
C422 VDD.n180 VSS 0.0112f
C423 VDD.n181 VSS 0.00381f
C424 VDD.n182 VSS 0.00762f
C425 VDD.n183 VSS 0.00925f
C426 VDD.n184 VSS 0.00472f
C427 VDD.n185 VSS 0.00671f
C428 VDD.n186 VSS 0.00542f
C429 VDD.n187 VSS 0.0043f
C430 VDD.n188 VSS 0.0105f
C431 VDD.n189 VSS 0.00643f
C432 VDD.n190 VSS 0.00664f
C433 VDD.n191 VSS 3.74e-19
C434 VDD.n192 VSS 0.00561f
C435 VDD.n193 VSS 5.44e-19
C436 VDD.n194 VSS 0.00399f
C437 VDD.n195 VSS 3.63e-19
C438 VDD.n196 VSS 0.012f
C439 VDD.n197 VSS 0.0148f
C440 VDD.n198 VSS 0.0112f
C441 VDD.n199 VSS 0.0112f
C442 VDD.n200 VSS 0.00381f
C443 VDD.n201 VSS 0.00762f
C444 VDD.n202 VSS 0.00925f
C445 VDD.n203 VSS 0.00381f
C446 VDD.n204 VSS 0.00472f
C447 VDD.n205 VSS 0.00671f
C448 VDD.n206 VSS -0.243f
C449 VDD.n207 VSS 0.0043f
C450 VDD.n208 VSS 0.0105f
C451 VDD.n209 VSS 0.00643f
C452 VDD.n210 VSS 0.00664f
C453 VDD.n211 VSS 3.74e-19
C454 VDD.n212 VSS 0.00561f
C455 VDD.n213 VSS 0.00916f
C456 VDD.n214 VSS 0.0043f
C457 VDD.n215 VSS 0.0105f
C458 VDD.n216 VSS 0.0105f
C459 VDD.n217 VSS 0.00561f
C460 VDD.n218 VSS 0.00505f
C461 VDD.n219 VSS 0.00925f
C462 VDD.n220 VSS 0.00381f
C463 VDD.n221 VSS 0.00762f
C464 VDD.n222 VSS 5.44e-19
C465 VDD.n223 VSS 0.00308f
C466 VDD.n224 VSS 0.0112f
C467 VDD.n225 VSS 0.0112f
C468 VDD.n226 VSS 0.00318f
C469 VDD.n227 VSS 0.00308f
C470 VDD.n228 VSS 3.63e-19
C471 VDD.n229 VSS 0.00308f
C472 VDD.n230 VSS 0.00399f
C473 VDD.n231 VSS 0.00308f
C474 VDD.n232 VSS 0.00381f
C475 VDD.n233 VSS 0.0112f
C476 VDD.n234 VSS 0.0148f
C477 VDD.n235 VSS 0.0112f
C478 VDD.n236 VSS 0.00308f
C479 VDD.n237 VSS 0.0112f
C480 VDD.n238 VSS 0.0105f
C481 VDD.n239 VSS 0.00399f
C482 VDD.n240 VSS 0.00472f
C483 VDD.n241 VSS 0.0043f
C484 VDD.n242 VSS 3.74e-19
C485 VDD.n243 VSS 0.00643f
C486 VDD.n244 VSS 0.00664f
C487 VDD.n245 VSS 3.74e-19
C488 VDD.n246 VSS 0.00561f
C489 VDD.n247 VSS 0.00916f
C490 VDD.n248 VSS 0.0107f
C491 VDD.n249 VSS 0.0105f
C492 VDD.n250 VSS 0.00643f
C493 VDD.n251 VSS 0.00399f
C494 VDD.n252 VSS 0.00561f
C495 VDD.n253 VSS 0.00308f
C496 VDD.n254 VSS 0.0148f
C497 VDD.n255 VSS 0.00318f
C498 VDD.n256 VSS 0.00308f
C499 VDD.n257 VSS 0.0337f
C500 VDD.n258 VSS 0.0299f
C501 VDD.n259 VSS 5.44e-19
C502 VDD.n260 VSS 0.00381f
C503 VDD.n261 VSS 0.00399f
C504 VDD.n262 VSS 0.00308f
C505 VDD.n263 VSS 0.00762f
C506 VDD.n264 VSS 0.00399f
C507 VDD.n265 VSS 0.00925f
C508 VDD.n266 VSS 0.00381f
C509 VDD.n267 VSS 0.00897f
C510 VDD.n268 VSS 0.00505f
C511 VDD.n269 VSS 0.00664f
C512 VDD.n270 VSS 0.00542f
C513 VDD.n271 VSS 0.00664f
C514 VDD.n272 VSS 0.0379f
C515 VDD.n273 VSS 0.0329f
C516 VDD.n274 VSS 0.0327f
C517 VDD.n275 VSS 0.0377f
C518 VDD.n276 VSS 0.00643f
C519 VDD.n277 VSS 3.74e-19
C520 VDD.n278 VSS -0.0864f
C521 VDD.n279 VSS 0.00381f
C522 VDD.n280 VSS 0.0105f
C523 VDD.n281 VSS 0.00472f
C524 VDD.n282 VSS 0.00671f
C525 VDD.n283 VSS -0.243f
C526 VDD.n284 VSS 0.00448f
C527 VDD.n285 VSS 0.0107f
C528 VDD.n286 VSS 0.0105f
C529 VDD.n287 VSS -0.224f
C530 VDD.n288 VSS 0.00561f
C531 VDD.n289 VSS 3.74e-19
C532 VDD.n290 VSS 0.00399f
C533 VDD.n291 VSS 0.00381f
C534 VDD.n292 VSS 0.00308f
C535 VDD.n293 VSS 0.0105f
C536 VDD.n294 VSS 0.00308f
C537 VDD.n295 VSS 0.00308f
C538 VDD.n296 VSS 0.00762f
C539 VDD.n297 VSS 0.00399f
C540 VDD.n298 VSS 0.00925f
C541 VDD.n299 VSS 0.00381f
C542 VDD.n300 VSS 0.00897f
C543 VDD.n301 VSS -0.0864f
C544 VDD.n302 VSS -0.099f
C545 VDD.n303 VSS 0.00664f
C546 VDD.n304 VSS 0.00505f
C547 VDD.n305 VSS 0.00472f
C548 VDD.n306 VSS 0.00671f
C549 VDD.n307 VSS 0.00561f
C550 VDD.n308 VSS 0.00448f
C551 VDD.n309 VSS 0.0107f
C552 VDD.n310 VSS 0.0105f
C553 VDD.n311 VSS 0.0105f
C554 VDD.n312 VSS -0.243f
C555 VDD.n313 VSS 3.74e-19
C556 VDD.n314 VSS 0.00399f
C557 VDD.n315 VSS 0.00381f
C558 VDD.n316 VSS 0.00308f
C559 VDD.n317 VSS 0.0105f
C560 VDD.n318 VSS 0.00308f
C561 VDD.n319 VSS 0.00308f
C562 VDD.n320 VSS 0.00762f
C563 VDD.n321 VSS 0.00399f
C564 VDD.n322 VSS 0.00925f
C565 VDD.n323 VSS 0.00381f
C566 VDD.n324 VSS 0.00897f
C567 VDD.n325 VSS 0.00505f
C568 VDD.n326 VSS 0.00643f
C569 VDD.n327 VSS 0.00664f
C570 VDD.n328 VSS 0.00505f
C571 VDD.n329 VSS 0.00472f
C572 VDD.n330 VSS 0.00671f
C573 VDD.n331 VSS 0.00561f
C574 VDD.n332 VSS 0.00448f
C575 VDD.n333 VSS 0.0107f
C576 VDD.n334 VSS -0.224f
C577 VDD.n335 VSS 0.00561f
C578 VDD.n336 VSS 0.00542f
C579 VDD.n337 VSS -0.107f
C580 VDD.n338 VSS 3.74e-19
C581 VDD.n339 VSS 0.00472f
C582 VDD.n340 VSS 0.00399f
C583 VDD.n341 VSS 0.00561f
C584 VDD.n342 VSS 0.0288f
C585 VDD.n343 VSS 0.0288f
C586 VDD.n344 VSS 0.00472f
C587 VDD.n345 VSS 0.0339f
C588 VDD.n346 VSS 0.0339f
C589 VDD.n347 VSS 0.00308f
C590 VDD.n348 VSS 3.63e-19
C591 VDD.n349 VSS 0.012f
C592 VDD.n350 VSS 0.00318f
C593 VDD.n351 VSS 0.00308f
C594 VDD.n352 VSS 0.0359f
C595 VDD.n353 VSS 0.0359f
C596 VDD.n354 VSS 0.00318f
C597 VDD.n355 VSS 0.00308f
C598 VDD.n356 VSS 0.0148f
C599 VDD.n357 VSS 0.0112f
C600 VDD.n358 VSS 0.0105f
C601 VDD.n359 VSS 0.00472f
C602 VDD.n360 VSS 0.0043f
C603 VDD.n361 VSS 3.74e-19
C604 VDD.n362 VSS 0.00916f
C605 VDD.n363 VSS -0.216f
C606 VDD.n364 VSS 0.0105f
C607 VDD.n365 VSS 0.00643f
C608 VDD.n366 VSS 0.00399f
C609 VDD.n367 VSS 0.00561f
C610 VDD.n368 VSS 0.00308f
C611 VDD.n369 VSS 0.00318f
C612 VDD.n370 VSS 0.00308f
C613 VDD.n371 VSS 0.0148f
C614 VDD.n372 VSS 0.0112f
C615 VDD.n373 VSS 0.0105f
C616 VDD.n374 VSS 0.00472f
C617 VDD.n375 VSS 0.0043f
C618 VDD.n376 VSS 3.74e-19
C619 VDD.n377 VSS 0.00664f
C620 VDD.n378 VSS 0.00916f
C621 VDD.n379 VSS 0.0107f
C622 VDD.n380 VSS 0.0105f
C623 VDD.n381 VSS 0.00643f
C624 VDD.n382 VSS 0.00399f
C625 VDD.n383 VSS 0.00561f
C626 VDD.n384 VSS 0.00308f
C627 VDD.n385 VSS 0.00318f
C628 VDD.n386 VSS 0.00308f
C629 VDD.n387 VSS 0.0148f
C630 VDD.n388 VSS 0.0112f
C631 VDD.n389 VSS 0.0105f
C632 VDD.n390 VSS 0.00472f
C633 VDD.n391 VSS 0.0043f
C634 VDD.n392 VSS 3.74e-19
C635 VDD.n393 VSS 0.00664f
C636 VDD.n394 VSS 0.00916f
C637 VDD.n395 VSS 0.0107f
C638 VDD.n396 VSS 0.0105f
C639 VDD.n397 VSS 0.00643f
C640 VDD.n398 VSS 0.00399f
C641 VDD.n399 VSS 0.00561f
C642 VDD.n400 VSS 0.00308f
C643 VDD.n401 VSS 0.00318f
C644 VDD.n402 VSS 0.00308f
C645 VDD.n403 VSS 0.0148f
C646 VDD.n404 VSS 0.0112f
C647 VDD.n405 VSS 0.0105f
C648 VDD.n406 VSS 0.00472f
C649 VDD.n407 VSS 0.0043f
C650 VDD.n408 VSS 3.74e-19
C651 VDD.n409 VSS -0.107f
C652 VDD.n410 VSS 0.00916f
C653 VDD.n411 VSS -0.216f
C654 VDD.n412 VSS 0.0105f
C655 VDD.n413 VSS 0.00643f
C656 VDD.n414 VSS 0.00399f
C657 VDD.n415 VSS 0.00561f
C658 VDD.n416 VSS 0.00308f
C659 VDD.n417 VSS 0.00308f
C660 VDD.n418 VSS 0.0112f
C661 VDD.n419 VSS 0.0105f
C662 VDD.n420 VSS 0.00472f
C663 VDD.n421 VSS 0.0043f
C664 VDD.n422 VSS 3.74e-19
C665 VDD.n423 VSS 0.00664f
C666 VDD.n424 VSS 0.00916f
C667 VDD.n425 VSS 0.0107f
C668 VDD.n426 VSS 0.0105f
C669 VDD.n427 VSS 0.00643f
C670 VDD.n428 VSS 0.00399f
C671 VDD.n429 VSS 0.00561f
C672 VDD.n430 VSS 0.00308f
C673 VDD.n431 VSS 0.0148f
C674 VDD.n432 VSS 0.00318f
C675 VDD.n433 VSS 0.00308f
C676 VDD.n434 VSS 0.0337f
C677 VDD.n435 VSS 0.0299f
C678 VDD.n436 VSS 5.44e-19
C679 VDD.n437 VSS 0.00381f
C680 VDD.n438 VSS 0.00399f
C681 VDD.n439 VSS 0.00308f
C682 VDD.n440 VSS 0.00762f
C683 VDD.n441 VSS 0.00399f
C684 VDD.n442 VSS 0.00925f
C685 VDD.n443 VSS 0.00381f
C686 VDD.n444 VSS 0.00897f
C687 VDD.n445 VSS 0.00505f
C688 VDD.n446 VSS 0.00664f
C689 VDD.n447 VSS 0.00542f
C690 VDD.n448 VSS 0.00664f
C691 VDD.n449 VSS 0.0379f
C692 VDD.n450 VSS 0.0329f
C693 VDD.n451 VSS 0.0327f
C694 VDD.n452 VSS 0.0377f
C695 VDD.n453 VSS 0.00643f
C696 VDD.n454 VSS 3.74e-19
C697 VDD.n455 VSS -0.0864f
C698 VDD.n456 VSS 0.00381f
C699 VDD.n457 VSS 0.0105f
C700 VDD.n458 VSS 0.00472f
C701 VDD.n459 VSS 0.00671f
C702 VDD.n460 VSS -0.243f
C703 VDD.n461 VSS 0.00448f
C704 VDD.n462 VSS 0.0107f
C705 VDD.n463 VSS 0.0105f
C706 VDD.n464 VSS -0.224f
C707 VDD.n465 VSS 0.00561f
C708 VDD.n466 VSS 3.74e-19
C709 VDD.n467 VSS 0.00399f
C710 VDD.n468 VSS 0.00381f
C711 VDD.n469 VSS 0.00308f
C712 VDD.n470 VSS 0.0105f
C713 VDD.n471 VSS 0.00308f
C714 VDD.n472 VSS 0.00308f
C715 VDD.n473 VSS 0.00762f
C716 VDD.n474 VSS 0.00399f
C717 VDD.n475 VSS 0.00925f
C718 VDD.n476 VSS 0.00381f
C719 VDD.n477 VSS 0.00897f
C720 VDD.n478 VSS -0.0864f
C721 VDD.n479 VSS -0.099f
C722 VDD.n480 VSS 0.00664f
C723 VDD.n481 VSS 0.00505f
C724 VDD.n482 VSS 0.00472f
C725 VDD.n483 VSS 0.00671f
C726 VDD.n484 VSS 0.00561f
C727 VDD.n485 VSS 0.00448f
C728 VDD.n486 VSS 0.0107f
C729 VDD.n487 VSS 0.0105f
C730 VDD.n488 VSS 0.0105f
C731 VDD.n489 VSS -0.243f
C732 VDD.n490 VSS 3.74e-19
C733 VDD.n491 VSS 0.00399f
C734 VDD.n492 VSS 0.00381f
C735 VDD.n493 VSS 0.00308f
C736 VDD.n494 VSS 0.0105f
C737 VDD.n495 VSS 0.00308f
C738 VDD.n496 VSS 0.00308f
C739 VDD.n497 VSS 0.00762f
C740 VDD.n498 VSS 0.00399f
C741 VDD.n499 VSS 0.00925f
C742 VDD.n500 VSS 0.00381f
C743 VDD.n501 VSS 0.00897f
C744 VDD.n502 VSS 0.00505f
C745 VDD.n503 VSS 0.00643f
C746 VDD.n504 VSS 0.00664f
C747 VDD.n505 VSS 0.00505f
C748 VDD.n506 VSS 0.00472f
C749 VDD.n507 VSS 0.00671f
C750 VDD.n508 VSS 0.00561f
C751 VDD.n509 VSS 0.00448f
C752 VDD.n510 VSS 0.0107f
C753 VDD.n511 VSS -0.224f
C754 VDD.n512 VSS 0.00561f
C755 VDD.n513 VSS 0.00542f
C756 VDD.n514 VSS -0.107f
C757 VDD.n515 VSS 3.74e-19
C758 VDD.n516 VSS 0.00472f
C759 VDD.n517 VSS 0.00399f
C760 VDD.n518 VSS 0.00561f
C761 VDD.n519 VSS 0.0288f
C762 VDD.n520 VSS 0.0288f
C763 VDD.n521 VSS 0.00472f
C764 VDD.n522 VSS 0.0339f
C765 VDD.n523 VSS 0.0339f
C766 VDD.n524 VSS 0.00308f
C767 VDD.n525 VSS 3.63e-19
C768 VDD.n526 VSS 0.012f
C769 VDD.n527 VSS 0.00318f
C770 VDD.n528 VSS 0.00308f
C771 VDD.n529 VSS 0.0359f
C772 VDD.n530 VSS 0.0359f
C773 VDD.n531 VSS 0.00318f
C774 VDD.n532 VSS 0.00308f
C775 VDD.n533 VSS 0.0148f
C776 VDD.n534 VSS 0.0112f
C777 VDD.n535 VSS 0.0105f
C778 VDD.n536 VSS 0.00472f
C779 VDD.n537 VSS 0.0043f
C780 VDD.n538 VSS 3.74e-19
C781 VDD.n539 VSS 0.00916f
C782 VDD.n540 VSS -0.216f
C783 VDD.n541 VSS 0.0105f
C784 VDD.n542 VSS 0.00643f
C785 VDD.n543 VSS 0.00399f
C786 VDD.n544 VSS 0.00561f
C787 VDD.n545 VSS 0.00308f
C788 VDD.n546 VSS 0.00318f
C789 VDD.n547 VSS 0.00308f
C790 VDD.n548 VSS 0.0148f
C791 VDD.n549 VSS 0.0112f
C792 VDD.n550 VSS 0.0105f
C793 VDD.n551 VSS 0.00472f
C794 VDD.n552 VSS 0.0043f
C795 VDD.n553 VSS 3.74e-19
C796 VDD.n554 VSS 0.00664f
C797 VDD.n555 VSS 0.00916f
C798 VDD.n556 VSS 0.0107f
C799 VDD.n557 VSS 0.0105f
C800 VDD.n558 VSS 0.00643f
C801 VDD.n559 VSS 0.00399f
C802 VDD.n560 VSS 0.00561f
C803 VDD.n561 VSS 0.00308f
C804 VDD.n562 VSS 0.00318f
C805 VDD.n563 VSS 0.00308f
C806 VDD.n564 VSS 0.0148f
C807 VDD.n565 VSS 0.0112f
C808 VDD.n566 VSS 0.0105f
C809 VDD.n567 VSS 0.00472f
C810 VDD.n568 VSS 0.0043f
C811 VDD.n569 VSS 3.74e-19
C812 VDD.n570 VSS 0.00664f
C813 VDD.n571 VSS 0.00916f
C814 VDD.n572 VSS 0.0107f
C815 VDD.n573 VSS 0.0105f
C816 VDD.n574 VSS 0.00643f
C817 VDD.n575 VSS 0.00399f
C818 VDD.n576 VSS 0.00561f
C819 VDD.n577 VSS 0.00308f
C820 VDD.n578 VSS 0.00318f
C821 VDD.n579 VSS 0.00308f
C822 VDD.n580 VSS 0.0148f
C823 VDD.n581 VSS 0.0112f
C824 VDD.n582 VSS 0.0105f
C825 VDD.n583 VSS 0.00472f
C826 VDD.n584 VSS 0.0043f
C827 VDD.n585 VSS 3.74e-19
C828 VDD.n586 VSS -0.107f
C829 VDD.n587 VSS 0.00916f
C830 VDD.n588 VSS -0.216f
C831 VDD.n589 VSS 0.0105f
C832 VDD.n590 VSS 0.00643f
C833 VDD.n591 VSS 0.00399f
C834 VDD.n592 VSS 0.00561f
C835 VDD.n593 VSS 0.00308f
C836 VDD.n594 VSS 0.00308f
C837 VDD.n595 VSS 0.0112f
C838 VDD.n596 VSS 0.0105f
C839 VDD.n597 VSS 0.00472f
C840 VDD.n598 VSS 0.0043f
C841 VDD.n599 VSS 3.74e-19
C842 VDD.n600 VSS 0.00664f
C843 VDD.n601 VSS 0.00916f
C844 VDD.n602 VSS 0.0107f
C845 VDD.n603 VSS 0.0105f
C846 VDD.n604 VSS 0.00643f
C847 VDD.n605 VSS 0.00399f
C848 VDD.n606 VSS 0.00561f
C849 VDD.n607 VSS 0.00308f
C850 VDD.n608 VSS 0.0148f
C851 VDD.n609 VSS 0.00318f
C852 VDD.n610 VSS 0.00308f
C853 VDD.n611 VSS 0.0337f
C854 VDD.n612 VSS 0.0299f
C855 VDD.n613 VSS 5.44e-19
C856 VDD.n614 VSS 0.00381f
C857 VDD.n615 VSS 0.00399f
C858 VDD.n616 VSS 0.00308f
C859 VDD.n617 VSS 0.00762f
C860 VDD.n618 VSS 0.00399f
C861 VDD.n619 VSS 0.00925f
C862 VDD.n620 VSS 0.00381f
C863 VDD.n621 VSS 0.00897f
C864 VDD.n622 VSS 0.00505f
C865 VDD.n623 VSS 0.00664f
C866 VDD.n624 VSS 0.00542f
C867 VDD.n625 VSS 0.00664f
C868 VDD.n626 VSS 0.0379f
C869 VDD.n627 VSS 0.0329f
C870 VDD.n628 VSS 0.0327f
C871 VDD.n629 VSS 0.0377f
C872 VDD.n630 VSS 0.00643f
C873 VDD.n631 VSS 3.74e-19
C874 VDD.n632 VSS -0.0864f
C875 VDD.n633 VSS 0.00381f
C876 VDD.n634 VSS 0.0105f
C877 VDD.n635 VSS 0.00472f
C878 VDD.n636 VSS 0.00671f
C879 VDD.n637 VSS -0.243f
C880 VDD.n638 VSS 0.00448f
C881 VDD.n639 VSS 0.0107f
C882 VDD.n640 VSS 0.0105f
C883 VDD.n641 VSS -0.224f
C884 VDD.n642 VSS 0.00561f
C885 VDD.n643 VSS 3.74e-19
C886 VDD.n644 VSS 0.00399f
C887 VDD.n645 VSS 0.00381f
C888 VDD.n646 VSS 0.00308f
C889 VDD.n647 VSS 0.0105f
C890 VDD.n648 VSS 0.00308f
C891 VDD.n649 VSS 0.00308f
C892 VDD.n650 VSS 0.00762f
C893 VDD.n651 VSS 0.00399f
C894 VDD.n652 VSS 0.00925f
C895 VDD.n653 VSS 0.00381f
C896 VDD.n654 VSS 0.00897f
C897 VDD.n655 VSS -0.0864f
C898 VDD.n656 VSS -0.099f
C899 VDD.n657 VSS 0.00664f
C900 VDD.n658 VSS 0.00505f
C901 VDD.n659 VSS 0.00472f
C902 VDD.n660 VSS 0.00671f
C903 VDD.n661 VSS 0.00561f
C904 VDD.n662 VSS 0.00448f
C905 VDD.n663 VSS 0.0107f
C906 VDD.n664 VSS 0.0105f
C907 VDD.n665 VSS 0.0105f
C908 VDD.n666 VSS -0.243f
C909 VDD.n667 VSS 3.74e-19
C910 VDD.n668 VSS 0.00399f
C911 VDD.n669 VSS 0.00381f
C912 VDD.n670 VSS 0.00308f
C913 VDD.n671 VSS 0.0105f
C914 VDD.n672 VSS 0.00308f
C915 VDD.n673 VSS 0.00308f
C916 VDD.n674 VSS 0.00762f
C917 VDD.n675 VSS 0.00399f
C918 VDD.n676 VSS 0.00925f
C919 VDD.n677 VSS 0.00381f
C920 VDD.n678 VSS 0.00897f
C921 VDD.n679 VSS 0.00505f
C922 VDD.n680 VSS 0.00643f
C923 VDD.n681 VSS 0.00664f
C924 VDD.n682 VSS 0.00505f
C925 VDD.n683 VSS 0.00472f
C926 VDD.n684 VSS 0.00671f
C927 VDD.n685 VSS 0.00561f
C928 VDD.n686 VSS 0.00448f
C929 VDD.n687 VSS 0.0107f
C930 VDD.n688 VSS -0.224f
C931 VDD.n689 VSS 0.00561f
C932 VDD.n690 VSS 0.00542f
C933 VDD.n691 VSS -0.107f
C934 VDD.n692 VSS 3.74e-19
C935 VDD.n693 VSS 0.00472f
C936 VDD.n694 VSS 0.00399f
C937 VDD.n695 VSS 0.00561f
C938 VDD.n696 VSS 0.0288f
C939 VDD.n697 VSS 0.0288f
C940 VDD.n698 VSS 0.00472f
C941 VDD.n699 VSS 0.0339f
C942 VDD.n700 VSS 0.0339f
C943 VDD.n701 VSS 0.00308f
C944 VDD.n702 VSS 3.63e-19
C945 VDD.n703 VSS 0.012f
C946 VDD.n704 VSS 0.00318f
C947 VDD.n705 VSS 0.00308f
C948 VDD.n706 VSS 0.0359f
C949 VDD.n707 VSS 0.0359f
C950 VDD.n708 VSS 0.00318f
C951 VDD.n709 VSS 0.00308f
C952 VDD.n710 VSS 0.0148f
C953 VDD.n711 VSS 0.0112f
C954 VDD.n712 VSS 0.0105f
C955 VDD.n713 VSS 0.00472f
C956 VDD.n714 VSS 0.0043f
C957 VDD.n715 VSS 3.74e-19
C958 VDD.n716 VSS 0.00916f
C959 VDD.n717 VSS -0.216f
C960 VDD.n718 VSS 0.0105f
C961 VDD.n719 VSS 0.00643f
C962 VDD.n720 VSS 0.00399f
C963 VDD.n721 VSS 0.00561f
C964 VDD.n722 VSS 0.00308f
C965 VDD.n723 VSS 0.00318f
C966 VDD.n724 VSS 0.00308f
C967 VDD.n725 VSS 0.0148f
C968 VDD.n726 VSS 0.0112f
C969 VDD.n727 VSS 0.0105f
C970 VDD.n728 VSS 0.00472f
C971 VDD.n729 VSS 0.0043f
C972 VDD.n730 VSS 3.74e-19
C973 VDD.n731 VSS 0.00664f
C974 VDD.n732 VSS 0.00916f
C975 VDD.n733 VSS 0.0107f
C976 VDD.n734 VSS 0.0105f
C977 VDD.n735 VSS 0.00643f
C978 VDD.n736 VSS 0.00399f
C979 VDD.n737 VSS 0.00561f
C980 VDD.n738 VSS 0.00308f
C981 VDD.n739 VSS 0.00318f
C982 VDD.n740 VSS 0.00308f
C983 VDD.n741 VSS 0.0148f
C984 VDD.n742 VSS 0.0112f
C985 VDD.n743 VSS 0.0105f
C986 VDD.n744 VSS 0.00472f
C987 VDD.n745 VSS 0.0043f
C988 VDD.n746 VSS 3.74e-19
C989 VDD.n747 VSS 0.00664f
C990 VDD.n748 VSS 0.00916f
C991 VDD.n749 VSS 0.0107f
C992 VDD.n750 VSS 0.0105f
C993 VDD.n751 VSS 0.00643f
C994 VDD.n752 VSS 0.00399f
C995 VDD.n753 VSS 0.00561f
C996 VDD.n754 VSS 0.00308f
C997 VDD.n755 VSS 0.00318f
C998 VDD.n756 VSS 0.00308f
C999 VDD.n757 VSS 0.0148f
C1000 VDD.n758 VSS 0.0112f
C1001 VDD.n759 VSS 0.0105f
C1002 VDD.n760 VSS 0.00472f
C1003 VDD.n761 VSS 0.0043f
C1004 VDD.n762 VSS 3.74e-19
C1005 VDD.n763 VSS -0.107f
C1006 VDD.n764 VSS 0.00916f
C1007 VDD.n765 VSS -0.216f
C1008 VDD.n766 VSS 0.0105f
C1009 VDD.n767 VSS 0.00643f
C1010 VDD.n768 VSS 0.00399f
C1011 VDD.n769 VSS 0.00561f
C1012 VDD.n770 VSS 0.00308f
C1013 VDD.n771 VSS 0.00308f
C1014 VDD.n772 VSS 0.0112f
C1015 VDD.n773 VSS 0.0105f
C1016 VDD.n774 VSS 0.00472f
C1017 VDD.n775 VSS 0.0043f
C1018 VDD.n776 VSS 3.74e-19
C1019 VDD.n777 VSS 0.00664f
C1020 VDD.n778 VSS 0.00916f
C1021 VDD.n779 VSS 0.0107f
C1022 VDD.n780 VSS 0.0105f
C1023 VDD.n781 VSS 0.00643f
C1024 VDD.n782 VSS 0.00399f
C1025 VDD.n783 VSS 0.00561f
C1026 VDD.n784 VSS 0.00308f
C1027 VDD.n785 VSS 0.0148f
C1028 VDD.n786 VSS 0.00318f
C1029 VDD.n787 VSS 0.00308f
C1030 VDD.n788 VSS 0.0337f
C1031 VDD.n789 VSS 0.0299f
C1032 VDD.n790 VSS 5.44e-19
C1033 VDD.n791 VSS 0.00381f
C1034 VDD.n792 VSS 0.00399f
C1035 VDD.n793 VSS 0.00308f
C1036 VDD.n794 VSS 0.00762f
C1037 VDD.n795 VSS 0.00399f
C1038 VDD.n796 VSS 0.00925f
C1039 VDD.n797 VSS 0.00381f
C1040 VDD.n798 VSS 0.00897f
C1041 VDD.n799 VSS 0.00505f
C1042 VDD.n800 VSS 0.00664f
C1043 VDD.n801 VSS 0.00542f
C1044 VDD.n802 VSS 0.00664f
C1045 VDD.n803 VSS 0.0379f
C1046 VDD.n804 VSS 0.0329f
C1047 VDD.n805 VSS 0.0327f
C1048 VDD.n806 VSS 0.0377f
C1049 VDD.n807 VSS 0.00643f
C1050 VDD.n808 VSS 3.74e-19
C1051 VDD.n809 VSS -0.0864f
C1052 VDD.n810 VSS 0.00381f
C1053 VDD.n811 VSS 0.0105f
C1054 VDD.n812 VSS 0.00472f
C1055 VDD.n813 VSS 0.00671f
C1056 VDD.n814 VSS -0.243f
C1057 VDD.n815 VSS 0.00448f
C1058 VDD.n816 VSS 0.0107f
C1059 VDD.n817 VSS 0.0105f
C1060 VDD.n818 VSS -0.224f
C1061 VDD.n819 VSS 0.00561f
C1062 VDD.n820 VSS 3.74e-19
C1063 VDD.n821 VSS 0.00399f
C1064 VDD.n822 VSS 0.00381f
C1065 VDD.n823 VSS 0.00308f
C1066 VDD.n824 VSS 0.0105f
C1067 VDD.n825 VSS 0.00308f
C1068 VDD.n826 VSS 0.00308f
C1069 VDD.n827 VSS 0.00762f
C1070 VDD.n828 VSS 0.00399f
C1071 VDD.n829 VSS 0.00925f
C1072 VDD.n830 VSS 0.00381f
C1073 VDD.n831 VSS 0.00897f
C1074 VDD.n832 VSS -0.0864f
C1075 VDD.n833 VSS -0.099f
C1076 VDD.n834 VSS 0.00664f
C1077 VDD.n835 VSS 0.00505f
C1078 VDD.n836 VSS 0.00472f
C1079 VDD.n837 VSS 0.00671f
C1080 VDD.n838 VSS 0.00561f
C1081 VDD.n839 VSS 0.00448f
C1082 VDD.n840 VSS 0.0107f
C1083 VDD.n841 VSS 0.0105f
C1084 VDD.n842 VSS 0.0105f
C1085 VDD.n843 VSS -0.243f
C1086 VDD.n844 VSS 3.74e-19
C1087 VDD.n845 VSS 0.00399f
C1088 VDD.n846 VSS 0.00381f
C1089 VDD.n847 VSS 0.00308f
C1090 VDD.n848 VSS 0.0105f
C1091 VDD.n849 VSS 0.00308f
C1092 VDD.n850 VSS 0.00308f
C1093 VDD.n851 VSS 0.00762f
C1094 VDD.n852 VSS 0.0592f
C1095 VDD.n853 VSS 0.0484f
C1096 VDD.n854 VSS 0.00925f
C1097 VDD.n855 VSS 0.00381f
C1098 VDD.n856 VSS 0.00897f
C1099 VDD.n857 VSS 0.00505f
C1100 VDD.n858 VSS 0.00643f
C1101 VDD.n859 VSS 0.00664f
C1102 VDD.n860 VSS 0.00505f
C1103 VDD.n861 VSS 0.00472f
C1104 VDD.n862 VSS 0.00671f
C1105 VDD.n863 VSS 0.00561f
C1106 VDD.n864 VSS 0.00448f
C1107 VDD.n865 VSS 0.0107f
C1108 VDD.n866 VSS -0.224f
C1109 VDD.n867 VSS 0.00667f
C1110 VDD.n868 VSS 3.74e-19
C1111 VDD.n869 VSS 0.0662f
C1112 VDD.n870 VSS 0.00472f
C1113 VDD.n871 VSS -0.243f
C1114 VDD.n872 VSS 0.0109f
C1115 VDD.n873 VSS 3.74e-19
C1116 VDD.n874 VSS 0.00399f
C1117 VDD.n875 VSS 0.00381f
C1118 VDD.n876 VSS 0.00308f
C1119 VDD.n877 VSS 0.0105f
C1120 VDD.n878 VSS 0.00308f
C1121 VDD.n879 VSS 0.00308f
C1122 VDD.n881 VSS 0.036f
C1123 VDD.n882 VSS 0.0271f
C1124 VDD.n883 VSS 0.00318f
C1125 VDD.n884 VSS 0.00308f
C1126 VDD.n885 VSS 0.0109f
C1127 VDD.n886 VSS 0.00671f
C1128 VDD.n887 VSS 0.00925f
C1129 VDD.n888 VSS 0.00762f
C1130 VDD.n889 VSS 0.00381f
C1131 VDD.n890 VSS 0.0112f
C1132 VDD.n891 VSS 0.0112f
C1133 VDD.n892 VSS 0.0148f
C1134 VDD.n893 VSS 0.012f
C1135 VDD.n894 VSS 0.00308f
C1136 VDD.n895 VSS 0.00762f
C1137 VDD.n896 VSS 0.00399f
C1138 VDD.n897 VSS 0.00925f
C1139 VDD.n898 VSS 0.00381f
C1140 VDD.n899 VSS 0.00897f
C1141 VDD.n900 VSS 0.00505f
C1142 VDD.n901 VSS 0.00667f
C1143 VDD.n902 VSS 0.0069f
C1144 VDD.n903 VSS 0.00505f
C1145 VDD.n904 VSS 0.00472f
C1146 VDD.n905 VSS 0.00671f
C1147 VDD.n906 VSS 0.00561f
C1148 VDD.n907 VSS 0.00448f
C1149 VDD.n908 VSS 0.0111f
C1150 VDD.n909 VSS -0.223f
C1151 VDD.n910 VSS 0.0109f
C1152 VDD.n911 VSS 0.00561f
C1153 VDD.n912 VSS 3.74e-19
C1154 VDD.n913 VSS 0.00399f
C1155 VDD.n914 VSS 0.00381f
C1156 VDD.n915 VSS 0.00308f
C1157 VDD.n916 VSS 0.0105f
C1158 VDD.n917 VSS 0.00308f
C1159 VDD.n918 VSS 0.00308f
C1160 VDD.n920 VSS 0.00318f
C1161 VDD.n921 VSS 3.63e-19
C1162 VDD.n922 VSS 0.00308f
C1163 VDD.n923 VSS 0.0105f
C1164 VDD.n924 VSS 0.00472f
C1165 VDD.n925 VSS 0.00671f
C1166 VDD.n926 VSS 0.00925f
C1167 VDD.n927 VSS 0.00762f
C1168 VDD.n928 VSS 0.00381f
C1169 VDD.n929 VSS 0.0112f
C1170 VDD.n930 VSS 0.0112f
C1171 VDD.n931 VSS 0.0148f
C1172 VDD.n932 VSS 0.012f
C1173 VDD.n933 VSS 0.00308f
C1174 VDD.n934 VSS 0.00762f
C1175 VDD.n935 VSS 0.00399f
C1176 VDD.n936 VSS 0.00925f
C1177 VDD.n937 VSS 0.00381f
C1178 VDD.n938 VSS 0.00897f
C1179 VDD.n939 VSS 0.00505f
C1180 VDD.n940 VSS 0.00667f
C1181 VDD.n941 VSS 0.0069f
C1182 VDD.n942 VSS -0.0864f
C1183 VDD.n943 VSS 0.00472f
C1184 VDD.n944 VSS 0.00671f
C1185 VDD.n945 VSS -0.243f
C1186 VDD.n946 VSS 0.00448f
C1187 VDD.n947 VSS 0.0111f
C1188 VDD.n948 VSS 0.0109f
C1189 VDD.n949 VSS -0.223f
C1190 VDD.n950 VSS 0.00561f
C1191 VDD.n951 VSS 3.74e-19
C1192 VDD.n952 VSS 0.00399f
C1193 VDD.n953 VSS 0.00381f
C1194 VDD.n954 VSS 0.00308f
C1195 VDD.n955 VSS 0.0181f
C1196 VDD.n956 VSS 0.00308f
C1197 VDD.n957 VSS 0.00347f
C1198 VDD.t6 VSS 0.0067f
C1199 VDD.n958 VSS 0.014f
C1200 VDD.n959 VSS 0.00851f
C1201 VDD.n960 VSS 0.00709f
C1202 VDD.n961 VSS 0.0305f
C1203 VDD.n962 VSS 0.00472f
C1204 VDD.n963 VSS 0.00895f
C1205 VDD.n964 VSS 0.00561f
C1206 VDD.n965 VSS -0.0987f
C1207 VDD.n966 VSS 0.00505f
C1208 VDD.n967 VSS 0.0069f
C1209 VDD.n968 VSS 0.00734f
C1210 VDD.n969 VSS 0.00881f
C1211 VDD.n970 VSS 0.00937f
C1212 VDD.n971 VSS 0.0149f
C1213 VDD.n972 VSS 0.0142f
C1214 VDD.n973 VSS 0.0128f
C1215 VDD.n974 VSS 0.00122f
C1216 VDD.n975 VSS 0.0199f
C1217 VDD.n976 VSS 0.0414f
C1218 VDD.n977 VSS 0.0665f
C1219 VDD.t5 VSS 0.29f
C1220 VDD.n978 VSS 0.00954f
C1221 VDD.n979 VSS 0.00939f
C1222 VDD.n980 VSS 0.0933f
C1223 VDD.n981 VSS 0.541f
C1224 VDD.t8 VSS 1.91f
C1225 VDD.n982 VSS 0.00954f
C1226 VDD.n983 VSS 0.00939f
C1227 VDD.n984 VSS 0.0933f
C1228 VDD.n985 VSS 0.00954f
C1229 VDD.n986 VSS 0.00939f
C1230 VDD.n987 VSS 0.0933f
C1231 VDD.n988 VSS 0.00954f
C1232 VDD.n989 VSS 0.00939f
C1233 VDD.n990 VSS 0.0933f
C1234 VDD.n991 VSS 2.38f
C1235 VDD.t7 VSS 2.9f
C1236 VDD.n992 VSS 2.38f
C1237 VDD.t4 VSS 2.59f
C1238 VDD.n993 VSS 2.31f
C1239 VDD.n994 VSS 0.353f
C1240 VDD.n995 VSS 0.0727f
C1241 VDD.n996 VSS 0.0117f
C1242 VDD.n997 VSS 0.0199f
C1243 VDD.n998 VSS 0.00318f
C1244 VDD.n1000 VSS 0.00318f
C1245 VDD.n1001 VSS 3.63e-19
C1246 VDD.n1002 VSS 0.00308f
C1247 VDD.n1003 VSS 0.0105f
C1248 VDD.n1004 VSS 0.00472f
C1249 VDD.n1005 VSS 0.00671f
C1250 VDD.n1006 VSS 0.00925f
C1251 VDD.n1007 VSS 0.00762f
C1252 VDD.n1008 VSS 0.00381f
C1253 VDD.n1009 VSS 0.0112f
C1254 VDD.n1010 VSS 0.0112f
C1255 VDD.n1011 VSS 0.0148f
C1256 VDD.n1013 VSS 0.012f
C1257 VDD.n1014 VSS 3.63e-19
C1258 VDD.n1015 VSS 0.00399f
C1259 VDD.n1016 VSS 5.44e-19
C1260 VDD.n1017 VSS 0.00542f
C1261 VDD.n1018 VSS 0.00897f
C1262 VDD.n1019 VSS 0.00448f
C1263 VDD.n1020 VSS 0.0111f
C1264 VDD.n1021 VSS 0.0069f
C1265 VDD.n1022 VSS 0.00667f
C1266 VDD.n1023 VSS 3.74e-19
C1267 VDD.n1024 VSS 0.00542f
C1268 VDD.n1025 VSS 5.44e-19
C1269 VDD.n1026 VSS 0.00399f
C1270 VDD.n1027 VSS 0.00308f
C1271 VDD.n1028 VSS 0.00381f
C1272 VDD.n1029 VSS 0.0112f
C1273 VDD.n1030 VSS 0.0112f
C1274 VDD.n1031 VSS 0.0148f
C1275 VDD.n1032 VSS 0.00318f
C1276 VDD.n1034 VSS 0.012f
C1277 VDD.n1035 VSS 3.63e-19
C1278 VDD.n1036 VSS 0.00399f
C1279 VDD.n1037 VSS 5.44e-19
C1280 VDD.n1038 VSS 0.00542f
C1281 VDD.n1039 VSS 0.00897f
C1282 VDD.n1040 VSS 0.00448f
C1283 VDD.n1041 VSS 0.0111f
C1284 VDD.n1042 VSS 0.0069f
C1285 VDD.n1043 VSS -0.0987f
C1286 VDD.n1044 VSS 3.74e-19
C1287 VDD.n1045 VSS 0.00542f
C1288 VDD.n1046 VSS 5.44e-19
C1289 VDD.n1047 VSS 0.00399f
C1290 VDD.n1048 VSS 0.00308f
C1291 VDD.n1049 VSS 0.00381f
C1292 VDD.n1050 VSS 0.0112f
C1293 VDD.n1051 VSS 0.0112f
C1294 VDD.n1052 VSS 0.0148f
C1295 VDD.n1053 VSS 0.00318f
C1296 VDD.n1055 VSS 0.012f
C1297 VDD.n1056 VSS 3.63e-19
C1298 VDD.n1057 VSS 0.00399f
C1299 VDD.n1058 VSS 5.44e-19
C1300 VDD.n1059 VSS 0.00542f
C1301 VDD.n1060 VSS 0.00897f
C1302 VDD.n1061 VSS 0.00448f
C1303 VDD.n1062 VSS 0.0111f
C1304 VDD.n1063 VSS 0.0069f
C1305 VDD.n1064 VSS -0.0864f
C1306 VDD.n1065 VSS 0.00381f
C1307 VDD.n1066 VSS 0.0497f
C1308 VDD.n1067 VSS 0.0504f
C1309 VDD.n1068 VSS 0.0447f
C1310 VDD.n1069 VSS 0.0447f
C1311 VDD.n1070 VSS 0.0457f
C1312 VDD.n1071 VSS 0.0283f
C1313 VDD.n1072 VSS 0.00664f
C1314 VDD.n1073 VSS -0.099f
C1315 VDD.n1074 VSS 3.74e-19
C1316 VDD.n1075 VSS 0.00542f
C1317 VDD.n1076 VSS 5.44e-19
C1318 VDD.n1077 VSS 0.00399f
C1319 VDD.n1078 VSS 0.00308f
C1320 VDD.n1079 VSS 0.00381f
C1321 VDD.n1080 VSS 0.0112f
C1322 VDD.n1081 VSS 0.0112f
C1323 VDD.n1082 VSS 0.0148f
C1324 VDD.n1083 VSS 0.00318f
C1325 VDD.n1084 VSS 0.00308f
C1326 VDD.n1085 VSS 3.63e-19
C1327 VDD.n1086 VSS 0.012f
C1328 VDD.n1087 VSS 0.00318f
C1329 VDD.n1088 VSS 0.00308f
C1330 VDD.n1089 VSS 0.0105f
C1331 VDD.n1090 VSS 0.00472f
C1332 VDD.n1091 VSS 0.00671f
C1333 VDD.n1092 VSS 0.00925f
C1334 VDD.n1093 VSS 0.00762f
C1335 VDD.n1094 VSS 0.00381f
C1336 VDD.n1095 VSS 0.0112f
C1337 VDD.n1096 VSS 0.0112f
C1338 VDD.n1097 VSS 0.0148f
C1339 VDD.n1098 VSS 0.012f
C1340 VDD.n1099 VSS 3.63e-19
C1341 VDD.n1100 VSS 0.00399f
C1342 VDD.n1101 VSS 5.44e-19
C1343 VDD.n1102 VSS 0.00542f
C1344 VDD.n1103 VSS 0.00897f
C1345 VDD.n1104 VSS 0.00448f
C1346 VDD.n1105 VSS 0.0107f
C1347 VDD.n1106 VSS 0.00664f
C1348 VDD.n1107 VSS 0.00643f
C1349 VDD.n1108 VSS 3.74e-19
C1350 VDD.n1109 VSS 0.00542f
C1351 VDD.n1110 VSS 5.44e-19
C1352 VDD.n1111 VSS 0.00399f
C1353 VDD.n1112 VSS 0.00308f
C1354 VDD.n1113 VSS 0.00381f
C1355 VDD.n1114 VSS 0.0112f
C1356 VDD.n1115 VSS 0.0112f
C1357 VDD.n1116 VSS 0.0148f
C1358 VDD.n1117 VSS 0.00318f
C1359 VDD.n1118 VSS 0.00308f
C1360 VDD.n1119 VSS 3.63e-19
C1361 VDD.n1120 VSS 0.012f
C1362 VDD.n1121 VSS 0.00318f
C1363 VDD.n1122 VSS 0.00308f
C1364 VDD.n1123 VSS 0.0105f
C1365 VDD.n1124 VSS 0.00472f
C1366 VDD.n1125 VSS 0.00671f
C1367 VDD.n1126 VSS 0.00925f
C1368 VDD.n1127 VSS 0.00762f
C1369 VDD.n1128 VSS 0.00381f
C1370 VDD.n1129 VSS 0.0112f
C1371 VDD.n1130 VSS 0.0112f
C1372 VDD.n1131 VSS 0.0148f
C1373 VDD.n1132 VSS 0.012f
C1374 VDD.n1133 VSS 3.63e-19
C1375 VDD.n1134 VSS 0.00399f
C1376 VDD.n1135 VSS 5.44e-19
C1377 VDD.n1136 VSS 0.00542f
C1378 VDD.n1137 VSS 0.00897f
C1379 VDD.n1138 VSS 0.00448f
C1380 VDD.n1139 VSS 0.0107f
C1381 VDD.n1140 VSS 0.00664f
C1382 VDD.n1141 VSS 0.00643f
C1383 VDD.n1142 VSS 3.74e-19
C1384 VDD.n1143 VSS 0.00542f
C1385 VDD.n1144 VSS 5.44e-19
C1386 VDD.n1145 VSS 0.00399f
C1387 VDD.n1146 VSS 0.00308f
C1388 VDD.n1147 VSS 0.00381f
C1389 VDD.n1148 VSS 0.0112f
C1390 VDD.n1149 VSS 0.0112f
C1391 VDD.n1150 VSS 0.0148f
C1392 VDD.n1151 VSS 0.00318f
C1393 VDD.n1152 VSS 0.00308f
C1394 VDD.n1153 VSS 6.06e-19
C1395 VDD.n1154 VSS 0.00308f
C1396 VDD.n1155 VSS 0.00308f
C1397 VDD.n1156 VSS 0.00399f
C1398 VDD.n1157 VSS 0.0328f
C1399 VDD.n1158 VSS 0.0328f
C1400 VDD.n1159 VSS 0.0299f
C1401 VDD.n1160 VSS 0.00381f
C1402 VDD.n1161 VSS 0.0337f
C1403 VDD.n1162 VSS 0.00308f
C1404 VDD.n1163 VSS 6.06e-19
C1405 VDD.n1164 VSS 0.00399f
C1406 VDD.n1165 VSS 5.44e-19
C1407 VDD.n1166 VSS 0.00381f
C1408 VDD.n1167 VSS -0.0864f
C1409 VDD.n1168 VSS -0.243f
C1410 VDD.n1169 VSS 0.00671f
C1411 VDD.n1170 VSS 0.00925f
C1412 VDD.n1171 VSS 0.00762f
C1413 VDD.n1172 VSS 0.00381f
C1414 VDD.n1173 VSS 0.0112f
C1415 VDD.n1174 VSS 0.00308f
C1416 VDD.n1175 VSS 0.00318f
C1417 VDD.n1176 VSS 0.012f
C1418 VDD.n1177 VSS 3.63e-19
C1419 VDD.n1178 VSS 0.00399f
C1420 VDD.n1179 VSS 5.44e-19
C1421 VDD.n1180 VSS 0.00381f
C1422 VDD.n1181 VSS 0.00505f
C1423 VDD.n1182 VSS 0.00542f
C1424 VDD.n1183 VSS 0.00671f
C1425 VDD.n1184 VSS 0.00925f
C1426 VDD.n1185 VSS 0.00762f
C1427 VDD.n1186 VSS 0.00381f
C1428 VDD.n1187 VSS 0.0112f
C1429 VDD.n1188 VSS 0.00308f
C1430 VDD.n1189 VSS 3.63e-19
C1431 VDD.n1190 VSS 0.00399f
C1432 VDD.n1191 VSS 5.44e-19
C1433 VDD.n1192 VSS 0.00381f
C1434 VDD.n1193 VSS 0.00505f
C1435 VDD.n1194 VSS 0.00542f
C1436 VDD.n1195 VSS 0.00671f
C1437 VDD.n1196 VSS 0.00925f
C1438 VDD.n1197 VSS 0.00762f
C1439 VDD.n1198 VSS 0.00381f
C1440 VDD.n1199 VSS 0.0112f
C1441 VDD.n1200 VSS 0.00308f
C1442 VDD.n1201 VSS 3.63e-19
C1443 VDD.n1202 VSS 0.00399f
C1444 VDD.n1203 VSS 5.44e-19
C1445 VDD.n1204 VSS 0.00381f
C1446 VDD.n1205 VSS -0.0864f
C1447 VDD.n1206 VSS -0.243f
C1448 VDD.n1207 VSS 0.00671f
C1449 VDD.n1208 VSS 0.00925f
C1450 VDD.n1209 VSS 0.00762f
C1451 VDD.n1210 VSS 0.00381f
C1452 VDD.n1211 VSS 0.0112f
C1453 VDD.n1212 VSS 0.00308f
C1454 VDD.n1213 VSS 3.63e-19
C1455 VDD.n1214 VSS 0.00399f
C1456 VDD.n1215 VSS 5.44e-19
C1457 VDD.n1216 VSS 0.00381f
C1458 VDD.n1217 VSS 0.00505f
C1459 VDD.n1218 VSS 0.00542f
C1460 VDD.n1219 VSS 0.00671f
C1461 VDD.n1220 VSS 0.00925f
C1462 VDD.n1221 VSS 0.00762f
C1463 VDD.n1222 VSS 0.00381f
C1464 VDD.n1223 VSS 0.0112f
C1465 VDD.n1224 VSS 0.00308f
C1466 VDD.n1225 VSS 3.63e-19
C1467 VDD.n1226 VSS 0.00399f
C1468 VDD.n1227 VSS 5.44e-19
C1469 VDD.n1228 VSS 0.00381f
C1470 VDD.n1229 VSS 0.00505f
C1471 VDD.n1230 VSS 0.00643f
C1472 VDD.n1231 VSS 0.00664f
C1473 VDD.n1232 VSS 0.0277f
C1474 VDD.n1233 VSS 0.0278f
C1475 VDD.n1234 VSS 0.0283f
C1476 VDD.n1235 VSS 0.00664f
C1477 VDD.n1236 VSS -0.099f
C1478 VDD.n1237 VSS 3.74e-19
C1479 VDD.n1238 VSS 0.00542f
C1480 VDD.n1239 VSS 5.44e-19
C1481 VDD.n1240 VSS 0.00399f
C1482 VDD.n1241 VSS 0.00308f
C1483 VDD.n1242 VSS 0.00381f
C1484 VDD.n1243 VSS 0.0112f
C1485 VDD.n1244 VSS 0.0112f
C1486 VDD.n1245 VSS 0.0148f
C1487 VDD.n1246 VSS 0.00318f
C1488 VDD.n1247 VSS 0.00308f
C1489 VDD.n1248 VSS 3.63e-19
C1490 VDD.n1249 VSS 0.012f
C1491 VDD.n1250 VSS 0.00318f
C1492 VDD.n1251 VSS 0.00308f
C1493 VDD.n1252 VSS 0.0105f
C1494 VDD.n1253 VSS 0.00472f
C1495 VDD.n1254 VSS 0.00671f
C1496 VDD.n1255 VSS 0.00925f
C1497 VDD.n1256 VSS 0.00762f
C1498 VDD.n1257 VSS 0.00381f
C1499 VDD.n1258 VSS 0.0112f
C1500 VDD.n1259 VSS 0.0112f
C1501 VDD.n1260 VSS 0.0148f
C1502 VDD.n1261 VSS 0.012f
C1503 VDD.n1262 VSS 3.63e-19
C1504 VDD.n1263 VSS 0.00399f
C1505 VDD.n1264 VSS 5.44e-19
C1506 VDD.n1265 VSS 0.00542f
C1507 VDD.n1266 VSS 0.00897f
C1508 VDD.n1267 VSS 0.00448f
C1509 VDD.n1268 VSS 0.0107f
C1510 VDD.n1269 VSS 0.00664f
C1511 VDD.n1270 VSS 0.00643f
C1512 VDD.n1271 VSS 3.74e-19
C1513 VDD.n1272 VSS 0.00542f
C1514 VDD.n1273 VSS 5.44e-19
C1515 VDD.n1274 VSS 0.00399f
C1516 VDD.n1275 VSS 0.00308f
C1517 VDD.n1276 VSS 0.00381f
C1518 VDD.n1277 VSS 0.0112f
C1519 VDD.n1278 VSS 0.0112f
C1520 VDD.n1279 VSS 0.0148f
C1521 VDD.n1280 VSS 0.00318f
C1522 VDD.n1281 VSS 0.00308f
C1523 VDD.n1282 VSS 3.63e-19
C1524 VDD.n1283 VSS 0.012f
C1525 VDD.n1284 VSS 0.00318f
C1526 VDD.n1285 VSS 0.00308f
C1527 VDD.n1286 VSS 0.0105f
C1528 VDD.n1287 VSS 0.00472f
C1529 VDD.n1288 VSS 0.00671f
C1530 VDD.n1289 VSS 0.00925f
C1531 VDD.n1290 VSS 0.00762f
C1532 VDD.n1291 VSS 0.00381f
C1533 VDD.n1292 VSS 0.0112f
C1534 VDD.n1293 VSS 0.0112f
C1535 VDD.n1294 VSS 0.0148f
C1536 VDD.n1295 VSS 0.012f
C1537 VDD.n1296 VSS 3.63e-19
C1538 VDD.n1297 VSS 0.00399f
C1539 VDD.n1298 VSS 5.44e-19
C1540 VDD.n1299 VSS 0.00542f
C1541 VDD.n1300 VSS 0.00897f
C1542 VDD.n1301 VSS 0.00448f
C1543 VDD.n1302 VSS 0.0107f
C1544 VDD.n1303 VSS 0.00664f
C1545 VDD.n1304 VSS 0.00643f
C1546 VDD.n1305 VSS 3.74e-19
C1547 VDD.n1306 VSS 0.00542f
C1548 VDD.n1307 VSS 5.44e-19
C1549 VDD.n1308 VSS 0.00399f
C1550 VDD.n1309 VSS 0.00308f
C1551 VDD.n1310 VSS 0.00381f
C1552 VDD.n1311 VSS 0.0112f
C1553 VDD.n1312 VSS 0.0112f
C1554 VDD.n1313 VSS 0.0148f
C1555 VDD.n1314 VSS 0.00318f
C1556 VDD.n1315 VSS 0.00308f
C1557 VDD.n1316 VSS 6.06e-19
C1558 VDD.n1317 VSS 0.00308f
C1559 VDD.n1318 VSS 0.00308f
C1560 VDD.n1319 VSS 0.00399f
C1561 VDD.n1320 VSS 0.0328f
C1562 VDD.n1321 VSS 0.0328f
C1563 VDD.n1322 VSS 0.0299f
C1564 VDD.n1323 VSS 0.00381f
C1565 VDD.n1324 VSS 0.0337f
C1566 VDD.n1325 VSS 0.00308f
C1567 VDD.n1326 VSS 6.06e-19
C1568 VDD.n1327 VSS 0.00399f
C1569 VDD.n1328 VSS 5.44e-19
C1570 VDD.n1329 VSS 0.00381f
C1571 VDD.n1330 VSS -0.0864f
C1572 VDD.n1331 VSS -0.243f
C1573 VDD.n1332 VSS 0.00671f
C1574 VDD.n1333 VSS 0.00925f
C1575 VDD.n1334 VSS 0.00762f
C1576 VDD.n1335 VSS 0.00381f
C1577 VDD.n1336 VSS 0.0112f
C1578 VDD.n1337 VSS 0.00308f
C1579 VDD.n1338 VSS 0.00318f
C1580 VDD.n1339 VSS 0.012f
C1581 VDD.n1340 VSS 3.63e-19
C1582 VDD.n1341 VSS 0.00399f
C1583 VDD.n1342 VSS 5.44e-19
C1584 VDD.n1343 VSS 0.00381f
C1585 VDD.n1344 VSS 0.00505f
C1586 VDD.n1345 VSS 0.00542f
C1587 VDD.n1346 VSS 0.00671f
C1588 VDD.n1347 VSS 0.00925f
C1589 VDD.n1348 VSS 0.00762f
C1590 VDD.n1349 VSS 0.00381f
C1591 VDD.n1350 VSS 0.0112f
C1592 VDD.n1351 VSS 0.00308f
C1593 VDD.n1352 VSS 3.63e-19
C1594 VDD.n1353 VSS 0.00399f
C1595 VDD.n1354 VSS 5.44e-19
C1596 VDD.n1355 VSS 0.00381f
C1597 VDD.n1356 VSS 0.00505f
C1598 VDD.n1357 VSS 0.00542f
C1599 VDD.n1358 VSS 0.00671f
C1600 VDD.n1359 VSS 0.00925f
C1601 VDD.n1360 VSS 0.00762f
C1602 VDD.n1361 VSS 0.00381f
C1603 VDD.n1362 VSS 0.0112f
C1604 VDD.n1363 VSS 0.00308f
C1605 VDD.n1364 VSS 3.63e-19
C1606 VDD.n1365 VSS 0.00399f
C1607 VDD.n1366 VSS 5.44e-19
C1608 VDD.n1367 VSS 0.00381f
C1609 VDD.n1368 VSS -0.0864f
C1610 VDD.n1369 VSS -0.243f
C1611 VDD.n1370 VSS 0.00671f
C1612 VDD.n1371 VSS 0.00925f
C1613 VDD.n1372 VSS 0.00762f
C1614 VDD.n1373 VSS 0.00381f
C1615 VDD.n1374 VSS 0.0112f
C1616 VDD.n1375 VSS 0.00308f
C1617 VDD.n1376 VSS 3.63e-19
C1618 VDD.n1377 VSS 0.00399f
C1619 VDD.n1378 VSS 5.44e-19
C1620 VDD.n1379 VSS 0.00381f
C1621 VDD.n1380 VSS 0.00505f
C1622 VDD.n1381 VSS 0.00542f
C1623 VDD.n1382 VSS 0.00671f
C1624 VDD.n1383 VSS 0.00925f
C1625 VDD.n1384 VSS 0.00762f
C1626 VDD.n1385 VSS 0.00381f
C1627 VDD.n1386 VSS 0.0112f
C1628 VDD.n1387 VSS 0.00308f
C1629 VDD.n1388 VSS 3.63e-19
C1630 VDD.n1389 VSS 0.00399f
C1631 VDD.n1390 VSS 5.44e-19
C1632 VDD.n1391 VSS 0.00381f
C1633 VDD.n1392 VSS 0.00505f
C1634 VDD.n1393 VSS 0.00643f
C1635 VDD.n1394 VSS 0.00664f
C1636 VDD.n1395 VSS 0.0277f
C1637 VDD.n1396 VSS 0.0278f
C1638 VDD.n1397 VSS 0.0283f
C1639 VDD.n1398 VSS 0.00664f
C1640 VDD.n1399 VSS -0.099f
C1641 VDD.n1400 VSS 3.74e-19
C1642 VDD.n1401 VSS 0.00542f
C1643 VDD.n1402 VSS 5.44e-19
C1644 VDD.n1403 VSS 0.00399f
C1645 VDD.n1404 VSS 0.00308f
C1646 VDD.n1405 VSS 0.00381f
C1647 VDD.n1406 VSS 0.0112f
C1648 VDD.n1407 VSS 0.0112f
C1649 VDD.n1408 VSS 0.0148f
C1650 VDD.n1409 VSS 0.00318f
C1651 VDD.n1410 VSS 0.00308f
C1652 VDD.n1411 VSS 3.63e-19
C1653 VDD.n1412 VSS 0.012f
C1654 VDD.n1413 VSS 0.00318f
C1655 VDD.n1414 VSS 0.00308f
C1656 VDD.n1415 VSS 0.0105f
C1657 VDD.n1416 VSS 0.00472f
C1658 VDD.n1417 VSS 0.00671f
C1659 VDD.n1418 VSS 0.00925f
C1660 VDD.n1419 VSS 0.00762f
C1661 VDD.n1420 VSS 0.00381f
C1662 VDD.n1421 VSS 0.0112f
C1663 VDD.n1422 VSS 0.0112f
C1664 VDD.n1423 VSS 0.0148f
C1665 VDD.n1424 VSS 0.012f
C1666 VDD.n1425 VSS 3.63e-19
C1667 VDD.n1426 VSS 0.00399f
C1668 VDD.n1427 VSS 5.44e-19
C1669 VDD.n1428 VSS 0.00542f
C1670 VDD.n1429 VSS 0.00897f
C1671 VDD.n1430 VSS 0.00448f
C1672 VDD.n1431 VSS 0.0107f
C1673 VDD.n1432 VSS 0.00664f
C1674 VDD.n1433 VSS 0.00643f
C1675 VDD.n1434 VSS 3.74e-19
C1676 VDD.n1435 VSS 0.00542f
C1677 VDD.n1436 VSS 5.44e-19
C1678 VDD.n1437 VSS 0.00399f
C1679 VDD.n1438 VSS 0.00308f
C1680 VDD.n1439 VSS 0.00381f
C1681 VDD.n1440 VSS 0.0112f
C1682 VDD.n1441 VSS 0.0112f
C1683 VDD.n1442 VSS 0.0148f
C1684 VDD.n1443 VSS 0.00318f
C1685 VDD.n1444 VSS 0.00308f
C1686 VDD.n1445 VSS 3.63e-19
C1687 VDD.n1446 VSS 0.012f
C1688 VDD.n1447 VSS 0.00318f
C1689 VDD.n1448 VSS 0.00308f
C1690 VDD.n1449 VSS 0.0105f
C1691 VDD.n1450 VSS 0.00472f
C1692 VDD.n1451 VSS 0.00671f
C1693 VDD.n1452 VSS 0.00925f
C1694 VDD.n1453 VSS 0.00762f
C1695 VDD.n1454 VSS 0.00381f
C1696 VDD.n1455 VSS 0.0112f
C1697 VDD.n1456 VSS 0.0112f
C1698 VDD.n1457 VSS 0.0148f
C1699 VDD.n1458 VSS 0.012f
C1700 VDD.n1459 VSS 3.63e-19
C1701 VDD.n1460 VSS 0.00399f
C1702 VDD.n1461 VSS 5.44e-19
C1703 VDD.n1462 VSS 0.00542f
C1704 VDD.n1463 VSS 0.00897f
C1705 VDD.n1464 VSS 0.00448f
C1706 VDD.n1465 VSS 0.0107f
C1707 VDD.n1466 VSS 0.00664f
C1708 VDD.n1467 VSS 0.00643f
C1709 VDD.n1468 VSS 3.74e-19
C1710 VDD.n1469 VSS 0.00542f
C1711 VDD.n1470 VSS 5.44e-19
C1712 VDD.n1471 VSS 0.00399f
C1713 VDD.n1472 VSS 0.00308f
C1714 VDD.n1473 VSS 0.00381f
C1715 VDD.n1474 VSS 0.0112f
C1716 VDD.n1475 VSS 0.0112f
C1717 VDD.n1476 VSS 0.0148f
C1718 VDD.n1477 VSS 0.00318f
C1719 VDD.n1478 VSS 0.00308f
C1720 VDD.n1479 VSS 6.06e-19
C1721 VDD.n1480 VSS 0.00308f
C1722 VDD.n1481 VSS 0.00308f
C1723 VDD.n1482 VSS 0.00399f
C1724 VDD.n1483 VSS 0.0328f
C1725 VDD.n1484 VSS 0.0328f
C1726 VDD.n1485 VSS 0.0299f
C1727 VDD.n1486 VSS 0.00381f
C1728 VDD.n1487 VSS 0.0337f
C1729 VDD.n1488 VSS 0.00308f
C1730 VDD.n1489 VSS 6.06e-19
C1731 VDD.n1490 VSS 0.00399f
C1732 VDD.n1491 VSS 5.44e-19
C1733 VDD.n1492 VSS 0.00381f
C1734 VDD.n1493 VSS -0.0864f
C1735 VDD.n1494 VSS -0.243f
C1736 VDD.n1495 VSS 0.00671f
C1737 VDD.n1496 VSS 0.00925f
C1738 VDD.n1497 VSS 0.00762f
C1739 VDD.n1498 VSS 0.00381f
C1740 VDD.n1499 VSS 0.0112f
C1741 VDD.n1500 VSS 0.00308f
C1742 VDD.n1501 VSS 0.00318f
C1743 VDD.n1502 VSS 0.012f
C1744 VDD.n1503 VSS 3.63e-19
C1745 VDD.n1504 VSS 0.00399f
C1746 VDD.n1505 VSS 5.44e-19
C1747 VDD.n1506 VSS 0.00381f
C1748 VDD.n1507 VSS 0.00505f
C1749 VDD.n1508 VSS 0.00542f
C1750 VDD.n1509 VSS 0.00671f
C1751 VDD.n1510 VSS 0.00925f
C1752 VDD.n1511 VSS 0.00762f
C1753 VDD.n1512 VSS 0.00381f
C1754 VDD.n1513 VSS 0.0112f
C1755 VDD.n1514 VSS 0.00308f
C1756 VDD.n1515 VSS 3.63e-19
C1757 VDD.n1516 VSS 0.00399f
C1758 VDD.n1517 VSS 5.44e-19
C1759 VDD.n1518 VSS 0.00381f
C1760 VDD.n1519 VSS 0.00505f
C1761 VDD.n1520 VSS 0.00542f
C1762 VDD.n1521 VSS 0.00671f
C1763 VDD.n1522 VSS 0.00925f
C1764 VDD.n1523 VSS 0.00762f
C1765 VDD.n1524 VSS 0.00381f
C1766 VDD.n1525 VSS 0.0112f
C1767 VDD.n1526 VSS 0.00308f
C1768 VDD.n1527 VSS 3.63e-19
C1769 VDD.n1528 VSS 0.00399f
C1770 VDD.n1529 VSS 5.44e-19
C1771 VDD.n1530 VSS 0.00381f
C1772 VDD.n1531 VSS -0.0864f
C1773 VDD.n1532 VSS -0.243f
C1774 VDD.n1533 VSS 0.00671f
C1775 VDD.n1534 VSS 0.00925f
C1776 VDD.n1535 VSS 0.00762f
C1777 VDD.n1536 VSS 0.00381f
C1778 VDD.n1537 VSS 0.0112f
C1779 VDD.n1538 VSS 0.00308f
C1780 VDD.n1539 VSS 3.63e-19
C1781 VDD.n1540 VSS 0.00399f
C1782 VDD.n1541 VSS 5.44e-19
C1783 VDD.n1542 VSS 0.00381f
C1784 VDD.n1543 VSS 0.00505f
C1785 VDD.n1544 VSS 0.00542f
C1786 VDD.n1545 VSS 0.00671f
C1787 VDD.n1546 VSS 0.00925f
C1788 VDD.n1547 VSS 0.00762f
C1789 VDD.n1548 VSS 0.00381f
C1790 VDD.n1549 VSS 0.0112f
C1791 VDD.n1550 VSS 0.00308f
C1792 VDD.n1551 VSS 3.63e-19
C1793 VDD.n1552 VSS 0.00399f
C1794 VDD.n1553 VSS 5.44e-19
C1795 VDD.n1554 VSS 0.00381f
C1796 VDD.n1555 VSS 0.00505f
C1797 VDD.n1556 VSS 0.00643f
C1798 VDD.n1557 VSS 0.00664f
C1799 VDD.n1558 VSS 0.0277f
C1800 VDD.n1559 VSS 0.0278f
C1801 VDD.n1560 VSS 0.0283f
C1802 VDD.n1561 VSS 0.00664f
C1803 VDD.n1562 VSS -0.099f
C1804 VDD.n1563 VSS 3.74e-19
C1805 VDD.n1564 VSS 0.00542f
C1806 VDD.n1565 VSS 5.44e-19
C1807 VDD.n1566 VSS 0.00399f
C1808 VDD.n1567 VSS 0.00308f
C1809 VDD.n1568 VSS 0.00381f
C1810 VDD.n1569 VSS 0.0112f
C1811 VDD.n1570 VSS 0.0112f
C1812 VDD.n1571 VSS 0.0148f
C1813 VDD.n1572 VSS 0.00318f
C1814 VDD.n1573 VSS 0.00308f
C1815 VDD.n1574 VSS 3.63e-19
C1816 VDD.n1575 VSS 0.012f
C1817 VDD.n1576 VSS 0.00318f
C1818 VDD.n1577 VSS 0.00308f
C1819 VDD.n1578 VSS 0.0105f
C1820 VDD.n1579 VSS 0.00472f
C1821 VDD.n1580 VSS 0.00671f
C1822 VDD.n1581 VSS 0.00925f
C1823 VDD.n1582 VSS 0.00762f
C1824 VDD.n1583 VSS 0.00381f
C1825 VDD.n1584 VSS 0.0112f
C1826 VDD.n1585 VSS 0.0112f
C1827 VDD.n1586 VSS 0.0148f
C1828 VDD.n1587 VSS 0.012f
C1829 VDD.n1588 VSS 3.63e-19
C1830 VDD.n1589 VSS 0.00399f
C1831 VDD.n1590 VSS 5.44e-19
C1832 VDD.n1591 VSS 0.00542f
C1833 VDD.n1592 VSS 0.00897f
C1834 VDD.n1593 VSS 0.00448f
C1835 VDD.n1594 VSS 0.0107f
C1836 VDD.n1595 VSS 0.00664f
C1837 VDD.n1596 VSS 0.00643f
C1838 VDD.n1597 VSS 3.74e-19
C1839 VDD.n1598 VSS 0.00542f
C1840 VDD.n1599 VSS 5.44e-19
C1841 VDD.n1600 VSS 0.00399f
C1842 VDD.n1601 VSS 0.00308f
C1843 VDD.n1602 VSS 0.00381f
C1844 VDD.n1603 VSS 0.0112f
C1845 VDD.n1604 VSS 0.0112f
C1846 VDD.n1605 VSS 0.0148f
C1847 VDD.n1606 VSS 0.00318f
C1848 VDD.n1607 VSS 0.00308f
C1849 VDD.n1608 VSS 3.63e-19
C1850 VDD.n1609 VSS 0.012f
C1851 VDD.n1610 VSS 0.00318f
C1852 VDD.n1611 VSS 0.00308f
C1853 VDD.n1612 VSS 0.0105f
C1854 VDD.n1613 VSS 0.00472f
C1855 VDD.n1614 VSS 0.00671f
C1856 VDD.n1615 VSS 0.00925f
C1857 VDD.n1616 VSS 0.00762f
C1858 VDD.n1617 VSS 0.00381f
C1859 VDD.n1618 VSS 0.0112f
C1860 VDD.n1619 VSS 0.0112f
C1861 VDD.n1620 VSS 0.0148f
C1862 VDD.n1621 VSS 0.012f
C1863 VDD.n1622 VSS 3.63e-19
C1864 VDD.n1623 VSS 0.00399f
C1865 VDD.n1624 VSS 5.44e-19
C1866 VDD.n1625 VSS 0.00542f
C1867 VDD.n1626 VSS 0.00897f
C1868 VDD.n1627 VSS 0.00448f
C1869 VDD.n1628 VSS 0.0107f
C1870 VDD.n1629 VSS 0.00664f
C1871 VDD.n1630 VSS 0.00643f
C1872 VDD.n1631 VSS 3.74e-19
C1873 VDD.n1632 VSS 0.00542f
C1874 VDD.n1633 VSS 5.44e-19
C1875 VDD.n1634 VSS 0.00399f
C1876 VDD.n1635 VSS 0.00308f
C1877 VDD.n1636 VSS 0.00381f
C1878 VDD.n1637 VSS 0.0112f
C1879 VDD.n1638 VSS 0.0112f
C1880 VDD.n1639 VSS 0.0148f
C1881 VDD.n1640 VSS 0.00318f
C1882 VDD.n1641 VSS 0.00308f
C1883 VDD.n1642 VSS 6.06e-19
C1884 VDD.n1643 VSS 0.00308f
C1885 VDD.n1644 VSS 0.00308f
C1886 VDD.n1645 VSS 0.00399f
C1887 VDD.n1646 VSS 0.0328f
C1888 VDD.n1647 VSS 0.0328f
C1889 VDD.n1648 VSS 0.0299f
C1890 VDD.n1649 VSS 0.00381f
C1891 VDD.n1650 VSS 0.0337f
C1892 VDD.n1651 VSS 0.00308f
C1893 VDD.n1652 VSS 6.06e-19
C1894 VDD.n1653 VSS 0.00399f
C1895 VDD.n1654 VSS 5.44e-19
C1896 VDD.n1655 VSS 0.00381f
C1897 VDD.n1656 VSS -0.0864f
C1898 VDD.n1657 VSS -0.243f
C1899 VDD.n1658 VSS 0.00671f
C1900 VDD.n1659 VSS 0.00925f
C1901 VDD.n1660 VSS 0.00762f
C1902 VDD.n1661 VSS 0.00381f
C1903 VDD.n1662 VSS 0.0112f
C1904 VDD.n1663 VSS 0.00308f
C1905 VDD.n1664 VSS 0.00318f
C1906 VDD.n1665 VSS 0.012f
C1907 VDD.n1666 VSS 3.63e-19
C1908 VDD.n1667 VSS 0.00399f
C1909 VDD.n1668 VSS 0.0105f
C1910 VDD.n1669 VSS 0.00472f
C1911 VDD.n1670 VSS 0.00671f
C1912 VDD.n1671 VSS 0.00542f
C1913 VDD.n1672 VSS 0.0043f
C1914 VDD.n1673 VSS 0.00916f
C1915 VDD.n1674 VSS -0.216f
C1916 VDD.n1675 VSS -0.107f
C1917 VDD.n1676 VSS 0.00643f
C1918 VDD.n1677 VSS 0.00505f
C1919 VDD.n1678 VSS 0.00381f
C1920 VDD.n1679 VSS 0.00472f
C1921 VDD.n1680 VSS 0.0105f
C1922 VDD.n1681 VSS 0.00762f
C1923 VDD.n1682 VSS 0.00925f
C1924 VDD.n1683 VSS 0.00399f
C1925 VDD.n1684 VSS 0.00308f
C1926 VDD.n1685 VSS 0.00399f
C1927 VDD.n1686 VSS 3.63e-19
C1928 VDD.n1687 VSS 0.012f
C1929 VDD.n1688 VSS 2.92f
C1930 VDD.n1689 VSS 0.0232f
C1931 VDD.n1690 VSS 0.0592f
C1932 VDD.n1691 VSS 0.0484f
C1933 VDD.n1692 VSS 0.0447f
C1934 VDD.n1693 VSS 0.0457f
C1935 VDD.n1694 VSS 0.00667f
C1936 VDD.n1695 VSS 0.176f
C1937 VDD.n1696 VSS 0.0125f
C1938 VDD.n1697 VSS 0.0996f
C1939 VDD.n1698 VSS 0.0996f
C1940 VDD.n1699 VSS 0.0125f
C1941 VDD.n1700 VSS 0.107f
C1942 VDD.n1701 VSS 0.107f
C1943 VDD.n1702 VSS 0.0125f
C1944 VDD.n1703 VSS 0.122f
C1945 VDD.n1704 VSS 0.122f
C1946 VDD.n1705 VSS 0.0125f
C1947 VDD.n1706 VSS 0.111f
C1948 VDD.n1707 VSS 0.0524f
C1949 VDD.n1708 VSS 0.111f
C1950 VDD.n1709 VSS 0.0125f
C1951 VDD.n1710 VSS 0.00728f
C1952 VDD.n1711 VSS 0.00939f
C1953 VDD.n1712 VSS 0.0933f
C1954 VDD.n1713 VSS 1.82f
C1955 VDD.t17 VSS 0.492f
C1956 VDD.t11 VSS 1.03f
C1957 VDD.n1714 VSS 0.0179f
C1958 VDD.t2 VSS 2.54f
C1959 VDD.t0 VSS 7.66f
C1960 VDD.t14 VSS 5.87f
C1961 VDD.n1715 VSS 1.05f
C1962 VDD.t9 VSS 0.143f
C1963 VDD.n1716 VSS 0.0726f
C1964 VDD.n1717 VSS 0.0361f
C1965 VDD.n1718 VSS 0.00915f
C1966 VDD.n1719 VSS 0.00448f
C1967 VDD.n1720 VSS 0.0126f
C1968 VDD.n1721 VSS 0.0122f
C1969 VDD.n1722 VSS 0.0314f
C1970 VDD.n1723 VSS 0.0198f
C1971 VDD.n1724 VSS 0.0227f
C1972 VDD.n1725 VSS 9.36e-19
C1973 VDD.n1726 VSS 0.03f
C1974 VDD.n1727 VSS 0.023f
C1975 VDD.n1728 VSS 0.0276f
C1976 VDD.n1729 VSS 0.00459f
C1977 VDD.n1730 VSS 0.0142f
C1978 VDD.n1731 VSS 0.00529f
C1979 VDD.n1732 VSS 0.00554f
C1980 VDD.n1733 VSS 0.00211f
C1981 VDD.n1734 VSS 0.00156f
C1982 VDD.n1735 VSS 0.0124f
C1983 VDD.n1736 VSS 0.00294f
C1984 VDD.n1737 VSS 0.00187f
C1985 VDD.n1738 VSS 0.0171f
C1986 VDD.n1739 VSS 0.0867f
C1987 VDD.t12 VSS 0.118f
C1988 VDD.n1740 VSS 0.107f
C1989 VDD.n1741 VSS 0.0232f
C1990 VDD.n1742 VSS 0.00915f
C1991 VDD.n1743 VSS 0.0638f
C1992 VDD.n1744 VSS 0.0258f
C1993 x5[7].floating.n0 VSS -7.97f
C1994 x5[7].floating.n1 VSS -28.8f
C1995 x5[7].floating.n2 VSS 3.82f
C1996 x5[7].floating.n3 VSS -7.06f
C1997 x5[7].floating.n4 VSS -28.3f
C1998 x5[7].floating.n5 VSS 52.6f
C1999 x5[7].floating.n6 VSS -28.3f
C2000 x5[7].floating.n7 VSS -7.06f
C2001 x5[7].floating.n8 VSS 3.82f
C2002 x5[7].floating.n9 VSS -28.8f
C2003 x5[7].floating.n10 VSS -8f
C2004 x5[7].floating.n11 VSS 2.2f
C2005 x5[7].floating.t5 VSS 0.857f
C2006 x5[7].floating.n12 VSS 6.64f
C2007 x5[7].floating.n13 VSS 1.21f
C2008 x5[7].floating.n14 VSS 1.16f
C2009 x5[7].floating.n15 VSS 2.18f
C2010 x5[7].floating.n16 VSS 1.06f
C2011 x5[7].floating.n17 VSS 0.365f
C2012 x5[7].floating.n18 VSS 1.06f
C2013 x5[7].floating.n19 VSS 2.8f
C2014 x5[7].floating.n20 VSS 51.3f
C2015 x5[7].floating.n21 VSS 2.78f
C2016 x5[7].floating.n22 VSS 1.06f
C2017 x5[7].floating.n23 VSS 0.363f
C2018 x5[7].floating.t2 VSS 0.857f
C2019 x5[7].floating.n24 VSS 6.47f
C2020 x5[7].floating.n25 VSS 1.15f
C2021 x5[7].floating.n26 VSS 1.36f
C2022 x5[7].floating.n27 VSS 2.2f
C2023 x5[7].floating.n28 VSS 1.06f
C2024 x5[7].floating.n29 VSS 2.22f
C2025 x5[7].floating.n30 VSS -7.97f
C2026 x5[7].floating.n31 VSS -28.8f
C2027 x5[7].floating.n32 VSS 3.82f
C2028 x5[7].floating.n33 VSS -7.06f
C2029 x5[7].floating.n34 VSS -28.3f
C2030 x5[7].floating.n35 VSS 52.6f
C2031 x5[7].floating.n36 VSS -28.3f
C2032 x5[7].floating.n37 VSS -7.06f
C2033 x5[7].floating.n38 VSS 3.82f
C2034 x5[7].floating.n39 VSS -28.8f
C2035 x5[7].floating.n40 VSS -8f
C2036 x5[7].floating.n41 VSS 2.2f
C2037 x5[7].floating.t1 VSS 0.857f
C2038 x5[7].floating.n42 VSS 6.64f
C2039 x5[7].floating.n43 VSS 1.21f
C2040 x5[7].floating.n44 VSS 1.16f
C2041 x5[7].floating.n45 VSS 2.18f
C2042 x5[7].floating.n46 VSS 1.06f
C2043 x5[7].floating.n47 VSS 0.365f
C2044 x5[7].floating.n48 VSS 1.06f
C2045 x5[7].floating.n49 VSS 2.8f
C2046 x5[7].floating.n50 VSS 51.3f
C2047 x5[7].floating.n51 VSS 2.78f
C2048 x5[7].floating.n52 VSS 1.06f
C2049 x5[7].floating.n53 VSS 0.363f
C2050 x5[7].floating.t3 VSS 0.857f
C2051 x5[7].floating.n54 VSS 6.47f
C2052 x5[7].floating.n55 VSS 1.15f
C2053 x5[7].floating.n56 VSS 1.36f
C2054 x5[7].floating.n57 VSS 2.2f
C2055 x5[7].floating.n58 VSS 1.06f
C2056 x5[7].floating.n59 VSS -15.2f
C2057 x5[7].floating.n60 VSS -15.1f
C2058 x5[7].floating.n61 VSS -41.5f
C2059 x5[7].floating.n62 VSS 0.765f
C2060 x5[7].floating.n63 VSS 2.46f
C2061 x5[7].floating.n64 VSS 51.4f
C2062 x5[7].floating.n65 VSS 2.46f
C2063 x5[7].floating.n66 VSS 0.765f
C2064 x5[7].floating.n67 VSS -33.4f
C2065 x5[7].floating.n68 VSS -4.55f
C2066 x5[7].floating.n69 VSS 3.82f
C2067 x5[7].floating.n70 VSS -28.8f
C2068 x5[7].floating.n71 VSS -7.06f
C2069 x5[7].floating.n72 VSS 2.68f
C2070 x5[7].floating.n73 VSS 51.9f
C2071 x5[7].floating.n74 VSS 3.23f
C2072 x5[7].floating.n75 VSS -7.82f
C2073 x5[7].floating.n76 VSS -28.8f
C2074 x5[7].floating.n77 VSS 3.82f
C2075 x5[7].floating.n78 VSS -5f
C2076 x5[7].floating.n79 VSS -32.9f
C2077 x5[7].floating.n80 VSS 0.765f
C2078 x5[7].floating.n81 VSS 2.46f
C2079 x5[7].floating.n82 VSS 2.68f
C2080 x5[7].floating.n83 VSS -7.06f
C2081 x5[7].floating.n84 VSS -28.8f
C2082 x5[7].floating.n85 VSS 3.82f
C2083 x5[7].floating.n86 VSS -4.55f
C2084 x5[7].floating.n87 VSS -33.4f
C2085 x5[7].floating.n88 VSS 0.765f
C2086 x5[7].floating.n89 VSS 2.46f
C2087 x5[7].floating.n90 VSS 51.4f
C2088 x5[7].floating.n91 VSS 51.3f
C2089 x5[7].floating.n92 VSS 2.8f
C2090 x5[7].floating.n93 VSS 1.06f
C2091 x5[7].floating.n94 VSS 0.365f
C2092 x5[7].floating.t7 VSS 0.857f
C2093 x5[7].floating.n95 VSS 6.64f
C2094 x5[7].floating.n96 VSS 1.21f
C2095 x5[7].floating.n97 VSS 1.16f
C2096 x5[7].floating.n98 VSS 2.18f
C2097 x5[7].floating.n99 VSS 1.06f
C2098 x5[7].floating.n100 VSS 2.2f
C2099 x5[7].floating.n101 VSS -8f
C2100 x5[7].floating.n102 VSS -28.8f
C2101 x5[7].floating.n103 VSS 3.82f
C2102 x5[7].floating.n104 VSS -7.06f
C2103 x5[7].floating.n105 VSS -28.3f
C2104 x5[7].floating.n106 VSS 2.78f
C2105 x5[7].floating.n107 VSS 1.06f
C2106 x5[7].floating.n108 VSS 0.363f
C2107 x5[7].floating.t6 VSS 0.857f
C2108 x5[7].floating.n109 VSS 6.47f
C2109 x5[7].floating.n110 VSS 1.15f
C2110 x5[7].floating.n111 VSS 1.36f
C2111 x5[7].floating.n112 VSS 2.2f
C2112 x5[7].floating.n113 VSS 1.06f
C2113 x5[7].floating.n114 VSS 2.22f
C2114 x5[7].floating.n115 VSS -7.97f
C2115 x5[7].floating.n116 VSS -28.8f
C2116 x5[7].floating.n117 VSS 3.82f
C2117 x5[7].floating.n118 VSS -7.06f
C2118 x5[7].floating.n119 VSS -28.3f
C2119 x5[7].floating.n120 VSS 52.6f
C2120 x5[7].floating.n121 VSS 51.9f
C2121 x5[7].floating.n122 VSS 3.23f
C2122 x5[7].floating.n123 VSS -7.82f
C2123 x5[7].floating.n124 VSS -28.8f
C2124 x5[7].floating.n125 VSS 3.82f
C2125 x5[7].floating.n126 VSS -5f
C2126 x5[7].floating.n127 VSS -32.9f
C2127 x5[7].floating.n128 VSS 0.765f
C2128 x5[7].floating.n129 VSS 2.46f
C2129 x5[7].floating.n130 VSS 51.4f
C2130 x5[7].floating.n131 VSS 2.46f
C2131 x5[7].floating.n132 VSS 0.765f
C2132 x5[7].floating.n133 VSS -33.4f
C2133 x5[7].floating.n134 VSS -4.55f
C2134 x5[7].floating.n135 VSS 3.82f
C2135 x5[7].floating.n136 VSS -28.8f
C2136 x5[7].floating.n137 VSS -7.06f
C2137 x5[7].floating.n138 VSS 2.68f
C2138 x5[7].floating.n139 VSS 51.9f
C2139 x5[7].floating.n140 VSS 3.23f
C2140 x5[7].floating.n141 VSS 2.22f
C2141 x5[7].floating.t4 VSS 0.857f
C2142 x5[7].floating.n142 VSS 6.47f
C2143 x5[7].floating.n143 VSS 1.15f
C2144 x5[7].floating.n144 VSS 1.36f
C2145 x5[7].floating.n145 VSS 2.2f
C2146 x5[7].floating.n146 VSS 1.06f
C2147 x5[7].floating.n147 VSS 0.363f
C2148 x5[7].floating.n148 VSS 1.06f
C2149 x5[7].floating.n149 VSS 2.78f
C2150 x5[7].floating.n150 VSS 51.3f
C2151 x5[7].floating.n151 VSS 2.8f
C2152 x5[7].floating.n152 VSS 1.06f
C2153 x5[7].floating.n153 VSS 0.365f
C2154 x5[7].floating.t0 VSS 0.857f
C2155 x5[7].floating.n154 VSS 7.14f
C2156 x5[7].floating.n155 VSS 1.21f
C2157 x5[7].floating.n156 VSS 1.16f
C2158 x5[7].floating.n157 VSS 1.67f
C2159 x5[7].floating.n158 VSS 1.06f
C2160 x5[7].floating.n159 VSS -17.3f
C2161 x5[7].floating.n160 VSS -17.2f
C2162 x5[7].floating.n161 VSS -43.5f
C2163 x5[7].floating.n162 VSS 0.765f
C2164 x5[7].floating.n163 VSS 2.46f
C2165 x5[7].floating.n164 VSS 51.4f
C2166 x5[7].floating.n165 VSS 2.46f
C2167 x5[7].floating.n166 VSS 0.765f
C2168 x5[7].floating.n167 VSS -32.9f
C2169 x5[7].floating.n168 VSS -5f
C2170 x5[7].floating.n169 VSS 3.82f
C2171 x5[7].floating.n170 VSS -28.8f
C2172 x5[7].floating.n171 VSS -7.82f
C2173 x10.Y.t0 VSS 0.0462f
C2174 x10.Y.t6 VSS 0.0167f
C2175 x10.Y.t8 VSS 0.0167f
C2176 x10.Y.t7 VSS 0.0167f
C2177 x10.Y.t2 VSS 0.0167f
C2178 x10.Y.t3 VSS 0.0167f
C2179 x10.Y.t4 VSS 0.0167f
C2180 x10.Y.t5 VSS 0.0167f
C2181 x10.Y.t9 VSS 0.0167f
C2182 x10.Y.n0 VSS 0.222f
C2183 x10.Y.n1 VSS 0.0366f
C2184 x10.Y.t1 VSS 0.0174f
C2185 x10.Y.n2 VSS 0.0188f
C2186 x10.Y.n3 VSS 0.0186f
C2187 x10.Y.n4 VSS 0.0151f
C2188 x10.Y.n5 VSS 0.0211f
.ends

