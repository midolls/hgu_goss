magic
tech sky130A
magscale 1 2
timestamp 1698045515
<< checkpaint >>
rect -1313 2170 1629 2329
rect -1313 -713 2736 2170
rect -206 -872 2736 -713
<< error_s >>
rect 298 999 333 1016
rect 299 998 333 999
rect 299 962 369 998
rect 129 931 187 937
rect 129 897 141 931
rect 316 928 387 962
rect 667 928 702 962
rect 129 891 187 897
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 928
rect 668 909 702 928
rect 498 860 556 866
rect 498 826 510 860
rect 498 820 556 826
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 687 530 702 909
rect 721 875 756 909
rect 721 530 755 875
rect 867 807 925 813
rect 867 773 879 807
rect 867 767 925 773
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 0
transform 1 0 527 0 1 746
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM2
timestamp 0
transform 1 0 158 0 1 808
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_L7T3GD  XM3
timestamp 0
transform 1 0 896 0 1 693
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM4
timestamp 0
transform 1 0 1265 0 1 649
box -211 -261 211 261
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 B
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
