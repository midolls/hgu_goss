magic
tech sky130A
magscale 1 2
timestamp 1697025759
<< nwell >>
rect -346 -299 346 299
<< pmos >>
rect -150 -80 150 80
<< pdiff >>
rect -208 68 -150 80
rect -208 -68 -196 68
rect -162 -68 -150 68
rect -208 -80 -150 -68
rect 150 68 208 80
rect 150 -68 162 68
rect 196 -68 208 68
rect 150 -80 208 -68
<< pdiffc >>
rect -196 -68 -162 68
rect 162 -68 196 68
<< nsubdiff >>
rect -310 229 -214 263
rect 214 229 310 263
rect -310 167 -276 229
rect 276 167 310 229
rect -310 -229 -276 -167
rect 276 -229 310 -167
rect -310 -263 -214 -229
rect 214 -263 310 -229
<< nsubdiffcont >>
rect -214 229 214 263
rect -310 -167 -276 167
rect 276 -167 310 167
rect -214 -263 214 -229
<< poly >>
rect -150 161 150 177
rect -150 127 -134 161
rect 134 127 150 161
rect -150 80 150 127
rect -150 -127 150 -80
rect -150 -161 -134 -127
rect 134 -161 150 -127
rect -150 -177 150 -161
<< polycont >>
rect -134 127 134 161
rect -134 -161 134 -127
<< locali >>
rect -310 229 -214 263
rect 214 229 310 263
rect -310 167 -276 229
rect 276 167 310 229
rect -150 127 -134 161
rect 134 127 150 161
rect -196 68 -162 84
rect -196 -84 -162 -68
rect 162 68 196 84
rect 162 -84 196 -68
rect -150 -161 -134 -127
rect 134 -161 150 -127
rect -310 -229 -276 -167
rect 276 -229 310 -167
rect -310 -263 -214 -229
rect 214 -263 310 -229
<< viali >>
rect -134 127 134 161
rect -196 -68 -162 68
rect 162 -68 196 68
rect -134 -161 134 -127
<< metal1 >>
rect -146 161 146 167
rect -146 127 -134 161
rect 134 127 146 161
rect -146 121 146 127
rect -202 68 -156 80
rect -202 -68 -196 68
rect -162 -68 -156 68
rect -202 -80 -156 -68
rect 156 68 202 80
rect 156 -68 162 68
rect 196 -68 202 68
rect 156 -80 202 -68
rect -146 -127 146 -121
rect -146 -161 -134 -127
rect 134 -161 146 -127
rect -146 -167 146 -161
<< properties >>
string FIXED_BBOX -293 -246 293 246
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 1.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
